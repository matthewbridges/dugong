----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:14:21 07/26/2012 
-- Design Name: 
-- Module Name:    test_program - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library UNISIM;
use UNISIM.Vcomponents.all;

entity inst_mem is
	generic(
		DATA_WIDTH : natural := 32;
		ADDR_WIDTH : natural := 9
	);
	port(
		--Wishbone Slave Lines
		CLK_I : in  STD_LOGIC;
		RST_I : in  STD_LOGIC;
		DAT_I : in  STD_LOGIC_VECTOR(DATA_WIDTH - 1 downto 0);
		DAT_O : out STD_LOGIC_VECTOR(DATA_WIDTH - 1 downto 0);
		ADR_I : in  STD_LOGIC_VECTOR(ADDR_WIDTH - 1 downto 0);
		WE_I  : in  STD_LOGIC;
		STB_I : in  STD_LOGIC
	--		CYC_I : in   STD_LOGIC;

	);
end inst_mem;

architecture Behavioral of inst_mem is
	signal adr : std_logic_vector(13 downto 0);
	signal we  : std_logic_vector(3 downto 0);

begin

	-- RAMB16BWER: 16k-bit Data and 2k-bit Parity Configurable Synchronous Dual Port Block RAM with Optional Output Registers
	--             Spartan-6
	-- Xilinx HDL Libraries Guide, version 14.1

	RAMB16BWER_inst : RAMB16BWER
		generic map(
			DATA_WIDTH_A        => 36,  -- Valid values are 0, 1, 2, 4, 9, 18, or 36
			DATA_WIDTH_B        => 0,   -- Valid values are 0, 1, 2, 4, 9, 18, or 36
			DOA_REG             => 0,   -- Specifies to enable=1/disable=0 port A output registers
			DOB_REG             => 0,   -- Specifies to enable=1/disable=0 port B output registers
			INIT_A              => X"000000000", -- Initial values on A output port
			INIT_B              => X"000000000", -- Initial values on B output port
			INIT_FILE           => "inst_mem_data.mem", -- INIT_FILE: Optional file used to specify initial RAM contents
			-- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
			EN_RSTRAM_A         => TRUE,
			EN_RSTRAM_B         => FALSE,
			-- RSTTYPE: "SYNC" or "ASYNC"
			RSTTYPE             => "SYNC",
			-- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR"
			RST_PRIORITY_A      => "CE",
			RST_PRIORITY_B      => "CE",
			SIM_COLLISION_CHECK => "ALL", -- Collision check enable "ALL", "WARNING_ONLY", 
			--                               "GENERATE_X_ONLY" or "NONE"
			SIM_DEVICE          => "SPARTAN6", -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behaviour
			SRVAL_A             => X"000000000", -- Port A output value upon SSR assertion
			SRVAL_B             => X"000000000", -- Port B output value upon SSR assertion
			WRITE_MODE_A        => "WRITE_FIRST", -- WRITE_FIRST, READ_FIRST or NO_CHANGE
			WRITE_MODE_B        => "WRITE_FIRST", -- WRITE_FIRST, READ_FIRST or NO_CHANGE
			-- INITP_00 to INITP_07: Initial memory contents.
			INITP_00            => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_01            => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_02            => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_03            => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_04            => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_05            => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_06            => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_07            => X"0000000000000000000000000000000000000000000000000000000000000000",
			-- INIT_00 to INIT_3F: Initial memory contents.
			INIT_00             => X"00000000000000000000000000000000000000000000000000000000400000D8", --0x00
			INIT_01             => X"801FAF081F080003801FAF081F080002801FAF081F080001801FAF081F080000", --0x08
			INIT_02             => X"801FAF081F080007801FAF081F080006801FAF081F080005801FAF081F080004", --0x10
			INIT_03             => X"801FAF081F08000B801FAF081F08000A801FAF081F080009801FAF081F080008", --0x18
			INIT_04             => X"801FAF081F08000F801FAF081F08000E801FAF081F08000D801FAF081F08000C", --0x20
			INIT_05             => X"801FAF081F08000C801FAF081F08000D801FAF081F08000E801FAF081F08000F", --0x28
			INIT_06             => X"801FAF081F080008801FAF081F080009801FAF081F08000A801FAF081F08000B", --0x30
			INIT_07             => X"801FAF081F080004801FAF081F080005801FAF081F080006801FAF081F080007", --0x38
			INIT_08             => X"801FAF081F080000801FAF081F080001801FAF081F080002801FAF081F080003", --0x40
			INIT_09             => X"801FAF081F080008801FAF081F080004801FAF081F080002801FAF081F080001", --0x48
			INIT_0A             => X"801FAF081F080080801FAF081F080040801FAF081F080020801FAF081F080010", --0x50
			INIT_0B             => X"801FAF081F080010801FAF081F080020801FAF081F080040801FAF081F080080", --0x58
			INIT_0C             => X"801FAF081F080001801FAF081F080002801FAF081F080004801FAF081F080008", --0x60
			INIT_0D             => X"000000000000000000000000000000000000000000000000400001081F080000", --0x68
			INIT_0E             => X"0000000082FAF0803F0800002F0100000000000082FAF0803F0800002F000000", --0x70
			INIT_0F             => X"0000000082FAF0803F0800002F0300000000000082FAF0803F0800002F020000", --0x78
			INIT_10             => X"0000000082FAF0803F0800002E0100000000000082FAF0803F0800002E000000", --0x80
			INIT_11             => X"0000000082FAF0803F0800002E0300000000000082FAF0803F0800002E020000", --0x88
			INIT_12             => X"000000000000000000000000000000000000000000000000400000981F080090", --0x90
			INIT_13             => X"180808FF180809FF18080AFF18080BFF18080CFF18080DFF18080EFF18080FFF", --0x98
			INIT_14             => X"180800FF180801FF180802FF180803FF180804FF180805FF180806FF180807FF", --0xA0
			INIT_15             => X"180806FF180805FF180804FF180803FF180802FF180801FF180800FF18080000", --0xA8
			INIT_16             => X"18080EFF18080DFF18080CFF18080BFF18080AFF180809FF180808FF180807FF", --0xB0
			INIT_17             => X"000000000000000000000000000000000000000000000000400000C01F0800B8", --0xB8
			INIT_18             => X"00000000000000000000000000000000400000C81F0800C2170800011F0800C0", --0xC0
			INIT_19             => X"00000000000000000000000000000000400000C938090000270A00001F0800C8", --0xC8
			INIT_1A             => X"0000000000000000400000D08000000F170820008000000F170810001F0800D0", --0xD0
			INIT_1B             => X"00000000400000E0820FAF08170800081F0800DB820FAF08170800011F0800D8", --0xD8
			INIT_1C             => X"00000000400000E8820FAF08170810801F0800E3820FAF08170800101F0800E0", --0xE0
			INIT_1D             => X"00000000400000F0820FAF08170808001F0800EB820FAF08170801001F0800E8", --0xE8
			INIT_1E             => X"00000000400000D8820FAF08170880001F0800F3820FAF08170810001F0800F0", --0xF0
			INIT_1F             => X"0000000000000000000000000000000000000000400000E0170810001F0800F8", --0xF8
			INIT_20             => X"0000000000000000000000000000000000000000400000E08FFFFFFF1F080100", --0x100
			INIT_21             => X"40000110820FAF083F08000021090000820FAF083F080000210800001F080108", --0x108
			INIT_22             => X"40000118820FAF083F080000210B0000820FAF083F080000210A00001F080110", --0x110
			INIT_23             => X"40000120820FAF083F080000210D0000820FAF083F080000210C00001F080118", --0x118
			INIT_24             => X"40000128820FAF083F080000210F0000820FAF083F080000210E00001F080120", --0x120
			INIT_25             => X"0000000000000000000000000000000000000000400001288FFFFFFF1F080128", --0x128
			INIT_26             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_27             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_28             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_29             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2A             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2B             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2C             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2D             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2E             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2F             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_30             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_31             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_32             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_33             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_34             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_35             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_36             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_37             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_38             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_39             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3A             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3B             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3C             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3D             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3E             => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3F             => X"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map(
			-- Port A Data: 32-bit (each) output: Port A data
			DOA    => DAT_O,            -- 32-bit output: A port data output
			--DOPA   => DOPA,             -- 4-bit output: A port parity output
			---- Port B Data: 32-bit (each) output: Port B data
			--DOB    => DOB,              -- 32-bit output: B port data output
			--DOPB   => DOPB,             -- 4-bit output: B port parity output
			-- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
			ADDRA  => adr,              -- 14-bit input: A port address input
			CLKA   => CLK_I,            -- 1-bit input: A port clock input
			ENA    => STB_I,            -- 1-bit input: A port enable input
			REGCEA => '0',              -- 1-bit input: A port register clock enable input
			RSTA   => RST_I,            -- 1-bit input: A port register set/reset input
			WEA    => we,               -- 4-bit input: Port A byte-wide write enable input
			-- Port A Data: 32-bit (each) input: Port A data
			DIA    => DAT_I,            -- 32-bit input: A port data input
			DIPA   => (others => '0'),  -- 4-bit input: A port parity input
			-- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
			ADDRB  => (others => '0'),  -- 14-bit input: B port address input
			CLKB   => '0',              -- 1-bit input: B port clock input
			ENB    => '0',              -- 1-bit input: B port enable input
			REGCEB => '0',              -- 1-bit input: B port register clock enable input
			RSTB   => '0',              -- 1-bit input: B port register set/reset input
			WEB    => (others => '0'),  -- 4-bit input: Port B byte-wide write enable input
			-- Port B Data: 32-bit (each) input: Port B data
			DIB    => (others => '0'),  -- 32-bit input: B port data input
			DIPB   => (others => '0')   -- 4-bit input: B port parity input
		);

	-- End of RAMB16BWER_inst instantiation

	adr <= ADR_I & "11111";
	we  <= WE_I & WE_I & WE_I & WE_I;
	
end Behavioral;

