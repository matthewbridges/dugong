----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:25:01 08/07/2012 
-- Design Name: 
-- Module Name:    wb_m - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity wb_m is
	generic(
		DATA_WIDTH : natural := 16;
		ADDR_WIDTH : natural := 32
	);
	port(
		--Wishbone Master Lines (inverted)
		CLK_I : out STD_LOGIC;
		RST_I : out STD_LOGIC;
		DAT_I : out STD_LOGIC_VECTOR(DATA_WIDTH - 1 downto 0);
		DAT_O : in  STD_LOGIC_VECTOR(DATA_WIDTH - 1 downto 0);
		ADR_O : in  STD_LOGIC_VECTOR(ADDR_WIDTH - 1 downto 0);
		WE_O  : in  STD_LOGIC;
		STB_O : in  STD_LOGIC;
		ACK_I : out STD_LOGIC;
		CYC_O : in  STD_LOGIC;
		--Master to WB
		WB_I  : in  STD_LOGIC_VECTOR(DATA_WIDTH downto 0);
		WB_O  : out STD_LOGIC_VECTOR(2 + ADDR_WIDTH + DATA_WIDTH downto 0)
	);
end wb_m;

architecture Behavioral of wb_m is
begin
	ACK_I <= WB_I(DATA_WIDTH);
	DAT_I <= WB_I(DATA_WIDTH - 1 downto 0);
	WB_O  <= (CYC_O & STB_O & WE_O & ADR_O & DAT_O);
end Behavioral;

