library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package sine_lut_pkg is

constant LUT_AMPL_WIDTH : natural := 16;
constant LUT_ADDR_WIDTH : natural := 15;

type lut_type is array (0 to 2 ** LUT_ADDR_WIDTH - 1) of signed(LUT_AMPL_WIDTH - 1 downto 0);
constant sine : lut_type := (
		0 => to_signed(0, LUT_AMPL_WIDTH),
		1 => to_signed(3, LUT_AMPL_WIDTH),
		2 => to_signed(6, LUT_AMPL_WIDTH),
		3 => to_signed(9, LUT_AMPL_WIDTH),
		4 => to_signed(13, LUT_AMPL_WIDTH),
		5 => to_signed(16, LUT_AMPL_WIDTH),
		6 => to_signed(19, LUT_AMPL_WIDTH),
		7 => to_signed(22, LUT_AMPL_WIDTH),
		8 => to_signed(25, LUT_AMPL_WIDTH),
		9 => to_signed(28, LUT_AMPL_WIDTH),
		10 => to_signed(31, LUT_AMPL_WIDTH),
		11 => to_signed(35, LUT_AMPL_WIDTH),
		12 => to_signed(38, LUT_AMPL_WIDTH),
		13 => to_signed(41, LUT_AMPL_WIDTH),
		14 => to_signed(44, LUT_AMPL_WIDTH),
		15 => to_signed(47, LUT_AMPL_WIDTH),
		16 => to_signed(50, LUT_AMPL_WIDTH),
		17 => to_signed(53, LUT_AMPL_WIDTH),
		18 => to_signed(57, LUT_AMPL_WIDTH),
		19 => to_signed(60, LUT_AMPL_WIDTH),
		20 => to_signed(63, LUT_AMPL_WIDTH),
		21 => to_signed(66, LUT_AMPL_WIDTH),
		22 => to_signed(69, LUT_AMPL_WIDTH),
		23 => to_signed(72, LUT_AMPL_WIDTH),
		24 => to_signed(75, LUT_AMPL_WIDTH),
		25 => to_signed(79, LUT_AMPL_WIDTH),
		26 => to_signed(82, LUT_AMPL_WIDTH),
		27 => to_signed(85, LUT_AMPL_WIDTH),
		28 => to_signed(88, LUT_AMPL_WIDTH),
		29 => to_signed(91, LUT_AMPL_WIDTH),
		30 => to_signed(94, LUT_AMPL_WIDTH),
		31 => to_signed(97, LUT_AMPL_WIDTH),
		32 => to_signed(101, LUT_AMPL_WIDTH),
		33 => to_signed(104, LUT_AMPL_WIDTH),
		34 => to_signed(107, LUT_AMPL_WIDTH),
		35 => to_signed(110, LUT_AMPL_WIDTH),
		36 => to_signed(113, LUT_AMPL_WIDTH),
		37 => to_signed(116, LUT_AMPL_WIDTH),
		38 => to_signed(119, LUT_AMPL_WIDTH),
		39 => to_signed(123, LUT_AMPL_WIDTH),
		40 => to_signed(126, LUT_AMPL_WIDTH),
		41 => to_signed(129, LUT_AMPL_WIDTH),
		42 => to_signed(132, LUT_AMPL_WIDTH),
		43 => to_signed(135, LUT_AMPL_WIDTH),
		44 => to_signed(138, LUT_AMPL_WIDTH),
		45 => to_signed(141, LUT_AMPL_WIDTH),
		46 => to_signed(145, LUT_AMPL_WIDTH),
		47 => to_signed(148, LUT_AMPL_WIDTH),
		48 => to_signed(151, LUT_AMPL_WIDTH),
		49 => to_signed(154, LUT_AMPL_WIDTH),
		50 => to_signed(157, LUT_AMPL_WIDTH),
		51 => to_signed(160, LUT_AMPL_WIDTH),
		52 => to_signed(163, LUT_AMPL_WIDTH),
		53 => to_signed(166, LUT_AMPL_WIDTH),
		54 => to_signed(170, LUT_AMPL_WIDTH),
		55 => to_signed(173, LUT_AMPL_WIDTH),
		56 => to_signed(176, LUT_AMPL_WIDTH),
		57 => to_signed(179, LUT_AMPL_WIDTH),
		58 => to_signed(182, LUT_AMPL_WIDTH),
		59 => to_signed(185, LUT_AMPL_WIDTH),
		60 => to_signed(188, LUT_AMPL_WIDTH),
		61 => to_signed(192, LUT_AMPL_WIDTH),
		62 => to_signed(195, LUT_AMPL_WIDTH),
		63 => to_signed(198, LUT_AMPL_WIDTH),
		64 => to_signed(201, LUT_AMPL_WIDTH),
		65 => to_signed(204, LUT_AMPL_WIDTH),
		66 => to_signed(207, LUT_AMPL_WIDTH),
		67 => to_signed(210, LUT_AMPL_WIDTH),
		68 => to_signed(214, LUT_AMPL_WIDTH),
		69 => to_signed(217, LUT_AMPL_WIDTH),
		70 => to_signed(220, LUT_AMPL_WIDTH),
		71 => to_signed(223, LUT_AMPL_WIDTH),
		72 => to_signed(226, LUT_AMPL_WIDTH),
		73 => to_signed(229, LUT_AMPL_WIDTH),
		74 => to_signed(232, LUT_AMPL_WIDTH),
		75 => to_signed(236, LUT_AMPL_WIDTH),
		76 => to_signed(239, LUT_AMPL_WIDTH),
		77 => to_signed(242, LUT_AMPL_WIDTH),
		78 => to_signed(245, LUT_AMPL_WIDTH),
		79 => to_signed(248, LUT_AMPL_WIDTH),
		80 => to_signed(251, LUT_AMPL_WIDTH),
		81 => to_signed(254, LUT_AMPL_WIDTH),
		82 => to_signed(258, LUT_AMPL_WIDTH),
		83 => to_signed(261, LUT_AMPL_WIDTH),
		84 => to_signed(264, LUT_AMPL_WIDTH),
		85 => to_signed(267, LUT_AMPL_WIDTH),
		86 => to_signed(270, LUT_AMPL_WIDTH),
		87 => to_signed(273, LUT_AMPL_WIDTH),
		88 => to_signed(276, LUT_AMPL_WIDTH),
		89 => to_signed(280, LUT_AMPL_WIDTH),
		90 => to_signed(283, LUT_AMPL_WIDTH),
		91 => to_signed(286, LUT_AMPL_WIDTH),
		92 => to_signed(289, LUT_AMPL_WIDTH),
		93 => to_signed(292, LUT_AMPL_WIDTH),
		94 => to_signed(295, LUT_AMPL_WIDTH),
		95 => to_signed(298, LUT_AMPL_WIDTH),
		96 => to_signed(302, LUT_AMPL_WIDTH),
		97 => to_signed(305, LUT_AMPL_WIDTH),
		98 => to_signed(308, LUT_AMPL_WIDTH),
		99 => to_signed(311, LUT_AMPL_WIDTH),
		100 => to_signed(314, LUT_AMPL_WIDTH),
		101 => to_signed(317, LUT_AMPL_WIDTH),
		102 => to_signed(320, LUT_AMPL_WIDTH),
		103 => to_signed(324, LUT_AMPL_WIDTH),
		104 => to_signed(327, LUT_AMPL_WIDTH),
		105 => to_signed(330, LUT_AMPL_WIDTH),
		106 => to_signed(333, LUT_AMPL_WIDTH),
		107 => to_signed(336, LUT_AMPL_WIDTH),
		108 => to_signed(339, LUT_AMPL_WIDTH),
		109 => to_signed(342, LUT_AMPL_WIDTH),
		110 => to_signed(346, LUT_AMPL_WIDTH),
		111 => to_signed(349, LUT_AMPL_WIDTH),
		112 => to_signed(352, LUT_AMPL_WIDTH),
		113 => to_signed(355, LUT_AMPL_WIDTH),
		114 => to_signed(358, LUT_AMPL_WIDTH),
		115 => to_signed(361, LUT_AMPL_WIDTH),
		116 => to_signed(364, LUT_AMPL_WIDTH),
		117 => to_signed(368, LUT_AMPL_WIDTH),
		118 => to_signed(371, LUT_AMPL_WIDTH),
		119 => to_signed(374, LUT_AMPL_WIDTH),
		120 => to_signed(377, LUT_AMPL_WIDTH),
		121 => to_signed(380, LUT_AMPL_WIDTH),
		122 => to_signed(383, LUT_AMPL_WIDTH),
		123 => to_signed(386, LUT_AMPL_WIDTH),
		124 => to_signed(390, LUT_AMPL_WIDTH),
		125 => to_signed(393, LUT_AMPL_WIDTH),
		126 => to_signed(396, LUT_AMPL_WIDTH),
		127 => to_signed(399, LUT_AMPL_WIDTH),
		128 => to_signed(402, LUT_AMPL_WIDTH),
		129 => to_signed(405, LUT_AMPL_WIDTH),
		130 => to_signed(408, LUT_AMPL_WIDTH),
		131 => to_signed(412, LUT_AMPL_WIDTH),
		132 => to_signed(415, LUT_AMPL_WIDTH),
		133 => to_signed(418, LUT_AMPL_WIDTH),
		134 => to_signed(421, LUT_AMPL_WIDTH),
		135 => to_signed(424, LUT_AMPL_WIDTH),
		136 => to_signed(427, LUT_AMPL_WIDTH),
		137 => to_signed(430, LUT_AMPL_WIDTH),
		138 => to_signed(434, LUT_AMPL_WIDTH),
		139 => to_signed(437, LUT_AMPL_WIDTH),
		140 => to_signed(440, LUT_AMPL_WIDTH),
		141 => to_signed(443, LUT_AMPL_WIDTH),
		142 => to_signed(446, LUT_AMPL_WIDTH),
		143 => to_signed(449, LUT_AMPL_WIDTH),
		144 => to_signed(452, LUT_AMPL_WIDTH),
		145 => to_signed(456, LUT_AMPL_WIDTH),
		146 => to_signed(459, LUT_AMPL_WIDTH),
		147 => to_signed(462, LUT_AMPL_WIDTH),
		148 => to_signed(465, LUT_AMPL_WIDTH),
		149 => to_signed(468, LUT_AMPL_WIDTH),
		150 => to_signed(471, LUT_AMPL_WIDTH),
		151 => to_signed(474, LUT_AMPL_WIDTH),
		152 => to_signed(477, LUT_AMPL_WIDTH),
		153 => to_signed(481, LUT_AMPL_WIDTH),
		154 => to_signed(484, LUT_AMPL_WIDTH),
		155 => to_signed(487, LUT_AMPL_WIDTH),
		156 => to_signed(490, LUT_AMPL_WIDTH),
		157 => to_signed(493, LUT_AMPL_WIDTH),
		158 => to_signed(496, LUT_AMPL_WIDTH),
		159 => to_signed(499, LUT_AMPL_WIDTH),
		160 => to_signed(503, LUT_AMPL_WIDTH),
		161 => to_signed(506, LUT_AMPL_WIDTH),
		162 => to_signed(509, LUT_AMPL_WIDTH),
		163 => to_signed(512, LUT_AMPL_WIDTH),
		164 => to_signed(515, LUT_AMPL_WIDTH),
		165 => to_signed(518, LUT_AMPL_WIDTH),
		166 => to_signed(521, LUT_AMPL_WIDTH),
		167 => to_signed(525, LUT_AMPL_WIDTH),
		168 => to_signed(528, LUT_AMPL_WIDTH),
		169 => to_signed(531, LUT_AMPL_WIDTH),
		170 => to_signed(534, LUT_AMPL_WIDTH),
		171 => to_signed(537, LUT_AMPL_WIDTH),
		172 => to_signed(540, LUT_AMPL_WIDTH),
		173 => to_signed(543, LUT_AMPL_WIDTH),
		174 => to_signed(547, LUT_AMPL_WIDTH),
		175 => to_signed(550, LUT_AMPL_WIDTH),
		176 => to_signed(553, LUT_AMPL_WIDTH),
		177 => to_signed(556, LUT_AMPL_WIDTH),
		178 => to_signed(559, LUT_AMPL_WIDTH),
		179 => to_signed(562, LUT_AMPL_WIDTH),
		180 => to_signed(565, LUT_AMPL_WIDTH),
		181 => to_signed(569, LUT_AMPL_WIDTH),
		182 => to_signed(572, LUT_AMPL_WIDTH),
		183 => to_signed(575, LUT_AMPL_WIDTH),
		184 => to_signed(578, LUT_AMPL_WIDTH),
		185 => to_signed(581, LUT_AMPL_WIDTH),
		186 => to_signed(584, LUT_AMPL_WIDTH),
		187 => to_signed(587, LUT_AMPL_WIDTH),
		188 => to_signed(591, LUT_AMPL_WIDTH),
		189 => to_signed(594, LUT_AMPL_WIDTH),
		190 => to_signed(597, LUT_AMPL_WIDTH),
		191 => to_signed(600, LUT_AMPL_WIDTH),
		192 => to_signed(603, LUT_AMPL_WIDTH),
		193 => to_signed(606, LUT_AMPL_WIDTH),
		194 => to_signed(609, LUT_AMPL_WIDTH),
		195 => to_signed(613, LUT_AMPL_WIDTH),
		196 => to_signed(616, LUT_AMPL_WIDTH),
		197 => to_signed(619, LUT_AMPL_WIDTH),
		198 => to_signed(622, LUT_AMPL_WIDTH),
		199 => to_signed(625, LUT_AMPL_WIDTH),
		200 => to_signed(628, LUT_AMPL_WIDTH),
		201 => to_signed(631, LUT_AMPL_WIDTH),
		202 => to_signed(635, LUT_AMPL_WIDTH),
		203 => to_signed(638, LUT_AMPL_WIDTH),
		204 => to_signed(641, LUT_AMPL_WIDTH),
		205 => to_signed(644, LUT_AMPL_WIDTH),
		206 => to_signed(647, LUT_AMPL_WIDTH),
		207 => to_signed(650, LUT_AMPL_WIDTH),
		208 => to_signed(653, LUT_AMPL_WIDTH),
		209 => to_signed(657, LUT_AMPL_WIDTH),
		210 => to_signed(660, LUT_AMPL_WIDTH),
		211 => to_signed(663, LUT_AMPL_WIDTH),
		212 => to_signed(666, LUT_AMPL_WIDTH),
		213 => to_signed(669, LUT_AMPL_WIDTH),
		214 => to_signed(672, LUT_AMPL_WIDTH),
		215 => to_signed(675, LUT_AMPL_WIDTH),
		216 => to_signed(679, LUT_AMPL_WIDTH),
		217 => to_signed(682, LUT_AMPL_WIDTH),
		218 => to_signed(685, LUT_AMPL_WIDTH),
		219 => to_signed(688, LUT_AMPL_WIDTH),
		220 => to_signed(691, LUT_AMPL_WIDTH),
		221 => to_signed(694, LUT_AMPL_WIDTH),
		222 => to_signed(697, LUT_AMPL_WIDTH),
		223 => to_signed(701, LUT_AMPL_WIDTH),
		224 => to_signed(704, LUT_AMPL_WIDTH),
		225 => to_signed(707, LUT_AMPL_WIDTH),
		226 => to_signed(710, LUT_AMPL_WIDTH),
		227 => to_signed(713, LUT_AMPL_WIDTH),
		228 => to_signed(716, LUT_AMPL_WIDTH),
		229 => to_signed(719, LUT_AMPL_WIDTH),
		230 => to_signed(722, LUT_AMPL_WIDTH),
		231 => to_signed(726, LUT_AMPL_WIDTH),
		232 => to_signed(729, LUT_AMPL_WIDTH),
		233 => to_signed(732, LUT_AMPL_WIDTH),
		234 => to_signed(735, LUT_AMPL_WIDTH),
		235 => to_signed(738, LUT_AMPL_WIDTH),
		236 => to_signed(741, LUT_AMPL_WIDTH),
		237 => to_signed(744, LUT_AMPL_WIDTH),
		238 => to_signed(748, LUT_AMPL_WIDTH),
		239 => to_signed(751, LUT_AMPL_WIDTH),
		240 => to_signed(754, LUT_AMPL_WIDTH),
		241 => to_signed(757, LUT_AMPL_WIDTH),
		242 => to_signed(760, LUT_AMPL_WIDTH),
		243 => to_signed(763, LUT_AMPL_WIDTH),
		244 => to_signed(766, LUT_AMPL_WIDTH),
		245 => to_signed(770, LUT_AMPL_WIDTH),
		246 => to_signed(773, LUT_AMPL_WIDTH),
		247 => to_signed(776, LUT_AMPL_WIDTH),
		248 => to_signed(779, LUT_AMPL_WIDTH),
		249 => to_signed(782, LUT_AMPL_WIDTH),
		250 => to_signed(785, LUT_AMPL_WIDTH),
		251 => to_signed(788, LUT_AMPL_WIDTH),
		252 => to_signed(792, LUT_AMPL_WIDTH),
		253 => to_signed(795, LUT_AMPL_WIDTH),
		254 => to_signed(798, LUT_AMPL_WIDTH),
		255 => to_signed(801, LUT_AMPL_WIDTH),
		256 => to_signed(804, LUT_AMPL_WIDTH),
		257 => to_signed(807, LUT_AMPL_WIDTH),
		258 => to_signed(810, LUT_AMPL_WIDTH),
		259 => to_signed(814, LUT_AMPL_WIDTH),
		260 => to_signed(817, LUT_AMPL_WIDTH),
		261 => to_signed(820, LUT_AMPL_WIDTH),
		262 => to_signed(823, LUT_AMPL_WIDTH),
		263 => to_signed(826, LUT_AMPL_WIDTH),
		264 => to_signed(829, LUT_AMPL_WIDTH),
		265 => to_signed(832, LUT_AMPL_WIDTH),
		266 => to_signed(836, LUT_AMPL_WIDTH),
		267 => to_signed(839, LUT_AMPL_WIDTH),
		268 => to_signed(842, LUT_AMPL_WIDTH),
		269 => to_signed(845, LUT_AMPL_WIDTH),
		270 => to_signed(848, LUT_AMPL_WIDTH),
		271 => to_signed(851, LUT_AMPL_WIDTH),
		272 => to_signed(854, LUT_AMPL_WIDTH),
		273 => to_signed(858, LUT_AMPL_WIDTH),
		274 => to_signed(861, LUT_AMPL_WIDTH),
		275 => to_signed(864, LUT_AMPL_WIDTH),
		276 => to_signed(867, LUT_AMPL_WIDTH),
		277 => to_signed(870, LUT_AMPL_WIDTH),
		278 => to_signed(873, LUT_AMPL_WIDTH),
		279 => to_signed(876, LUT_AMPL_WIDTH),
		280 => to_signed(880, LUT_AMPL_WIDTH),
		281 => to_signed(883, LUT_AMPL_WIDTH),
		282 => to_signed(886, LUT_AMPL_WIDTH),
		283 => to_signed(889, LUT_AMPL_WIDTH),
		284 => to_signed(892, LUT_AMPL_WIDTH),
		285 => to_signed(895, LUT_AMPL_WIDTH),
		286 => to_signed(898, LUT_AMPL_WIDTH),
		287 => to_signed(901, LUT_AMPL_WIDTH),
		288 => to_signed(905, LUT_AMPL_WIDTH),
		289 => to_signed(908, LUT_AMPL_WIDTH),
		290 => to_signed(911, LUT_AMPL_WIDTH),
		291 => to_signed(914, LUT_AMPL_WIDTH),
		292 => to_signed(917, LUT_AMPL_WIDTH),
		293 => to_signed(920, LUT_AMPL_WIDTH),
		294 => to_signed(923, LUT_AMPL_WIDTH),
		295 => to_signed(927, LUT_AMPL_WIDTH),
		296 => to_signed(930, LUT_AMPL_WIDTH),
		297 => to_signed(933, LUT_AMPL_WIDTH),
		298 => to_signed(936, LUT_AMPL_WIDTH),
		299 => to_signed(939, LUT_AMPL_WIDTH),
		300 => to_signed(942, LUT_AMPL_WIDTH),
		301 => to_signed(945, LUT_AMPL_WIDTH),
		302 => to_signed(949, LUT_AMPL_WIDTH),
		303 => to_signed(952, LUT_AMPL_WIDTH),
		304 => to_signed(955, LUT_AMPL_WIDTH),
		305 => to_signed(958, LUT_AMPL_WIDTH),
		306 => to_signed(961, LUT_AMPL_WIDTH),
		307 => to_signed(964, LUT_AMPL_WIDTH),
		308 => to_signed(967, LUT_AMPL_WIDTH),
		309 => to_signed(971, LUT_AMPL_WIDTH),
		310 => to_signed(974, LUT_AMPL_WIDTH),
		311 => to_signed(977, LUT_AMPL_WIDTH),
		312 => to_signed(980, LUT_AMPL_WIDTH),
		313 => to_signed(983, LUT_AMPL_WIDTH),
		314 => to_signed(986, LUT_AMPL_WIDTH),
		315 => to_signed(989, LUT_AMPL_WIDTH),
		316 => to_signed(993, LUT_AMPL_WIDTH),
		317 => to_signed(996, LUT_AMPL_WIDTH),
		318 => to_signed(999, LUT_AMPL_WIDTH),
		319 => to_signed(1002, LUT_AMPL_WIDTH),
		320 => to_signed(1005, LUT_AMPL_WIDTH),
		321 => to_signed(1008, LUT_AMPL_WIDTH),
		322 => to_signed(1011, LUT_AMPL_WIDTH),
		323 => to_signed(1015, LUT_AMPL_WIDTH),
		324 => to_signed(1018, LUT_AMPL_WIDTH),
		325 => to_signed(1021, LUT_AMPL_WIDTH),
		326 => to_signed(1024, LUT_AMPL_WIDTH),
		327 => to_signed(1027, LUT_AMPL_WIDTH),
		328 => to_signed(1030, LUT_AMPL_WIDTH),
		329 => to_signed(1033, LUT_AMPL_WIDTH),
		330 => to_signed(1037, LUT_AMPL_WIDTH),
		331 => to_signed(1040, LUT_AMPL_WIDTH),
		332 => to_signed(1043, LUT_AMPL_WIDTH),
		333 => to_signed(1046, LUT_AMPL_WIDTH),
		334 => to_signed(1049, LUT_AMPL_WIDTH),
		335 => to_signed(1052, LUT_AMPL_WIDTH),
		336 => to_signed(1055, LUT_AMPL_WIDTH),
		337 => to_signed(1059, LUT_AMPL_WIDTH),
		338 => to_signed(1062, LUT_AMPL_WIDTH),
		339 => to_signed(1065, LUT_AMPL_WIDTH),
		340 => to_signed(1068, LUT_AMPL_WIDTH),
		341 => to_signed(1071, LUT_AMPL_WIDTH),
		342 => to_signed(1074, LUT_AMPL_WIDTH),
		343 => to_signed(1077, LUT_AMPL_WIDTH),
		344 => to_signed(1080, LUT_AMPL_WIDTH),
		345 => to_signed(1084, LUT_AMPL_WIDTH),
		346 => to_signed(1087, LUT_AMPL_WIDTH),
		347 => to_signed(1090, LUT_AMPL_WIDTH),
		348 => to_signed(1093, LUT_AMPL_WIDTH),
		349 => to_signed(1096, LUT_AMPL_WIDTH),
		350 => to_signed(1099, LUT_AMPL_WIDTH),
		351 => to_signed(1102, LUT_AMPL_WIDTH),
		352 => to_signed(1106, LUT_AMPL_WIDTH),
		353 => to_signed(1109, LUT_AMPL_WIDTH),
		354 => to_signed(1112, LUT_AMPL_WIDTH),
		355 => to_signed(1115, LUT_AMPL_WIDTH),
		356 => to_signed(1118, LUT_AMPL_WIDTH),
		357 => to_signed(1121, LUT_AMPL_WIDTH),
		358 => to_signed(1124, LUT_AMPL_WIDTH),
		359 => to_signed(1128, LUT_AMPL_WIDTH),
		360 => to_signed(1131, LUT_AMPL_WIDTH),
		361 => to_signed(1134, LUT_AMPL_WIDTH),
		362 => to_signed(1137, LUT_AMPL_WIDTH),
		363 => to_signed(1140, LUT_AMPL_WIDTH),
		364 => to_signed(1143, LUT_AMPL_WIDTH),
		365 => to_signed(1146, LUT_AMPL_WIDTH),
		366 => to_signed(1150, LUT_AMPL_WIDTH),
		367 => to_signed(1153, LUT_AMPL_WIDTH),
		368 => to_signed(1156, LUT_AMPL_WIDTH),
		369 => to_signed(1159, LUT_AMPL_WIDTH),
		370 => to_signed(1162, LUT_AMPL_WIDTH),
		371 => to_signed(1165, LUT_AMPL_WIDTH),
		372 => to_signed(1168, LUT_AMPL_WIDTH),
		373 => to_signed(1172, LUT_AMPL_WIDTH),
		374 => to_signed(1175, LUT_AMPL_WIDTH),
		375 => to_signed(1178, LUT_AMPL_WIDTH),
		376 => to_signed(1181, LUT_AMPL_WIDTH),
		377 => to_signed(1184, LUT_AMPL_WIDTH),
		378 => to_signed(1187, LUT_AMPL_WIDTH),
		379 => to_signed(1190, LUT_AMPL_WIDTH),
		380 => to_signed(1194, LUT_AMPL_WIDTH),
		381 => to_signed(1197, LUT_AMPL_WIDTH),
		382 => to_signed(1200, LUT_AMPL_WIDTH),
		383 => to_signed(1203, LUT_AMPL_WIDTH),
		384 => to_signed(1206, LUT_AMPL_WIDTH),
		385 => to_signed(1209, LUT_AMPL_WIDTH),
		386 => to_signed(1212, LUT_AMPL_WIDTH),
		387 => to_signed(1215, LUT_AMPL_WIDTH),
		388 => to_signed(1219, LUT_AMPL_WIDTH),
		389 => to_signed(1222, LUT_AMPL_WIDTH),
		390 => to_signed(1225, LUT_AMPL_WIDTH),
		391 => to_signed(1228, LUT_AMPL_WIDTH),
		392 => to_signed(1231, LUT_AMPL_WIDTH),
		393 => to_signed(1234, LUT_AMPL_WIDTH),
		394 => to_signed(1237, LUT_AMPL_WIDTH),
		395 => to_signed(1241, LUT_AMPL_WIDTH),
		396 => to_signed(1244, LUT_AMPL_WIDTH),
		397 => to_signed(1247, LUT_AMPL_WIDTH),
		398 => to_signed(1250, LUT_AMPL_WIDTH),
		399 => to_signed(1253, LUT_AMPL_WIDTH),
		400 => to_signed(1256, LUT_AMPL_WIDTH),
		401 => to_signed(1259, LUT_AMPL_WIDTH),
		402 => to_signed(1263, LUT_AMPL_WIDTH),
		403 => to_signed(1266, LUT_AMPL_WIDTH),
		404 => to_signed(1269, LUT_AMPL_WIDTH),
		405 => to_signed(1272, LUT_AMPL_WIDTH),
		406 => to_signed(1275, LUT_AMPL_WIDTH),
		407 => to_signed(1278, LUT_AMPL_WIDTH),
		408 => to_signed(1281, LUT_AMPL_WIDTH),
		409 => to_signed(1285, LUT_AMPL_WIDTH),
		410 => to_signed(1288, LUT_AMPL_WIDTH),
		411 => to_signed(1291, LUT_AMPL_WIDTH),
		412 => to_signed(1294, LUT_AMPL_WIDTH),
		413 => to_signed(1297, LUT_AMPL_WIDTH),
		414 => to_signed(1300, LUT_AMPL_WIDTH),
		415 => to_signed(1303, LUT_AMPL_WIDTH),
		416 => to_signed(1307, LUT_AMPL_WIDTH),
		417 => to_signed(1310, LUT_AMPL_WIDTH),
		418 => to_signed(1313, LUT_AMPL_WIDTH),
		419 => to_signed(1316, LUT_AMPL_WIDTH),
		420 => to_signed(1319, LUT_AMPL_WIDTH),
		421 => to_signed(1322, LUT_AMPL_WIDTH),
		422 => to_signed(1325, LUT_AMPL_WIDTH),
		423 => to_signed(1328, LUT_AMPL_WIDTH),
		424 => to_signed(1332, LUT_AMPL_WIDTH),
		425 => to_signed(1335, LUT_AMPL_WIDTH),
		426 => to_signed(1338, LUT_AMPL_WIDTH),
		427 => to_signed(1341, LUT_AMPL_WIDTH),
		428 => to_signed(1344, LUT_AMPL_WIDTH),
		429 => to_signed(1347, LUT_AMPL_WIDTH),
		430 => to_signed(1350, LUT_AMPL_WIDTH),
		431 => to_signed(1354, LUT_AMPL_WIDTH),
		432 => to_signed(1357, LUT_AMPL_WIDTH),
		433 => to_signed(1360, LUT_AMPL_WIDTH),
		434 => to_signed(1363, LUT_AMPL_WIDTH),
		435 => to_signed(1366, LUT_AMPL_WIDTH),
		436 => to_signed(1369, LUT_AMPL_WIDTH),
		437 => to_signed(1372, LUT_AMPL_WIDTH),
		438 => to_signed(1376, LUT_AMPL_WIDTH),
		439 => to_signed(1379, LUT_AMPL_WIDTH),
		440 => to_signed(1382, LUT_AMPL_WIDTH),
		441 => to_signed(1385, LUT_AMPL_WIDTH),
		442 => to_signed(1388, LUT_AMPL_WIDTH),
		443 => to_signed(1391, LUT_AMPL_WIDTH),
		444 => to_signed(1394, LUT_AMPL_WIDTH),
		445 => to_signed(1398, LUT_AMPL_WIDTH),
		446 => to_signed(1401, LUT_AMPL_WIDTH),
		447 => to_signed(1404, LUT_AMPL_WIDTH),
		448 => to_signed(1407, LUT_AMPL_WIDTH),
		449 => to_signed(1410, LUT_AMPL_WIDTH),
		450 => to_signed(1413, LUT_AMPL_WIDTH),
		451 => to_signed(1416, LUT_AMPL_WIDTH),
		452 => to_signed(1420, LUT_AMPL_WIDTH),
		453 => to_signed(1423, LUT_AMPL_WIDTH),
		454 => to_signed(1426, LUT_AMPL_WIDTH),
		455 => to_signed(1429, LUT_AMPL_WIDTH),
		456 => to_signed(1432, LUT_AMPL_WIDTH),
		457 => to_signed(1435, LUT_AMPL_WIDTH),
		458 => to_signed(1438, LUT_AMPL_WIDTH),
		459 => to_signed(1441, LUT_AMPL_WIDTH),
		460 => to_signed(1445, LUT_AMPL_WIDTH),
		461 => to_signed(1448, LUT_AMPL_WIDTH),
		462 => to_signed(1451, LUT_AMPL_WIDTH),
		463 => to_signed(1454, LUT_AMPL_WIDTH),
		464 => to_signed(1457, LUT_AMPL_WIDTH),
		465 => to_signed(1460, LUT_AMPL_WIDTH),
		466 => to_signed(1463, LUT_AMPL_WIDTH),
		467 => to_signed(1467, LUT_AMPL_WIDTH),
		468 => to_signed(1470, LUT_AMPL_WIDTH),
		469 => to_signed(1473, LUT_AMPL_WIDTH),
		470 => to_signed(1476, LUT_AMPL_WIDTH),
		471 => to_signed(1479, LUT_AMPL_WIDTH),
		472 => to_signed(1482, LUT_AMPL_WIDTH),
		473 => to_signed(1485, LUT_AMPL_WIDTH),
		474 => to_signed(1489, LUT_AMPL_WIDTH),
		475 => to_signed(1492, LUT_AMPL_WIDTH),
		476 => to_signed(1495, LUT_AMPL_WIDTH),
		477 => to_signed(1498, LUT_AMPL_WIDTH),
		478 => to_signed(1501, LUT_AMPL_WIDTH),
		479 => to_signed(1504, LUT_AMPL_WIDTH),
		480 => to_signed(1507, LUT_AMPL_WIDTH),
		481 => to_signed(1511, LUT_AMPL_WIDTH),
		482 => to_signed(1514, LUT_AMPL_WIDTH),
		483 => to_signed(1517, LUT_AMPL_WIDTH),
		484 => to_signed(1520, LUT_AMPL_WIDTH),
		485 => to_signed(1523, LUT_AMPL_WIDTH),
		486 => to_signed(1526, LUT_AMPL_WIDTH),
		487 => to_signed(1529, LUT_AMPL_WIDTH),
		488 => to_signed(1532, LUT_AMPL_WIDTH),
		489 => to_signed(1536, LUT_AMPL_WIDTH),
		490 => to_signed(1539, LUT_AMPL_WIDTH),
		491 => to_signed(1542, LUT_AMPL_WIDTH),
		492 => to_signed(1545, LUT_AMPL_WIDTH),
		493 => to_signed(1548, LUT_AMPL_WIDTH),
		494 => to_signed(1551, LUT_AMPL_WIDTH),
		495 => to_signed(1554, LUT_AMPL_WIDTH),
		496 => to_signed(1558, LUT_AMPL_WIDTH),
		497 => to_signed(1561, LUT_AMPL_WIDTH),
		498 => to_signed(1564, LUT_AMPL_WIDTH),
		499 => to_signed(1567, LUT_AMPL_WIDTH),
		500 => to_signed(1570, LUT_AMPL_WIDTH),
		501 => to_signed(1573, LUT_AMPL_WIDTH),
		502 => to_signed(1576, LUT_AMPL_WIDTH),
		503 => to_signed(1580, LUT_AMPL_WIDTH),
		504 => to_signed(1583, LUT_AMPL_WIDTH),
		505 => to_signed(1586, LUT_AMPL_WIDTH),
		506 => to_signed(1589, LUT_AMPL_WIDTH),
		507 => to_signed(1592, LUT_AMPL_WIDTH),
		508 => to_signed(1595, LUT_AMPL_WIDTH),
		509 => to_signed(1598, LUT_AMPL_WIDTH),
		510 => to_signed(1602, LUT_AMPL_WIDTH),
		511 => to_signed(1605, LUT_AMPL_WIDTH),
		512 => to_signed(1608, LUT_AMPL_WIDTH),
		513 => to_signed(1611, LUT_AMPL_WIDTH),
		514 => to_signed(1614, LUT_AMPL_WIDTH),
		515 => to_signed(1617, LUT_AMPL_WIDTH),
		516 => to_signed(1620, LUT_AMPL_WIDTH),
		517 => to_signed(1623, LUT_AMPL_WIDTH),
		518 => to_signed(1627, LUT_AMPL_WIDTH),
		519 => to_signed(1630, LUT_AMPL_WIDTH),
		520 => to_signed(1633, LUT_AMPL_WIDTH),
		521 => to_signed(1636, LUT_AMPL_WIDTH),
		522 => to_signed(1639, LUT_AMPL_WIDTH),
		523 => to_signed(1642, LUT_AMPL_WIDTH),
		524 => to_signed(1645, LUT_AMPL_WIDTH),
		525 => to_signed(1649, LUT_AMPL_WIDTH),
		526 => to_signed(1652, LUT_AMPL_WIDTH),
		527 => to_signed(1655, LUT_AMPL_WIDTH),
		528 => to_signed(1658, LUT_AMPL_WIDTH),
		529 => to_signed(1661, LUT_AMPL_WIDTH),
		530 => to_signed(1664, LUT_AMPL_WIDTH),
		531 => to_signed(1667, LUT_AMPL_WIDTH),
		532 => to_signed(1671, LUT_AMPL_WIDTH),
		533 => to_signed(1674, LUT_AMPL_WIDTH),
		534 => to_signed(1677, LUT_AMPL_WIDTH),
		535 => to_signed(1680, LUT_AMPL_WIDTH),
		536 => to_signed(1683, LUT_AMPL_WIDTH),
		537 => to_signed(1686, LUT_AMPL_WIDTH),
		538 => to_signed(1689, LUT_AMPL_WIDTH),
		539 => to_signed(1693, LUT_AMPL_WIDTH),
		540 => to_signed(1696, LUT_AMPL_WIDTH),
		541 => to_signed(1699, LUT_AMPL_WIDTH),
		542 => to_signed(1702, LUT_AMPL_WIDTH),
		543 => to_signed(1705, LUT_AMPL_WIDTH),
		544 => to_signed(1708, LUT_AMPL_WIDTH),
		545 => to_signed(1711, LUT_AMPL_WIDTH),
		546 => to_signed(1714, LUT_AMPL_WIDTH),
		547 => to_signed(1718, LUT_AMPL_WIDTH),
		548 => to_signed(1721, LUT_AMPL_WIDTH),
		549 => to_signed(1724, LUT_AMPL_WIDTH),
		550 => to_signed(1727, LUT_AMPL_WIDTH),
		551 => to_signed(1730, LUT_AMPL_WIDTH),
		552 => to_signed(1733, LUT_AMPL_WIDTH),
		553 => to_signed(1736, LUT_AMPL_WIDTH),
		554 => to_signed(1740, LUT_AMPL_WIDTH),
		555 => to_signed(1743, LUT_AMPL_WIDTH),
		556 => to_signed(1746, LUT_AMPL_WIDTH),
		557 => to_signed(1749, LUT_AMPL_WIDTH),
		558 => to_signed(1752, LUT_AMPL_WIDTH),
		559 => to_signed(1755, LUT_AMPL_WIDTH),
		560 => to_signed(1758, LUT_AMPL_WIDTH),
		561 => to_signed(1762, LUT_AMPL_WIDTH),
		562 => to_signed(1765, LUT_AMPL_WIDTH),
		563 => to_signed(1768, LUT_AMPL_WIDTH),
		564 => to_signed(1771, LUT_AMPL_WIDTH),
		565 => to_signed(1774, LUT_AMPL_WIDTH),
		566 => to_signed(1777, LUT_AMPL_WIDTH),
		567 => to_signed(1780, LUT_AMPL_WIDTH),
		568 => to_signed(1783, LUT_AMPL_WIDTH),
		569 => to_signed(1787, LUT_AMPL_WIDTH),
		570 => to_signed(1790, LUT_AMPL_WIDTH),
		571 => to_signed(1793, LUT_AMPL_WIDTH),
		572 => to_signed(1796, LUT_AMPL_WIDTH),
		573 => to_signed(1799, LUT_AMPL_WIDTH),
		574 => to_signed(1802, LUT_AMPL_WIDTH),
		575 => to_signed(1805, LUT_AMPL_WIDTH),
		576 => to_signed(1809, LUT_AMPL_WIDTH),
		577 => to_signed(1812, LUT_AMPL_WIDTH),
		578 => to_signed(1815, LUT_AMPL_WIDTH),
		579 => to_signed(1818, LUT_AMPL_WIDTH),
		580 => to_signed(1821, LUT_AMPL_WIDTH),
		581 => to_signed(1824, LUT_AMPL_WIDTH),
		582 => to_signed(1827, LUT_AMPL_WIDTH),
		583 => to_signed(1831, LUT_AMPL_WIDTH),
		584 => to_signed(1834, LUT_AMPL_WIDTH),
		585 => to_signed(1837, LUT_AMPL_WIDTH),
		586 => to_signed(1840, LUT_AMPL_WIDTH),
		587 => to_signed(1843, LUT_AMPL_WIDTH),
		588 => to_signed(1846, LUT_AMPL_WIDTH),
		589 => to_signed(1849, LUT_AMPL_WIDTH),
		590 => to_signed(1852, LUT_AMPL_WIDTH),
		591 => to_signed(1856, LUT_AMPL_WIDTH),
		592 => to_signed(1859, LUT_AMPL_WIDTH),
		593 => to_signed(1862, LUT_AMPL_WIDTH),
		594 => to_signed(1865, LUT_AMPL_WIDTH),
		595 => to_signed(1868, LUT_AMPL_WIDTH),
		596 => to_signed(1871, LUT_AMPL_WIDTH),
		597 => to_signed(1874, LUT_AMPL_WIDTH),
		598 => to_signed(1878, LUT_AMPL_WIDTH),
		599 => to_signed(1881, LUT_AMPL_WIDTH),
		600 => to_signed(1884, LUT_AMPL_WIDTH),
		601 => to_signed(1887, LUT_AMPL_WIDTH),
		602 => to_signed(1890, LUT_AMPL_WIDTH),
		603 => to_signed(1893, LUT_AMPL_WIDTH),
		604 => to_signed(1896, LUT_AMPL_WIDTH),
		605 => to_signed(1900, LUT_AMPL_WIDTH),
		606 => to_signed(1903, LUT_AMPL_WIDTH),
		607 => to_signed(1906, LUT_AMPL_WIDTH),
		608 => to_signed(1909, LUT_AMPL_WIDTH),
		609 => to_signed(1912, LUT_AMPL_WIDTH),
		610 => to_signed(1915, LUT_AMPL_WIDTH),
		611 => to_signed(1918, LUT_AMPL_WIDTH),
		612 => to_signed(1921, LUT_AMPL_WIDTH),
		613 => to_signed(1925, LUT_AMPL_WIDTH),
		614 => to_signed(1928, LUT_AMPL_WIDTH),
		615 => to_signed(1931, LUT_AMPL_WIDTH),
		616 => to_signed(1934, LUT_AMPL_WIDTH),
		617 => to_signed(1937, LUT_AMPL_WIDTH),
		618 => to_signed(1940, LUT_AMPL_WIDTH),
		619 => to_signed(1943, LUT_AMPL_WIDTH),
		620 => to_signed(1947, LUT_AMPL_WIDTH),
		621 => to_signed(1950, LUT_AMPL_WIDTH),
		622 => to_signed(1953, LUT_AMPL_WIDTH),
		623 => to_signed(1956, LUT_AMPL_WIDTH),
		624 => to_signed(1959, LUT_AMPL_WIDTH),
		625 => to_signed(1962, LUT_AMPL_WIDTH),
		626 => to_signed(1965, LUT_AMPL_WIDTH),
		627 => to_signed(1969, LUT_AMPL_WIDTH),
		628 => to_signed(1972, LUT_AMPL_WIDTH),
		629 => to_signed(1975, LUT_AMPL_WIDTH),
		630 => to_signed(1978, LUT_AMPL_WIDTH),
		631 => to_signed(1981, LUT_AMPL_WIDTH),
		632 => to_signed(1984, LUT_AMPL_WIDTH),
		633 => to_signed(1987, LUT_AMPL_WIDTH),
		634 => to_signed(1990, LUT_AMPL_WIDTH),
		635 => to_signed(1994, LUT_AMPL_WIDTH),
		636 => to_signed(1997, LUT_AMPL_WIDTH),
		637 => to_signed(2000, LUT_AMPL_WIDTH),
		638 => to_signed(2003, LUT_AMPL_WIDTH),
		639 => to_signed(2006, LUT_AMPL_WIDTH),
		640 => to_signed(2009, LUT_AMPL_WIDTH),
		641 => to_signed(2012, LUT_AMPL_WIDTH),
		642 => to_signed(2016, LUT_AMPL_WIDTH),
		643 => to_signed(2019, LUT_AMPL_WIDTH),
		644 => to_signed(2022, LUT_AMPL_WIDTH),
		645 => to_signed(2025, LUT_AMPL_WIDTH),
		646 => to_signed(2028, LUT_AMPL_WIDTH),
		647 => to_signed(2031, LUT_AMPL_WIDTH),
		648 => to_signed(2034, LUT_AMPL_WIDTH),
		649 => to_signed(2038, LUT_AMPL_WIDTH),
		650 => to_signed(2041, LUT_AMPL_WIDTH),
		651 => to_signed(2044, LUT_AMPL_WIDTH),
		652 => to_signed(2047, LUT_AMPL_WIDTH),
		653 => to_signed(2050, LUT_AMPL_WIDTH),
		654 => to_signed(2053, LUT_AMPL_WIDTH),
		655 => to_signed(2056, LUT_AMPL_WIDTH),
		656 => to_signed(2059, LUT_AMPL_WIDTH),
		657 => to_signed(2063, LUT_AMPL_WIDTH),
		658 => to_signed(2066, LUT_AMPL_WIDTH),
		659 => to_signed(2069, LUT_AMPL_WIDTH),
		660 => to_signed(2072, LUT_AMPL_WIDTH),
		661 => to_signed(2075, LUT_AMPL_WIDTH),
		662 => to_signed(2078, LUT_AMPL_WIDTH),
		663 => to_signed(2081, LUT_AMPL_WIDTH),
		664 => to_signed(2085, LUT_AMPL_WIDTH),
		665 => to_signed(2088, LUT_AMPL_WIDTH),
		666 => to_signed(2091, LUT_AMPL_WIDTH),
		667 => to_signed(2094, LUT_AMPL_WIDTH),
		668 => to_signed(2097, LUT_AMPL_WIDTH),
		669 => to_signed(2100, LUT_AMPL_WIDTH),
		670 => to_signed(2103, LUT_AMPL_WIDTH),
		671 => to_signed(2106, LUT_AMPL_WIDTH),
		672 => to_signed(2110, LUT_AMPL_WIDTH),
		673 => to_signed(2113, LUT_AMPL_WIDTH),
		674 => to_signed(2116, LUT_AMPL_WIDTH),
		675 => to_signed(2119, LUT_AMPL_WIDTH),
		676 => to_signed(2122, LUT_AMPL_WIDTH),
		677 => to_signed(2125, LUT_AMPL_WIDTH),
		678 => to_signed(2128, LUT_AMPL_WIDTH),
		679 => to_signed(2132, LUT_AMPL_WIDTH),
		680 => to_signed(2135, LUT_AMPL_WIDTH),
		681 => to_signed(2138, LUT_AMPL_WIDTH),
		682 => to_signed(2141, LUT_AMPL_WIDTH),
		683 => to_signed(2144, LUT_AMPL_WIDTH),
		684 => to_signed(2147, LUT_AMPL_WIDTH),
		685 => to_signed(2150, LUT_AMPL_WIDTH),
		686 => to_signed(2154, LUT_AMPL_WIDTH),
		687 => to_signed(2157, LUT_AMPL_WIDTH),
		688 => to_signed(2160, LUT_AMPL_WIDTH),
		689 => to_signed(2163, LUT_AMPL_WIDTH),
		690 => to_signed(2166, LUT_AMPL_WIDTH),
		691 => to_signed(2169, LUT_AMPL_WIDTH),
		692 => to_signed(2172, LUT_AMPL_WIDTH),
		693 => to_signed(2175, LUT_AMPL_WIDTH),
		694 => to_signed(2179, LUT_AMPL_WIDTH),
		695 => to_signed(2182, LUT_AMPL_WIDTH),
		696 => to_signed(2185, LUT_AMPL_WIDTH),
		697 => to_signed(2188, LUT_AMPL_WIDTH),
		698 => to_signed(2191, LUT_AMPL_WIDTH),
		699 => to_signed(2194, LUT_AMPL_WIDTH),
		700 => to_signed(2197, LUT_AMPL_WIDTH),
		701 => to_signed(2201, LUT_AMPL_WIDTH),
		702 => to_signed(2204, LUT_AMPL_WIDTH),
		703 => to_signed(2207, LUT_AMPL_WIDTH),
		704 => to_signed(2210, LUT_AMPL_WIDTH),
		705 => to_signed(2213, LUT_AMPL_WIDTH),
		706 => to_signed(2216, LUT_AMPL_WIDTH),
		707 => to_signed(2219, LUT_AMPL_WIDTH),
		708 => to_signed(2222, LUT_AMPL_WIDTH),
		709 => to_signed(2226, LUT_AMPL_WIDTH),
		710 => to_signed(2229, LUT_AMPL_WIDTH),
		711 => to_signed(2232, LUT_AMPL_WIDTH),
		712 => to_signed(2235, LUT_AMPL_WIDTH),
		713 => to_signed(2238, LUT_AMPL_WIDTH),
		714 => to_signed(2241, LUT_AMPL_WIDTH),
		715 => to_signed(2244, LUT_AMPL_WIDTH),
		716 => to_signed(2248, LUT_AMPL_WIDTH),
		717 => to_signed(2251, LUT_AMPL_WIDTH),
		718 => to_signed(2254, LUT_AMPL_WIDTH),
		719 => to_signed(2257, LUT_AMPL_WIDTH),
		720 => to_signed(2260, LUT_AMPL_WIDTH),
		721 => to_signed(2263, LUT_AMPL_WIDTH),
		722 => to_signed(2266, LUT_AMPL_WIDTH),
		723 => to_signed(2269, LUT_AMPL_WIDTH),
		724 => to_signed(2273, LUT_AMPL_WIDTH),
		725 => to_signed(2276, LUT_AMPL_WIDTH),
		726 => to_signed(2279, LUT_AMPL_WIDTH),
		727 => to_signed(2282, LUT_AMPL_WIDTH),
		728 => to_signed(2285, LUT_AMPL_WIDTH),
		729 => to_signed(2288, LUT_AMPL_WIDTH),
		730 => to_signed(2291, LUT_AMPL_WIDTH),
		731 => to_signed(2295, LUT_AMPL_WIDTH),
		732 => to_signed(2298, LUT_AMPL_WIDTH),
		733 => to_signed(2301, LUT_AMPL_WIDTH),
		734 => to_signed(2304, LUT_AMPL_WIDTH),
		735 => to_signed(2307, LUT_AMPL_WIDTH),
		736 => to_signed(2310, LUT_AMPL_WIDTH),
		737 => to_signed(2313, LUT_AMPL_WIDTH),
		738 => to_signed(2316, LUT_AMPL_WIDTH),
		739 => to_signed(2320, LUT_AMPL_WIDTH),
		740 => to_signed(2323, LUT_AMPL_WIDTH),
		741 => to_signed(2326, LUT_AMPL_WIDTH),
		742 => to_signed(2329, LUT_AMPL_WIDTH),
		743 => to_signed(2332, LUT_AMPL_WIDTH),
		744 => to_signed(2335, LUT_AMPL_WIDTH),
		745 => to_signed(2338, LUT_AMPL_WIDTH),
		746 => to_signed(2342, LUT_AMPL_WIDTH),
		747 => to_signed(2345, LUT_AMPL_WIDTH),
		748 => to_signed(2348, LUT_AMPL_WIDTH),
		749 => to_signed(2351, LUT_AMPL_WIDTH),
		750 => to_signed(2354, LUT_AMPL_WIDTH),
		751 => to_signed(2357, LUT_AMPL_WIDTH),
		752 => to_signed(2360, LUT_AMPL_WIDTH),
		753 => to_signed(2363, LUT_AMPL_WIDTH),
		754 => to_signed(2367, LUT_AMPL_WIDTH),
		755 => to_signed(2370, LUT_AMPL_WIDTH),
		756 => to_signed(2373, LUT_AMPL_WIDTH),
		757 => to_signed(2376, LUT_AMPL_WIDTH),
		758 => to_signed(2379, LUT_AMPL_WIDTH),
		759 => to_signed(2382, LUT_AMPL_WIDTH),
		760 => to_signed(2385, LUT_AMPL_WIDTH),
		761 => to_signed(2389, LUT_AMPL_WIDTH),
		762 => to_signed(2392, LUT_AMPL_WIDTH),
		763 => to_signed(2395, LUT_AMPL_WIDTH),
		764 => to_signed(2398, LUT_AMPL_WIDTH),
		765 => to_signed(2401, LUT_AMPL_WIDTH),
		766 => to_signed(2404, LUT_AMPL_WIDTH),
		767 => to_signed(2407, LUT_AMPL_WIDTH),
		768 => to_signed(2410, LUT_AMPL_WIDTH),
		769 => to_signed(2414, LUT_AMPL_WIDTH),
		770 => to_signed(2417, LUT_AMPL_WIDTH),
		771 => to_signed(2420, LUT_AMPL_WIDTH),
		772 => to_signed(2423, LUT_AMPL_WIDTH),
		773 => to_signed(2426, LUT_AMPL_WIDTH),
		774 => to_signed(2429, LUT_AMPL_WIDTH),
		775 => to_signed(2432, LUT_AMPL_WIDTH),
		776 => to_signed(2436, LUT_AMPL_WIDTH),
		777 => to_signed(2439, LUT_AMPL_WIDTH),
		778 => to_signed(2442, LUT_AMPL_WIDTH),
		779 => to_signed(2445, LUT_AMPL_WIDTH),
		780 => to_signed(2448, LUT_AMPL_WIDTH),
		781 => to_signed(2451, LUT_AMPL_WIDTH),
		782 => to_signed(2454, LUT_AMPL_WIDTH),
		783 => to_signed(2457, LUT_AMPL_WIDTH),
		784 => to_signed(2461, LUT_AMPL_WIDTH),
		785 => to_signed(2464, LUT_AMPL_WIDTH),
		786 => to_signed(2467, LUT_AMPL_WIDTH),
		787 => to_signed(2470, LUT_AMPL_WIDTH),
		788 => to_signed(2473, LUT_AMPL_WIDTH),
		789 => to_signed(2476, LUT_AMPL_WIDTH),
		790 => to_signed(2479, LUT_AMPL_WIDTH),
		791 => to_signed(2483, LUT_AMPL_WIDTH),
		792 => to_signed(2486, LUT_AMPL_WIDTH),
		793 => to_signed(2489, LUT_AMPL_WIDTH),
		794 => to_signed(2492, LUT_AMPL_WIDTH),
		795 => to_signed(2495, LUT_AMPL_WIDTH),
		796 => to_signed(2498, LUT_AMPL_WIDTH),
		797 => to_signed(2501, LUT_AMPL_WIDTH),
		798 => to_signed(2504, LUT_AMPL_WIDTH),
		799 => to_signed(2508, LUT_AMPL_WIDTH),
		800 => to_signed(2511, LUT_AMPL_WIDTH),
		801 => to_signed(2514, LUT_AMPL_WIDTH),
		802 => to_signed(2517, LUT_AMPL_WIDTH),
		803 => to_signed(2520, LUT_AMPL_WIDTH),
		804 => to_signed(2523, LUT_AMPL_WIDTH),
		805 => to_signed(2526, LUT_AMPL_WIDTH),
		806 => to_signed(2530, LUT_AMPL_WIDTH),
		807 => to_signed(2533, LUT_AMPL_WIDTH),
		808 => to_signed(2536, LUT_AMPL_WIDTH),
		809 => to_signed(2539, LUT_AMPL_WIDTH),
		810 => to_signed(2542, LUT_AMPL_WIDTH),
		811 => to_signed(2545, LUT_AMPL_WIDTH),
		812 => to_signed(2548, LUT_AMPL_WIDTH),
		813 => to_signed(2551, LUT_AMPL_WIDTH),
		814 => to_signed(2555, LUT_AMPL_WIDTH),
		815 => to_signed(2558, LUT_AMPL_WIDTH),
		816 => to_signed(2561, LUT_AMPL_WIDTH),
		817 => to_signed(2564, LUT_AMPL_WIDTH),
		818 => to_signed(2567, LUT_AMPL_WIDTH),
		819 => to_signed(2570, LUT_AMPL_WIDTH),
		820 => to_signed(2573, LUT_AMPL_WIDTH),
		821 => to_signed(2577, LUT_AMPL_WIDTH),
		822 => to_signed(2580, LUT_AMPL_WIDTH),
		823 => to_signed(2583, LUT_AMPL_WIDTH),
		824 => to_signed(2586, LUT_AMPL_WIDTH),
		825 => to_signed(2589, LUT_AMPL_WIDTH),
		826 => to_signed(2592, LUT_AMPL_WIDTH),
		827 => to_signed(2595, LUT_AMPL_WIDTH),
		828 => to_signed(2598, LUT_AMPL_WIDTH),
		829 => to_signed(2602, LUT_AMPL_WIDTH),
		830 => to_signed(2605, LUT_AMPL_WIDTH),
		831 => to_signed(2608, LUT_AMPL_WIDTH),
		832 => to_signed(2611, LUT_AMPL_WIDTH),
		833 => to_signed(2614, LUT_AMPL_WIDTH),
		834 => to_signed(2617, LUT_AMPL_WIDTH),
		835 => to_signed(2620, LUT_AMPL_WIDTH),
		836 => to_signed(2623, LUT_AMPL_WIDTH),
		837 => to_signed(2627, LUT_AMPL_WIDTH),
		838 => to_signed(2630, LUT_AMPL_WIDTH),
		839 => to_signed(2633, LUT_AMPL_WIDTH),
		840 => to_signed(2636, LUT_AMPL_WIDTH),
		841 => to_signed(2639, LUT_AMPL_WIDTH),
		842 => to_signed(2642, LUT_AMPL_WIDTH),
		843 => to_signed(2645, LUT_AMPL_WIDTH),
		844 => to_signed(2649, LUT_AMPL_WIDTH),
		845 => to_signed(2652, LUT_AMPL_WIDTH),
		846 => to_signed(2655, LUT_AMPL_WIDTH),
		847 => to_signed(2658, LUT_AMPL_WIDTH),
		848 => to_signed(2661, LUT_AMPL_WIDTH),
		849 => to_signed(2664, LUT_AMPL_WIDTH),
		850 => to_signed(2667, LUT_AMPL_WIDTH),
		851 => to_signed(2670, LUT_AMPL_WIDTH),
		852 => to_signed(2674, LUT_AMPL_WIDTH),
		853 => to_signed(2677, LUT_AMPL_WIDTH),
		854 => to_signed(2680, LUT_AMPL_WIDTH),
		855 => to_signed(2683, LUT_AMPL_WIDTH),
		856 => to_signed(2686, LUT_AMPL_WIDTH),
		857 => to_signed(2689, LUT_AMPL_WIDTH),
		858 => to_signed(2692, LUT_AMPL_WIDTH),
		859 => to_signed(2695, LUT_AMPL_WIDTH),
		860 => to_signed(2699, LUT_AMPL_WIDTH),
		861 => to_signed(2702, LUT_AMPL_WIDTH),
		862 => to_signed(2705, LUT_AMPL_WIDTH),
		863 => to_signed(2708, LUT_AMPL_WIDTH),
		864 => to_signed(2711, LUT_AMPL_WIDTH),
		865 => to_signed(2714, LUT_AMPL_WIDTH),
		866 => to_signed(2717, LUT_AMPL_WIDTH),
		867 => to_signed(2721, LUT_AMPL_WIDTH),
		868 => to_signed(2724, LUT_AMPL_WIDTH),
		869 => to_signed(2727, LUT_AMPL_WIDTH),
		870 => to_signed(2730, LUT_AMPL_WIDTH),
		871 => to_signed(2733, LUT_AMPL_WIDTH),
		872 => to_signed(2736, LUT_AMPL_WIDTH),
		873 => to_signed(2739, LUT_AMPL_WIDTH),
		874 => to_signed(2742, LUT_AMPL_WIDTH),
		875 => to_signed(2746, LUT_AMPL_WIDTH),
		876 => to_signed(2749, LUT_AMPL_WIDTH),
		877 => to_signed(2752, LUT_AMPL_WIDTH),
		878 => to_signed(2755, LUT_AMPL_WIDTH),
		879 => to_signed(2758, LUT_AMPL_WIDTH),
		880 => to_signed(2761, LUT_AMPL_WIDTH),
		881 => to_signed(2764, LUT_AMPL_WIDTH),
		882 => to_signed(2767, LUT_AMPL_WIDTH),
		883 => to_signed(2771, LUT_AMPL_WIDTH),
		884 => to_signed(2774, LUT_AMPL_WIDTH),
		885 => to_signed(2777, LUT_AMPL_WIDTH),
		886 => to_signed(2780, LUT_AMPL_WIDTH),
		887 => to_signed(2783, LUT_AMPL_WIDTH),
		888 => to_signed(2786, LUT_AMPL_WIDTH),
		889 => to_signed(2789, LUT_AMPL_WIDTH),
		890 => to_signed(2793, LUT_AMPL_WIDTH),
		891 => to_signed(2796, LUT_AMPL_WIDTH),
		892 => to_signed(2799, LUT_AMPL_WIDTH),
		893 => to_signed(2802, LUT_AMPL_WIDTH),
		894 => to_signed(2805, LUT_AMPL_WIDTH),
		895 => to_signed(2808, LUT_AMPL_WIDTH),
		896 => to_signed(2811, LUT_AMPL_WIDTH),
		897 => to_signed(2814, LUT_AMPL_WIDTH),
		898 => to_signed(2818, LUT_AMPL_WIDTH),
		899 => to_signed(2821, LUT_AMPL_WIDTH),
		900 => to_signed(2824, LUT_AMPL_WIDTH),
		901 => to_signed(2827, LUT_AMPL_WIDTH),
		902 => to_signed(2830, LUT_AMPL_WIDTH),
		903 => to_signed(2833, LUT_AMPL_WIDTH),
		904 => to_signed(2836, LUT_AMPL_WIDTH),
		905 => to_signed(2839, LUT_AMPL_WIDTH),
		906 => to_signed(2843, LUT_AMPL_WIDTH),
		907 => to_signed(2846, LUT_AMPL_WIDTH),
		908 => to_signed(2849, LUT_AMPL_WIDTH),
		909 => to_signed(2852, LUT_AMPL_WIDTH),
		910 => to_signed(2855, LUT_AMPL_WIDTH),
		911 => to_signed(2858, LUT_AMPL_WIDTH),
		912 => to_signed(2861, LUT_AMPL_WIDTH),
		913 => to_signed(2865, LUT_AMPL_WIDTH),
		914 => to_signed(2868, LUT_AMPL_WIDTH),
		915 => to_signed(2871, LUT_AMPL_WIDTH),
		916 => to_signed(2874, LUT_AMPL_WIDTH),
		917 => to_signed(2877, LUT_AMPL_WIDTH),
		918 => to_signed(2880, LUT_AMPL_WIDTH),
		919 => to_signed(2883, LUT_AMPL_WIDTH),
		920 => to_signed(2886, LUT_AMPL_WIDTH),
		921 => to_signed(2890, LUT_AMPL_WIDTH),
		922 => to_signed(2893, LUT_AMPL_WIDTH),
		923 => to_signed(2896, LUT_AMPL_WIDTH),
		924 => to_signed(2899, LUT_AMPL_WIDTH),
		925 => to_signed(2902, LUT_AMPL_WIDTH),
		926 => to_signed(2905, LUT_AMPL_WIDTH),
		927 => to_signed(2908, LUT_AMPL_WIDTH),
		928 => to_signed(2911, LUT_AMPL_WIDTH),
		929 => to_signed(2915, LUT_AMPL_WIDTH),
		930 => to_signed(2918, LUT_AMPL_WIDTH),
		931 => to_signed(2921, LUT_AMPL_WIDTH),
		932 => to_signed(2924, LUT_AMPL_WIDTH),
		933 => to_signed(2927, LUT_AMPL_WIDTH),
		934 => to_signed(2930, LUT_AMPL_WIDTH),
		935 => to_signed(2933, LUT_AMPL_WIDTH),
		936 => to_signed(2936, LUT_AMPL_WIDTH),
		937 => to_signed(2940, LUT_AMPL_WIDTH),
		938 => to_signed(2943, LUT_AMPL_WIDTH),
		939 => to_signed(2946, LUT_AMPL_WIDTH),
		940 => to_signed(2949, LUT_AMPL_WIDTH),
		941 => to_signed(2952, LUT_AMPL_WIDTH),
		942 => to_signed(2955, LUT_AMPL_WIDTH),
		943 => to_signed(2958, LUT_AMPL_WIDTH),
		944 => to_signed(2962, LUT_AMPL_WIDTH),
		945 => to_signed(2965, LUT_AMPL_WIDTH),
		946 => to_signed(2968, LUT_AMPL_WIDTH),
		947 => to_signed(2971, LUT_AMPL_WIDTH),
		948 => to_signed(2974, LUT_AMPL_WIDTH),
		949 => to_signed(2977, LUT_AMPL_WIDTH),
		950 => to_signed(2980, LUT_AMPL_WIDTH),
		951 => to_signed(2983, LUT_AMPL_WIDTH),
		952 => to_signed(2987, LUT_AMPL_WIDTH),
		953 => to_signed(2990, LUT_AMPL_WIDTH),
		954 => to_signed(2993, LUT_AMPL_WIDTH),
		955 => to_signed(2996, LUT_AMPL_WIDTH),
		956 => to_signed(2999, LUT_AMPL_WIDTH),
		957 => to_signed(3002, LUT_AMPL_WIDTH),
		958 => to_signed(3005, LUT_AMPL_WIDTH),
		959 => to_signed(3008, LUT_AMPL_WIDTH),
		960 => to_signed(3012, LUT_AMPL_WIDTH),
		961 => to_signed(3015, LUT_AMPL_WIDTH),
		962 => to_signed(3018, LUT_AMPL_WIDTH),
		963 => to_signed(3021, LUT_AMPL_WIDTH),
		964 => to_signed(3024, LUT_AMPL_WIDTH),
		965 => to_signed(3027, LUT_AMPL_WIDTH),
		966 => to_signed(3030, LUT_AMPL_WIDTH),
		967 => to_signed(3033, LUT_AMPL_WIDTH),
		968 => to_signed(3037, LUT_AMPL_WIDTH),
		969 => to_signed(3040, LUT_AMPL_WIDTH),
		970 => to_signed(3043, LUT_AMPL_WIDTH),
		971 => to_signed(3046, LUT_AMPL_WIDTH),
		972 => to_signed(3049, LUT_AMPL_WIDTH),
		973 => to_signed(3052, LUT_AMPL_WIDTH),
		974 => to_signed(3055, LUT_AMPL_WIDTH),
		975 => to_signed(3059, LUT_AMPL_WIDTH),
		976 => to_signed(3062, LUT_AMPL_WIDTH),
		977 => to_signed(3065, LUT_AMPL_WIDTH),
		978 => to_signed(3068, LUT_AMPL_WIDTH),
		979 => to_signed(3071, LUT_AMPL_WIDTH),
		980 => to_signed(3074, LUT_AMPL_WIDTH),
		981 => to_signed(3077, LUT_AMPL_WIDTH),
		982 => to_signed(3080, LUT_AMPL_WIDTH),
		983 => to_signed(3084, LUT_AMPL_WIDTH),
		984 => to_signed(3087, LUT_AMPL_WIDTH),
		985 => to_signed(3090, LUT_AMPL_WIDTH),
		986 => to_signed(3093, LUT_AMPL_WIDTH),
		987 => to_signed(3096, LUT_AMPL_WIDTH),
		988 => to_signed(3099, LUT_AMPL_WIDTH),
		989 => to_signed(3102, LUT_AMPL_WIDTH),
		990 => to_signed(3105, LUT_AMPL_WIDTH),
		991 => to_signed(3109, LUT_AMPL_WIDTH),
		992 => to_signed(3112, LUT_AMPL_WIDTH),
		993 => to_signed(3115, LUT_AMPL_WIDTH),
		994 => to_signed(3118, LUT_AMPL_WIDTH),
		995 => to_signed(3121, LUT_AMPL_WIDTH),
		996 => to_signed(3124, LUT_AMPL_WIDTH),
		997 => to_signed(3127, LUT_AMPL_WIDTH),
		998 => to_signed(3130, LUT_AMPL_WIDTH),
		999 => to_signed(3134, LUT_AMPL_WIDTH),
		1000 => to_signed(3137, LUT_AMPL_WIDTH),
		1001 => to_signed(3140, LUT_AMPL_WIDTH),
		1002 => to_signed(3143, LUT_AMPL_WIDTH),
		1003 => to_signed(3146, LUT_AMPL_WIDTH),
		1004 => to_signed(3149, LUT_AMPL_WIDTH),
		1005 => to_signed(3152, LUT_AMPL_WIDTH),
		1006 => to_signed(3155, LUT_AMPL_WIDTH),
		1007 => to_signed(3159, LUT_AMPL_WIDTH),
		1008 => to_signed(3162, LUT_AMPL_WIDTH),
		1009 => to_signed(3165, LUT_AMPL_WIDTH),
		1010 => to_signed(3168, LUT_AMPL_WIDTH),
		1011 => to_signed(3171, LUT_AMPL_WIDTH),
		1012 => to_signed(3174, LUT_AMPL_WIDTH),
		1013 => to_signed(3177, LUT_AMPL_WIDTH),
		1014 => to_signed(3180, LUT_AMPL_WIDTH),
		1015 => to_signed(3184, LUT_AMPL_WIDTH),
		1016 => to_signed(3187, LUT_AMPL_WIDTH),
		1017 => to_signed(3190, LUT_AMPL_WIDTH),
		1018 => to_signed(3193, LUT_AMPL_WIDTH),
		1019 => to_signed(3196, LUT_AMPL_WIDTH),
		1020 => to_signed(3199, LUT_AMPL_WIDTH),
		1021 => to_signed(3202, LUT_AMPL_WIDTH),
		1022 => to_signed(3205, LUT_AMPL_WIDTH),
		1023 => to_signed(3209, LUT_AMPL_WIDTH),
		1024 => to_signed(3212, LUT_AMPL_WIDTH),
		1025 => to_signed(3215, LUT_AMPL_WIDTH),
		1026 => to_signed(3218, LUT_AMPL_WIDTH),
		1027 => to_signed(3221, LUT_AMPL_WIDTH),
		1028 => to_signed(3224, LUT_AMPL_WIDTH),
		1029 => to_signed(3227, LUT_AMPL_WIDTH),
		1030 => to_signed(3230, LUT_AMPL_WIDTH),
		1031 => to_signed(3234, LUT_AMPL_WIDTH),
		1032 => to_signed(3237, LUT_AMPL_WIDTH),
		1033 => to_signed(3240, LUT_AMPL_WIDTH),
		1034 => to_signed(3243, LUT_AMPL_WIDTH),
		1035 => to_signed(3246, LUT_AMPL_WIDTH),
		1036 => to_signed(3249, LUT_AMPL_WIDTH),
		1037 => to_signed(3252, LUT_AMPL_WIDTH),
		1038 => to_signed(3255, LUT_AMPL_WIDTH),
		1039 => to_signed(3259, LUT_AMPL_WIDTH),
		1040 => to_signed(3262, LUT_AMPL_WIDTH),
		1041 => to_signed(3265, LUT_AMPL_WIDTH),
		1042 => to_signed(3268, LUT_AMPL_WIDTH),
		1043 => to_signed(3271, LUT_AMPL_WIDTH),
		1044 => to_signed(3274, LUT_AMPL_WIDTH),
		1045 => to_signed(3277, LUT_AMPL_WIDTH),
		1046 => to_signed(3281, LUT_AMPL_WIDTH),
		1047 => to_signed(3284, LUT_AMPL_WIDTH),
		1048 => to_signed(3287, LUT_AMPL_WIDTH),
		1049 => to_signed(3290, LUT_AMPL_WIDTH),
		1050 => to_signed(3293, LUT_AMPL_WIDTH),
		1051 => to_signed(3296, LUT_AMPL_WIDTH),
		1052 => to_signed(3299, LUT_AMPL_WIDTH),
		1053 => to_signed(3302, LUT_AMPL_WIDTH),
		1054 => to_signed(3306, LUT_AMPL_WIDTH),
		1055 => to_signed(3309, LUT_AMPL_WIDTH),
		1056 => to_signed(3312, LUT_AMPL_WIDTH),
		1057 => to_signed(3315, LUT_AMPL_WIDTH),
		1058 => to_signed(3318, LUT_AMPL_WIDTH),
		1059 => to_signed(3321, LUT_AMPL_WIDTH),
		1060 => to_signed(3324, LUT_AMPL_WIDTH),
		1061 => to_signed(3327, LUT_AMPL_WIDTH),
		1062 => to_signed(3331, LUT_AMPL_WIDTH),
		1063 => to_signed(3334, LUT_AMPL_WIDTH),
		1064 => to_signed(3337, LUT_AMPL_WIDTH),
		1065 => to_signed(3340, LUT_AMPL_WIDTH),
		1066 => to_signed(3343, LUT_AMPL_WIDTH),
		1067 => to_signed(3346, LUT_AMPL_WIDTH),
		1068 => to_signed(3349, LUT_AMPL_WIDTH),
		1069 => to_signed(3352, LUT_AMPL_WIDTH),
		1070 => to_signed(3356, LUT_AMPL_WIDTH),
		1071 => to_signed(3359, LUT_AMPL_WIDTH),
		1072 => to_signed(3362, LUT_AMPL_WIDTH),
		1073 => to_signed(3365, LUT_AMPL_WIDTH),
		1074 => to_signed(3368, LUT_AMPL_WIDTH),
		1075 => to_signed(3371, LUT_AMPL_WIDTH),
		1076 => to_signed(3374, LUT_AMPL_WIDTH),
		1077 => to_signed(3377, LUT_AMPL_WIDTH),
		1078 => to_signed(3381, LUT_AMPL_WIDTH),
		1079 => to_signed(3384, LUT_AMPL_WIDTH),
		1080 => to_signed(3387, LUT_AMPL_WIDTH),
		1081 => to_signed(3390, LUT_AMPL_WIDTH),
		1082 => to_signed(3393, LUT_AMPL_WIDTH),
		1083 => to_signed(3396, LUT_AMPL_WIDTH),
		1084 => to_signed(3399, LUT_AMPL_WIDTH),
		1085 => to_signed(3402, LUT_AMPL_WIDTH),
		1086 => to_signed(3406, LUT_AMPL_WIDTH),
		1087 => to_signed(3409, LUT_AMPL_WIDTH),
		1088 => to_signed(3412, LUT_AMPL_WIDTH),
		1089 => to_signed(3415, LUT_AMPL_WIDTH),
		1090 => to_signed(3418, LUT_AMPL_WIDTH),
		1091 => to_signed(3421, LUT_AMPL_WIDTH),
		1092 => to_signed(3424, LUT_AMPL_WIDTH),
		1093 => to_signed(3427, LUT_AMPL_WIDTH),
		1094 => to_signed(3430, LUT_AMPL_WIDTH),
		1095 => to_signed(3434, LUT_AMPL_WIDTH),
		1096 => to_signed(3437, LUT_AMPL_WIDTH),
		1097 => to_signed(3440, LUT_AMPL_WIDTH),
		1098 => to_signed(3443, LUT_AMPL_WIDTH),
		1099 => to_signed(3446, LUT_AMPL_WIDTH),
		1100 => to_signed(3449, LUT_AMPL_WIDTH),
		1101 => to_signed(3452, LUT_AMPL_WIDTH),
		1102 => to_signed(3455, LUT_AMPL_WIDTH),
		1103 => to_signed(3459, LUT_AMPL_WIDTH),
		1104 => to_signed(3462, LUT_AMPL_WIDTH),
		1105 => to_signed(3465, LUT_AMPL_WIDTH),
		1106 => to_signed(3468, LUT_AMPL_WIDTH),
		1107 => to_signed(3471, LUT_AMPL_WIDTH),
		1108 => to_signed(3474, LUT_AMPL_WIDTH),
		1109 => to_signed(3477, LUT_AMPL_WIDTH),
		1110 => to_signed(3480, LUT_AMPL_WIDTH),
		1111 => to_signed(3484, LUT_AMPL_WIDTH),
		1112 => to_signed(3487, LUT_AMPL_WIDTH),
		1113 => to_signed(3490, LUT_AMPL_WIDTH),
		1114 => to_signed(3493, LUT_AMPL_WIDTH),
		1115 => to_signed(3496, LUT_AMPL_WIDTH),
		1116 => to_signed(3499, LUT_AMPL_WIDTH),
		1117 => to_signed(3502, LUT_AMPL_WIDTH),
		1118 => to_signed(3505, LUT_AMPL_WIDTH),
		1119 => to_signed(3509, LUT_AMPL_WIDTH),
		1120 => to_signed(3512, LUT_AMPL_WIDTH),
		1121 => to_signed(3515, LUT_AMPL_WIDTH),
		1122 => to_signed(3518, LUT_AMPL_WIDTH),
		1123 => to_signed(3521, LUT_AMPL_WIDTH),
		1124 => to_signed(3524, LUT_AMPL_WIDTH),
		1125 => to_signed(3527, LUT_AMPL_WIDTH),
		1126 => to_signed(3530, LUT_AMPL_WIDTH),
		1127 => to_signed(3534, LUT_AMPL_WIDTH),
		1128 => to_signed(3537, LUT_AMPL_WIDTH),
		1129 => to_signed(3540, LUT_AMPL_WIDTH),
		1130 => to_signed(3543, LUT_AMPL_WIDTH),
		1131 => to_signed(3546, LUT_AMPL_WIDTH),
		1132 => to_signed(3549, LUT_AMPL_WIDTH),
		1133 => to_signed(3552, LUT_AMPL_WIDTH),
		1134 => to_signed(3555, LUT_AMPL_WIDTH),
		1135 => to_signed(3559, LUT_AMPL_WIDTH),
		1136 => to_signed(3562, LUT_AMPL_WIDTH),
		1137 => to_signed(3565, LUT_AMPL_WIDTH),
		1138 => to_signed(3568, LUT_AMPL_WIDTH),
		1139 => to_signed(3571, LUT_AMPL_WIDTH),
		1140 => to_signed(3574, LUT_AMPL_WIDTH),
		1141 => to_signed(3577, LUT_AMPL_WIDTH),
		1142 => to_signed(3580, LUT_AMPL_WIDTH),
		1143 => to_signed(3584, LUT_AMPL_WIDTH),
		1144 => to_signed(3587, LUT_AMPL_WIDTH),
		1145 => to_signed(3590, LUT_AMPL_WIDTH),
		1146 => to_signed(3593, LUT_AMPL_WIDTH),
		1147 => to_signed(3596, LUT_AMPL_WIDTH),
		1148 => to_signed(3599, LUT_AMPL_WIDTH),
		1149 => to_signed(3602, LUT_AMPL_WIDTH),
		1150 => to_signed(3605, LUT_AMPL_WIDTH),
		1151 => to_signed(3609, LUT_AMPL_WIDTH),
		1152 => to_signed(3612, LUT_AMPL_WIDTH),
		1153 => to_signed(3615, LUT_AMPL_WIDTH),
		1154 => to_signed(3618, LUT_AMPL_WIDTH),
		1155 => to_signed(3621, LUT_AMPL_WIDTH),
		1156 => to_signed(3624, LUT_AMPL_WIDTH),
		1157 => to_signed(3627, LUT_AMPL_WIDTH),
		1158 => to_signed(3630, LUT_AMPL_WIDTH),
		1159 => to_signed(3634, LUT_AMPL_WIDTH),
		1160 => to_signed(3637, LUT_AMPL_WIDTH),
		1161 => to_signed(3640, LUT_AMPL_WIDTH),
		1162 => to_signed(3643, LUT_AMPL_WIDTH),
		1163 => to_signed(3646, LUT_AMPL_WIDTH),
		1164 => to_signed(3649, LUT_AMPL_WIDTH),
		1165 => to_signed(3652, LUT_AMPL_WIDTH),
		1166 => to_signed(3655, LUT_AMPL_WIDTH),
		1167 => to_signed(3658, LUT_AMPL_WIDTH),
		1168 => to_signed(3662, LUT_AMPL_WIDTH),
		1169 => to_signed(3665, LUT_AMPL_WIDTH),
		1170 => to_signed(3668, LUT_AMPL_WIDTH),
		1171 => to_signed(3671, LUT_AMPL_WIDTH),
		1172 => to_signed(3674, LUT_AMPL_WIDTH),
		1173 => to_signed(3677, LUT_AMPL_WIDTH),
		1174 => to_signed(3680, LUT_AMPL_WIDTH),
		1175 => to_signed(3683, LUT_AMPL_WIDTH),
		1176 => to_signed(3687, LUT_AMPL_WIDTH),
		1177 => to_signed(3690, LUT_AMPL_WIDTH),
		1178 => to_signed(3693, LUT_AMPL_WIDTH),
		1179 => to_signed(3696, LUT_AMPL_WIDTH),
		1180 => to_signed(3699, LUT_AMPL_WIDTH),
		1181 => to_signed(3702, LUT_AMPL_WIDTH),
		1182 => to_signed(3705, LUT_AMPL_WIDTH),
		1183 => to_signed(3708, LUT_AMPL_WIDTH),
		1184 => to_signed(3712, LUT_AMPL_WIDTH),
		1185 => to_signed(3715, LUT_AMPL_WIDTH),
		1186 => to_signed(3718, LUT_AMPL_WIDTH),
		1187 => to_signed(3721, LUT_AMPL_WIDTH),
		1188 => to_signed(3724, LUT_AMPL_WIDTH),
		1189 => to_signed(3727, LUT_AMPL_WIDTH),
		1190 => to_signed(3730, LUT_AMPL_WIDTH),
		1191 => to_signed(3733, LUT_AMPL_WIDTH),
		1192 => to_signed(3737, LUT_AMPL_WIDTH),
		1193 => to_signed(3740, LUT_AMPL_WIDTH),
		1194 => to_signed(3743, LUT_AMPL_WIDTH),
		1195 => to_signed(3746, LUT_AMPL_WIDTH),
		1196 => to_signed(3749, LUT_AMPL_WIDTH),
		1197 => to_signed(3752, LUT_AMPL_WIDTH),
		1198 => to_signed(3755, LUT_AMPL_WIDTH),
		1199 => to_signed(3758, LUT_AMPL_WIDTH),
		1200 => to_signed(3761, LUT_AMPL_WIDTH),
		1201 => to_signed(3765, LUT_AMPL_WIDTH),
		1202 => to_signed(3768, LUT_AMPL_WIDTH),
		1203 => to_signed(3771, LUT_AMPL_WIDTH),
		1204 => to_signed(3774, LUT_AMPL_WIDTH),
		1205 => to_signed(3777, LUT_AMPL_WIDTH),
		1206 => to_signed(3780, LUT_AMPL_WIDTH),
		1207 => to_signed(3783, LUT_AMPL_WIDTH),
		1208 => to_signed(3786, LUT_AMPL_WIDTH),
		1209 => to_signed(3790, LUT_AMPL_WIDTH),
		1210 => to_signed(3793, LUT_AMPL_WIDTH),
		1211 => to_signed(3796, LUT_AMPL_WIDTH),
		1212 => to_signed(3799, LUT_AMPL_WIDTH),
		1213 => to_signed(3802, LUT_AMPL_WIDTH),
		1214 => to_signed(3805, LUT_AMPL_WIDTH),
		1215 => to_signed(3808, LUT_AMPL_WIDTH),
		1216 => to_signed(3811, LUT_AMPL_WIDTH),
		1217 => to_signed(3815, LUT_AMPL_WIDTH),
		1218 => to_signed(3818, LUT_AMPL_WIDTH),
		1219 => to_signed(3821, LUT_AMPL_WIDTH),
		1220 => to_signed(3824, LUT_AMPL_WIDTH),
		1221 => to_signed(3827, LUT_AMPL_WIDTH),
		1222 => to_signed(3830, LUT_AMPL_WIDTH),
		1223 => to_signed(3833, LUT_AMPL_WIDTH),
		1224 => to_signed(3836, LUT_AMPL_WIDTH),
		1225 => to_signed(3839, LUT_AMPL_WIDTH),
		1226 => to_signed(3843, LUT_AMPL_WIDTH),
		1227 => to_signed(3846, LUT_AMPL_WIDTH),
		1228 => to_signed(3849, LUT_AMPL_WIDTH),
		1229 => to_signed(3852, LUT_AMPL_WIDTH),
		1230 => to_signed(3855, LUT_AMPL_WIDTH),
		1231 => to_signed(3858, LUT_AMPL_WIDTH),
		1232 => to_signed(3861, LUT_AMPL_WIDTH),
		1233 => to_signed(3864, LUT_AMPL_WIDTH),
		1234 => to_signed(3868, LUT_AMPL_WIDTH),
		1235 => to_signed(3871, LUT_AMPL_WIDTH),
		1236 => to_signed(3874, LUT_AMPL_WIDTH),
		1237 => to_signed(3877, LUT_AMPL_WIDTH),
		1238 => to_signed(3880, LUT_AMPL_WIDTH),
		1239 => to_signed(3883, LUT_AMPL_WIDTH),
		1240 => to_signed(3886, LUT_AMPL_WIDTH),
		1241 => to_signed(3889, LUT_AMPL_WIDTH),
		1242 => to_signed(3893, LUT_AMPL_WIDTH),
		1243 => to_signed(3896, LUT_AMPL_WIDTH),
		1244 => to_signed(3899, LUT_AMPL_WIDTH),
		1245 => to_signed(3902, LUT_AMPL_WIDTH),
		1246 => to_signed(3905, LUT_AMPL_WIDTH),
		1247 => to_signed(3908, LUT_AMPL_WIDTH),
		1248 => to_signed(3911, LUT_AMPL_WIDTH),
		1249 => to_signed(3914, LUT_AMPL_WIDTH),
		1250 => to_signed(3917, LUT_AMPL_WIDTH),
		1251 => to_signed(3921, LUT_AMPL_WIDTH),
		1252 => to_signed(3924, LUT_AMPL_WIDTH),
		1253 => to_signed(3927, LUT_AMPL_WIDTH),
		1254 => to_signed(3930, LUT_AMPL_WIDTH),
		1255 => to_signed(3933, LUT_AMPL_WIDTH),
		1256 => to_signed(3936, LUT_AMPL_WIDTH),
		1257 => to_signed(3939, LUT_AMPL_WIDTH),
		1258 => to_signed(3942, LUT_AMPL_WIDTH),
		1259 => to_signed(3946, LUT_AMPL_WIDTH),
		1260 => to_signed(3949, LUT_AMPL_WIDTH),
		1261 => to_signed(3952, LUT_AMPL_WIDTH),
		1262 => to_signed(3955, LUT_AMPL_WIDTH),
		1263 => to_signed(3958, LUT_AMPL_WIDTH),
		1264 => to_signed(3961, LUT_AMPL_WIDTH),
		1265 => to_signed(3964, LUT_AMPL_WIDTH),
		1266 => to_signed(3967, LUT_AMPL_WIDTH),
		1267 => to_signed(3970, LUT_AMPL_WIDTH),
		1268 => to_signed(3974, LUT_AMPL_WIDTH),
		1269 => to_signed(3977, LUT_AMPL_WIDTH),
		1270 => to_signed(3980, LUT_AMPL_WIDTH),
		1271 => to_signed(3983, LUT_AMPL_WIDTH),
		1272 => to_signed(3986, LUT_AMPL_WIDTH),
		1273 => to_signed(3989, LUT_AMPL_WIDTH),
		1274 => to_signed(3992, LUT_AMPL_WIDTH),
		1275 => to_signed(3995, LUT_AMPL_WIDTH),
		1276 => to_signed(3999, LUT_AMPL_WIDTH),
		1277 => to_signed(4002, LUT_AMPL_WIDTH),
		1278 => to_signed(4005, LUT_AMPL_WIDTH),
		1279 => to_signed(4008, LUT_AMPL_WIDTH),
		1280 => to_signed(4011, LUT_AMPL_WIDTH),
		1281 => to_signed(4014, LUT_AMPL_WIDTH),
		1282 => to_signed(4017, LUT_AMPL_WIDTH),
		1283 => to_signed(4020, LUT_AMPL_WIDTH),
		1284 => to_signed(4024, LUT_AMPL_WIDTH),
		1285 => to_signed(4027, LUT_AMPL_WIDTH),
		1286 => to_signed(4030, LUT_AMPL_WIDTH),
		1287 => to_signed(4033, LUT_AMPL_WIDTH),
		1288 => to_signed(4036, LUT_AMPL_WIDTH),
		1289 => to_signed(4039, LUT_AMPL_WIDTH),
		1290 => to_signed(4042, LUT_AMPL_WIDTH),
		1291 => to_signed(4045, LUT_AMPL_WIDTH),
		1292 => to_signed(4048, LUT_AMPL_WIDTH),
		1293 => to_signed(4052, LUT_AMPL_WIDTH),
		1294 => to_signed(4055, LUT_AMPL_WIDTH),
		1295 => to_signed(4058, LUT_AMPL_WIDTH),
		1296 => to_signed(4061, LUT_AMPL_WIDTH),
		1297 => to_signed(4064, LUT_AMPL_WIDTH),
		1298 => to_signed(4067, LUT_AMPL_WIDTH),
		1299 => to_signed(4070, LUT_AMPL_WIDTH),
		1300 => to_signed(4073, LUT_AMPL_WIDTH),
		1301 => to_signed(4076, LUT_AMPL_WIDTH),
		1302 => to_signed(4080, LUT_AMPL_WIDTH),
		1303 => to_signed(4083, LUT_AMPL_WIDTH),
		1304 => to_signed(4086, LUT_AMPL_WIDTH),
		1305 => to_signed(4089, LUT_AMPL_WIDTH),
		1306 => to_signed(4092, LUT_AMPL_WIDTH),
		1307 => to_signed(4095, LUT_AMPL_WIDTH),
		1308 => to_signed(4098, LUT_AMPL_WIDTH),
		1309 => to_signed(4101, LUT_AMPL_WIDTH),
		1310 => to_signed(4105, LUT_AMPL_WIDTH),
		1311 => to_signed(4108, LUT_AMPL_WIDTH),
		1312 => to_signed(4111, LUT_AMPL_WIDTH),
		1313 => to_signed(4114, LUT_AMPL_WIDTH),
		1314 => to_signed(4117, LUT_AMPL_WIDTH),
		1315 => to_signed(4120, LUT_AMPL_WIDTH),
		1316 => to_signed(4123, LUT_AMPL_WIDTH),
		1317 => to_signed(4126, LUT_AMPL_WIDTH),
		1318 => to_signed(4129, LUT_AMPL_WIDTH),
		1319 => to_signed(4133, LUT_AMPL_WIDTH),
		1320 => to_signed(4136, LUT_AMPL_WIDTH),
		1321 => to_signed(4139, LUT_AMPL_WIDTH),
		1322 => to_signed(4142, LUT_AMPL_WIDTH),
		1323 => to_signed(4145, LUT_AMPL_WIDTH),
		1324 => to_signed(4148, LUT_AMPL_WIDTH),
		1325 => to_signed(4151, LUT_AMPL_WIDTH),
		1326 => to_signed(4154, LUT_AMPL_WIDTH),
		1327 => to_signed(4158, LUT_AMPL_WIDTH),
		1328 => to_signed(4161, LUT_AMPL_WIDTH),
		1329 => to_signed(4164, LUT_AMPL_WIDTH),
		1330 => to_signed(4167, LUT_AMPL_WIDTH),
		1331 => to_signed(4170, LUT_AMPL_WIDTH),
		1332 => to_signed(4173, LUT_AMPL_WIDTH),
		1333 => to_signed(4176, LUT_AMPL_WIDTH),
		1334 => to_signed(4179, LUT_AMPL_WIDTH),
		1335 => to_signed(4182, LUT_AMPL_WIDTH),
		1336 => to_signed(4186, LUT_AMPL_WIDTH),
		1337 => to_signed(4189, LUT_AMPL_WIDTH),
		1338 => to_signed(4192, LUT_AMPL_WIDTH),
		1339 => to_signed(4195, LUT_AMPL_WIDTH),
		1340 => to_signed(4198, LUT_AMPL_WIDTH),
		1341 => to_signed(4201, LUT_AMPL_WIDTH),
		1342 => to_signed(4204, LUT_AMPL_WIDTH),
		1343 => to_signed(4207, LUT_AMPL_WIDTH),
		1344 => to_signed(4210, LUT_AMPL_WIDTH),
		1345 => to_signed(4214, LUT_AMPL_WIDTH),
		1346 => to_signed(4217, LUT_AMPL_WIDTH),
		1347 => to_signed(4220, LUT_AMPL_WIDTH),
		1348 => to_signed(4223, LUT_AMPL_WIDTH),
		1349 => to_signed(4226, LUT_AMPL_WIDTH),
		1350 => to_signed(4229, LUT_AMPL_WIDTH),
		1351 => to_signed(4232, LUT_AMPL_WIDTH),
		1352 => to_signed(4235, LUT_AMPL_WIDTH),
		1353 => to_signed(4239, LUT_AMPL_WIDTH),
		1354 => to_signed(4242, LUT_AMPL_WIDTH),
		1355 => to_signed(4245, LUT_AMPL_WIDTH),
		1356 => to_signed(4248, LUT_AMPL_WIDTH),
		1357 => to_signed(4251, LUT_AMPL_WIDTH),
		1358 => to_signed(4254, LUT_AMPL_WIDTH),
		1359 => to_signed(4257, LUT_AMPL_WIDTH),
		1360 => to_signed(4260, LUT_AMPL_WIDTH),
		1361 => to_signed(4263, LUT_AMPL_WIDTH),
		1362 => to_signed(4267, LUT_AMPL_WIDTH),
		1363 => to_signed(4270, LUT_AMPL_WIDTH),
		1364 => to_signed(4273, LUT_AMPL_WIDTH),
		1365 => to_signed(4276, LUT_AMPL_WIDTH),
		1366 => to_signed(4279, LUT_AMPL_WIDTH),
		1367 => to_signed(4282, LUT_AMPL_WIDTH),
		1368 => to_signed(4285, LUT_AMPL_WIDTH),
		1369 => to_signed(4288, LUT_AMPL_WIDTH),
		1370 => to_signed(4291, LUT_AMPL_WIDTH),
		1371 => to_signed(4295, LUT_AMPL_WIDTH),
		1372 => to_signed(4298, LUT_AMPL_WIDTH),
		1373 => to_signed(4301, LUT_AMPL_WIDTH),
		1374 => to_signed(4304, LUT_AMPL_WIDTH),
		1375 => to_signed(4307, LUT_AMPL_WIDTH),
		1376 => to_signed(4310, LUT_AMPL_WIDTH),
		1377 => to_signed(4313, LUT_AMPL_WIDTH),
		1378 => to_signed(4316, LUT_AMPL_WIDTH),
		1379 => to_signed(4320, LUT_AMPL_WIDTH),
		1380 => to_signed(4323, LUT_AMPL_WIDTH),
		1381 => to_signed(4326, LUT_AMPL_WIDTH),
		1382 => to_signed(4329, LUT_AMPL_WIDTH),
		1383 => to_signed(4332, LUT_AMPL_WIDTH),
		1384 => to_signed(4335, LUT_AMPL_WIDTH),
		1385 => to_signed(4338, LUT_AMPL_WIDTH),
		1386 => to_signed(4341, LUT_AMPL_WIDTH),
		1387 => to_signed(4344, LUT_AMPL_WIDTH),
		1388 => to_signed(4348, LUT_AMPL_WIDTH),
		1389 => to_signed(4351, LUT_AMPL_WIDTH),
		1390 => to_signed(4354, LUT_AMPL_WIDTH),
		1391 => to_signed(4357, LUT_AMPL_WIDTH),
		1392 => to_signed(4360, LUT_AMPL_WIDTH),
		1393 => to_signed(4363, LUT_AMPL_WIDTH),
		1394 => to_signed(4366, LUT_AMPL_WIDTH),
		1395 => to_signed(4369, LUT_AMPL_WIDTH),
		1396 => to_signed(4372, LUT_AMPL_WIDTH),
		1397 => to_signed(4376, LUT_AMPL_WIDTH),
		1398 => to_signed(4379, LUT_AMPL_WIDTH),
		1399 => to_signed(4382, LUT_AMPL_WIDTH),
		1400 => to_signed(4385, LUT_AMPL_WIDTH),
		1401 => to_signed(4388, LUT_AMPL_WIDTH),
		1402 => to_signed(4391, LUT_AMPL_WIDTH),
		1403 => to_signed(4394, LUT_AMPL_WIDTH),
		1404 => to_signed(4397, LUT_AMPL_WIDTH),
		1405 => to_signed(4400, LUT_AMPL_WIDTH),
		1406 => to_signed(4404, LUT_AMPL_WIDTH),
		1407 => to_signed(4407, LUT_AMPL_WIDTH),
		1408 => to_signed(4410, LUT_AMPL_WIDTH),
		1409 => to_signed(4413, LUT_AMPL_WIDTH),
		1410 => to_signed(4416, LUT_AMPL_WIDTH),
		1411 => to_signed(4419, LUT_AMPL_WIDTH),
		1412 => to_signed(4422, LUT_AMPL_WIDTH),
		1413 => to_signed(4425, LUT_AMPL_WIDTH),
		1414 => to_signed(4428, LUT_AMPL_WIDTH),
		1415 => to_signed(4432, LUT_AMPL_WIDTH),
		1416 => to_signed(4435, LUT_AMPL_WIDTH),
		1417 => to_signed(4438, LUT_AMPL_WIDTH),
		1418 => to_signed(4441, LUT_AMPL_WIDTH),
		1419 => to_signed(4444, LUT_AMPL_WIDTH),
		1420 => to_signed(4447, LUT_AMPL_WIDTH),
		1421 => to_signed(4450, LUT_AMPL_WIDTH),
		1422 => to_signed(4453, LUT_AMPL_WIDTH),
		1423 => to_signed(4456, LUT_AMPL_WIDTH),
		1424 => to_signed(4460, LUT_AMPL_WIDTH),
		1425 => to_signed(4463, LUT_AMPL_WIDTH),
		1426 => to_signed(4466, LUT_AMPL_WIDTH),
		1427 => to_signed(4469, LUT_AMPL_WIDTH),
		1428 => to_signed(4472, LUT_AMPL_WIDTH),
		1429 => to_signed(4475, LUT_AMPL_WIDTH),
		1430 => to_signed(4478, LUT_AMPL_WIDTH),
		1431 => to_signed(4481, LUT_AMPL_WIDTH),
		1432 => to_signed(4485, LUT_AMPL_WIDTH),
		1433 => to_signed(4488, LUT_AMPL_WIDTH),
		1434 => to_signed(4491, LUT_AMPL_WIDTH),
		1435 => to_signed(4494, LUT_AMPL_WIDTH),
		1436 => to_signed(4497, LUT_AMPL_WIDTH),
		1437 => to_signed(4500, LUT_AMPL_WIDTH),
		1438 => to_signed(4503, LUT_AMPL_WIDTH),
		1439 => to_signed(4506, LUT_AMPL_WIDTH),
		1440 => to_signed(4509, LUT_AMPL_WIDTH),
		1441 => to_signed(4513, LUT_AMPL_WIDTH),
		1442 => to_signed(4516, LUT_AMPL_WIDTH),
		1443 => to_signed(4519, LUT_AMPL_WIDTH),
		1444 => to_signed(4522, LUT_AMPL_WIDTH),
		1445 => to_signed(4525, LUT_AMPL_WIDTH),
		1446 => to_signed(4528, LUT_AMPL_WIDTH),
		1447 => to_signed(4531, LUT_AMPL_WIDTH),
		1448 => to_signed(4534, LUT_AMPL_WIDTH),
		1449 => to_signed(4537, LUT_AMPL_WIDTH),
		1450 => to_signed(4541, LUT_AMPL_WIDTH),
		1451 => to_signed(4544, LUT_AMPL_WIDTH),
		1452 => to_signed(4547, LUT_AMPL_WIDTH),
		1453 => to_signed(4550, LUT_AMPL_WIDTH),
		1454 => to_signed(4553, LUT_AMPL_WIDTH),
		1455 => to_signed(4556, LUT_AMPL_WIDTH),
		1456 => to_signed(4559, LUT_AMPL_WIDTH),
		1457 => to_signed(4562, LUT_AMPL_WIDTH),
		1458 => to_signed(4565, LUT_AMPL_WIDTH),
		1459 => to_signed(4569, LUT_AMPL_WIDTH),
		1460 => to_signed(4572, LUT_AMPL_WIDTH),
		1461 => to_signed(4575, LUT_AMPL_WIDTH),
		1462 => to_signed(4578, LUT_AMPL_WIDTH),
		1463 => to_signed(4581, LUT_AMPL_WIDTH),
		1464 => to_signed(4584, LUT_AMPL_WIDTH),
		1465 => to_signed(4587, LUT_AMPL_WIDTH),
		1466 => to_signed(4590, LUT_AMPL_WIDTH),
		1467 => to_signed(4593, LUT_AMPL_WIDTH),
		1468 => to_signed(4597, LUT_AMPL_WIDTH),
		1469 => to_signed(4600, LUT_AMPL_WIDTH),
		1470 => to_signed(4603, LUT_AMPL_WIDTH),
		1471 => to_signed(4606, LUT_AMPL_WIDTH),
		1472 => to_signed(4609, LUT_AMPL_WIDTH),
		1473 => to_signed(4612, LUT_AMPL_WIDTH),
		1474 => to_signed(4615, LUT_AMPL_WIDTH),
		1475 => to_signed(4618, LUT_AMPL_WIDTH),
		1476 => to_signed(4621, LUT_AMPL_WIDTH),
		1477 => to_signed(4624, LUT_AMPL_WIDTH),
		1478 => to_signed(4628, LUT_AMPL_WIDTH),
		1479 => to_signed(4631, LUT_AMPL_WIDTH),
		1480 => to_signed(4634, LUT_AMPL_WIDTH),
		1481 => to_signed(4637, LUT_AMPL_WIDTH),
		1482 => to_signed(4640, LUT_AMPL_WIDTH),
		1483 => to_signed(4643, LUT_AMPL_WIDTH),
		1484 => to_signed(4646, LUT_AMPL_WIDTH),
		1485 => to_signed(4649, LUT_AMPL_WIDTH),
		1486 => to_signed(4652, LUT_AMPL_WIDTH),
		1487 => to_signed(4656, LUT_AMPL_WIDTH),
		1488 => to_signed(4659, LUT_AMPL_WIDTH),
		1489 => to_signed(4662, LUT_AMPL_WIDTH),
		1490 => to_signed(4665, LUT_AMPL_WIDTH),
		1491 => to_signed(4668, LUT_AMPL_WIDTH),
		1492 => to_signed(4671, LUT_AMPL_WIDTH),
		1493 => to_signed(4674, LUT_AMPL_WIDTH),
		1494 => to_signed(4677, LUT_AMPL_WIDTH),
		1495 => to_signed(4680, LUT_AMPL_WIDTH),
		1496 => to_signed(4684, LUT_AMPL_WIDTH),
		1497 => to_signed(4687, LUT_AMPL_WIDTH),
		1498 => to_signed(4690, LUT_AMPL_WIDTH),
		1499 => to_signed(4693, LUT_AMPL_WIDTH),
		1500 => to_signed(4696, LUT_AMPL_WIDTH),
		1501 => to_signed(4699, LUT_AMPL_WIDTH),
		1502 => to_signed(4702, LUT_AMPL_WIDTH),
		1503 => to_signed(4705, LUT_AMPL_WIDTH),
		1504 => to_signed(4708, LUT_AMPL_WIDTH),
		1505 => to_signed(4712, LUT_AMPL_WIDTH),
		1506 => to_signed(4715, LUT_AMPL_WIDTH),
		1507 => to_signed(4718, LUT_AMPL_WIDTH),
		1508 => to_signed(4721, LUT_AMPL_WIDTH),
		1509 => to_signed(4724, LUT_AMPL_WIDTH),
		1510 => to_signed(4727, LUT_AMPL_WIDTH),
		1511 => to_signed(4730, LUT_AMPL_WIDTH),
		1512 => to_signed(4733, LUT_AMPL_WIDTH),
		1513 => to_signed(4736, LUT_AMPL_WIDTH),
		1514 => to_signed(4740, LUT_AMPL_WIDTH),
		1515 => to_signed(4743, LUT_AMPL_WIDTH),
		1516 => to_signed(4746, LUT_AMPL_WIDTH),
		1517 => to_signed(4749, LUT_AMPL_WIDTH),
		1518 => to_signed(4752, LUT_AMPL_WIDTH),
		1519 => to_signed(4755, LUT_AMPL_WIDTH),
		1520 => to_signed(4758, LUT_AMPL_WIDTH),
		1521 => to_signed(4761, LUT_AMPL_WIDTH),
		1522 => to_signed(4764, LUT_AMPL_WIDTH),
		1523 => to_signed(4768, LUT_AMPL_WIDTH),
		1524 => to_signed(4771, LUT_AMPL_WIDTH),
		1525 => to_signed(4774, LUT_AMPL_WIDTH),
		1526 => to_signed(4777, LUT_AMPL_WIDTH),
		1527 => to_signed(4780, LUT_AMPL_WIDTH),
		1528 => to_signed(4783, LUT_AMPL_WIDTH),
		1529 => to_signed(4786, LUT_AMPL_WIDTH),
		1530 => to_signed(4789, LUT_AMPL_WIDTH),
		1531 => to_signed(4792, LUT_AMPL_WIDTH),
		1532 => to_signed(4795, LUT_AMPL_WIDTH),
		1533 => to_signed(4799, LUT_AMPL_WIDTH),
		1534 => to_signed(4802, LUT_AMPL_WIDTH),
		1535 => to_signed(4805, LUT_AMPL_WIDTH),
		1536 => to_signed(4808, LUT_AMPL_WIDTH),
		1537 => to_signed(4811, LUT_AMPL_WIDTH),
		1538 => to_signed(4814, LUT_AMPL_WIDTH),
		1539 => to_signed(4817, LUT_AMPL_WIDTH),
		1540 => to_signed(4820, LUT_AMPL_WIDTH),
		1541 => to_signed(4823, LUT_AMPL_WIDTH),
		1542 => to_signed(4827, LUT_AMPL_WIDTH),
		1543 => to_signed(4830, LUT_AMPL_WIDTH),
		1544 => to_signed(4833, LUT_AMPL_WIDTH),
		1545 => to_signed(4836, LUT_AMPL_WIDTH),
		1546 => to_signed(4839, LUT_AMPL_WIDTH),
		1547 => to_signed(4842, LUT_AMPL_WIDTH),
		1548 => to_signed(4845, LUT_AMPL_WIDTH),
		1549 => to_signed(4848, LUT_AMPL_WIDTH),
		1550 => to_signed(4851, LUT_AMPL_WIDTH),
		1551 => to_signed(4855, LUT_AMPL_WIDTH),
		1552 => to_signed(4858, LUT_AMPL_WIDTH),
		1553 => to_signed(4861, LUT_AMPL_WIDTH),
		1554 => to_signed(4864, LUT_AMPL_WIDTH),
		1555 => to_signed(4867, LUT_AMPL_WIDTH),
		1556 => to_signed(4870, LUT_AMPL_WIDTH),
		1557 => to_signed(4873, LUT_AMPL_WIDTH),
		1558 => to_signed(4876, LUT_AMPL_WIDTH),
		1559 => to_signed(4879, LUT_AMPL_WIDTH),
		1560 => to_signed(4882, LUT_AMPL_WIDTH),
		1561 => to_signed(4886, LUT_AMPL_WIDTH),
		1562 => to_signed(4889, LUT_AMPL_WIDTH),
		1563 => to_signed(4892, LUT_AMPL_WIDTH),
		1564 => to_signed(4895, LUT_AMPL_WIDTH),
		1565 => to_signed(4898, LUT_AMPL_WIDTH),
		1566 => to_signed(4901, LUT_AMPL_WIDTH),
		1567 => to_signed(4904, LUT_AMPL_WIDTH),
		1568 => to_signed(4907, LUT_AMPL_WIDTH),
		1569 => to_signed(4910, LUT_AMPL_WIDTH),
		1570 => to_signed(4914, LUT_AMPL_WIDTH),
		1571 => to_signed(4917, LUT_AMPL_WIDTH),
		1572 => to_signed(4920, LUT_AMPL_WIDTH),
		1573 => to_signed(4923, LUT_AMPL_WIDTH),
		1574 => to_signed(4926, LUT_AMPL_WIDTH),
		1575 => to_signed(4929, LUT_AMPL_WIDTH),
		1576 => to_signed(4932, LUT_AMPL_WIDTH),
		1577 => to_signed(4935, LUT_AMPL_WIDTH),
		1578 => to_signed(4938, LUT_AMPL_WIDTH),
		1579 => to_signed(4941, LUT_AMPL_WIDTH),
		1580 => to_signed(4945, LUT_AMPL_WIDTH),
		1581 => to_signed(4948, LUT_AMPL_WIDTH),
		1582 => to_signed(4951, LUT_AMPL_WIDTH),
		1583 => to_signed(4954, LUT_AMPL_WIDTH),
		1584 => to_signed(4957, LUT_AMPL_WIDTH),
		1585 => to_signed(4960, LUT_AMPL_WIDTH),
		1586 => to_signed(4963, LUT_AMPL_WIDTH),
		1587 => to_signed(4966, LUT_AMPL_WIDTH),
		1588 => to_signed(4969, LUT_AMPL_WIDTH),
		1589 => to_signed(4973, LUT_AMPL_WIDTH),
		1590 => to_signed(4976, LUT_AMPL_WIDTH),
		1591 => to_signed(4979, LUT_AMPL_WIDTH),
		1592 => to_signed(4982, LUT_AMPL_WIDTH),
		1593 => to_signed(4985, LUT_AMPL_WIDTH),
		1594 => to_signed(4988, LUT_AMPL_WIDTH),
		1595 => to_signed(4991, LUT_AMPL_WIDTH),
		1596 => to_signed(4994, LUT_AMPL_WIDTH),
		1597 => to_signed(4997, LUT_AMPL_WIDTH),
		1598 => to_signed(5000, LUT_AMPL_WIDTH),
		1599 => to_signed(5004, LUT_AMPL_WIDTH),
		1600 => to_signed(5007, LUT_AMPL_WIDTH),
		1601 => to_signed(5010, LUT_AMPL_WIDTH),
		1602 => to_signed(5013, LUT_AMPL_WIDTH),
		1603 => to_signed(5016, LUT_AMPL_WIDTH),
		1604 => to_signed(5019, LUT_AMPL_WIDTH),
		1605 => to_signed(5022, LUT_AMPL_WIDTH),
		1606 => to_signed(5025, LUT_AMPL_WIDTH),
		1607 => to_signed(5028, LUT_AMPL_WIDTH),
		1608 => to_signed(5032, LUT_AMPL_WIDTH),
		1609 => to_signed(5035, LUT_AMPL_WIDTH),
		1610 => to_signed(5038, LUT_AMPL_WIDTH),
		1611 => to_signed(5041, LUT_AMPL_WIDTH),
		1612 => to_signed(5044, LUT_AMPL_WIDTH),
		1613 => to_signed(5047, LUT_AMPL_WIDTH),
		1614 => to_signed(5050, LUT_AMPL_WIDTH),
		1615 => to_signed(5053, LUT_AMPL_WIDTH),
		1616 => to_signed(5056, LUT_AMPL_WIDTH),
		1617 => to_signed(5059, LUT_AMPL_WIDTH),
		1618 => to_signed(5063, LUT_AMPL_WIDTH),
		1619 => to_signed(5066, LUT_AMPL_WIDTH),
		1620 => to_signed(5069, LUT_AMPL_WIDTH),
		1621 => to_signed(5072, LUT_AMPL_WIDTH),
		1622 => to_signed(5075, LUT_AMPL_WIDTH),
		1623 => to_signed(5078, LUT_AMPL_WIDTH),
		1624 => to_signed(5081, LUT_AMPL_WIDTH),
		1625 => to_signed(5084, LUT_AMPL_WIDTH),
		1626 => to_signed(5087, LUT_AMPL_WIDTH),
		1627 => to_signed(5091, LUT_AMPL_WIDTH),
		1628 => to_signed(5094, LUT_AMPL_WIDTH),
		1629 => to_signed(5097, LUT_AMPL_WIDTH),
		1630 => to_signed(5100, LUT_AMPL_WIDTH),
		1631 => to_signed(5103, LUT_AMPL_WIDTH),
		1632 => to_signed(5106, LUT_AMPL_WIDTH),
		1633 => to_signed(5109, LUT_AMPL_WIDTH),
		1634 => to_signed(5112, LUT_AMPL_WIDTH),
		1635 => to_signed(5115, LUT_AMPL_WIDTH),
		1636 => to_signed(5118, LUT_AMPL_WIDTH),
		1637 => to_signed(5122, LUT_AMPL_WIDTH),
		1638 => to_signed(5125, LUT_AMPL_WIDTH),
		1639 => to_signed(5128, LUT_AMPL_WIDTH),
		1640 => to_signed(5131, LUT_AMPL_WIDTH),
		1641 => to_signed(5134, LUT_AMPL_WIDTH),
		1642 => to_signed(5137, LUT_AMPL_WIDTH),
		1643 => to_signed(5140, LUT_AMPL_WIDTH),
		1644 => to_signed(5143, LUT_AMPL_WIDTH),
		1645 => to_signed(5146, LUT_AMPL_WIDTH),
		1646 => to_signed(5149, LUT_AMPL_WIDTH),
		1647 => to_signed(5153, LUT_AMPL_WIDTH),
		1648 => to_signed(5156, LUT_AMPL_WIDTH),
		1649 => to_signed(5159, LUT_AMPL_WIDTH),
		1650 => to_signed(5162, LUT_AMPL_WIDTH),
		1651 => to_signed(5165, LUT_AMPL_WIDTH),
		1652 => to_signed(5168, LUT_AMPL_WIDTH),
		1653 => to_signed(5171, LUT_AMPL_WIDTH),
		1654 => to_signed(5174, LUT_AMPL_WIDTH),
		1655 => to_signed(5177, LUT_AMPL_WIDTH),
		1656 => to_signed(5180, LUT_AMPL_WIDTH),
		1657 => to_signed(5184, LUT_AMPL_WIDTH),
		1658 => to_signed(5187, LUT_AMPL_WIDTH),
		1659 => to_signed(5190, LUT_AMPL_WIDTH),
		1660 => to_signed(5193, LUT_AMPL_WIDTH),
		1661 => to_signed(5196, LUT_AMPL_WIDTH),
		1662 => to_signed(5199, LUT_AMPL_WIDTH),
		1663 => to_signed(5202, LUT_AMPL_WIDTH),
		1664 => to_signed(5205, LUT_AMPL_WIDTH),
		1665 => to_signed(5208, LUT_AMPL_WIDTH),
		1666 => to_signed(5212, LUT_AMPL_WIDTH),
		1667 => to_signed(5215, LUT_AMPL_WIDTH),
		1668 => to_signed(5218, LUT_AMPL_WIDTH),
		1669 => to_signed(5221, LUT_AMPL_WIDTH),
		1670 => to_signed(5224, LUT_AMPL_WIDTH),
		1671 => to_signed(5227, LUT_AMPL_WIDTH),
		1672 => to_signed(5230, LUT_AMPL_WIDTH),
		1673 => to_signed(5233, LUT_AMPL_WIDTH),
		1674 => to_signed(5236, LUT_AMPL_WIDTH),
		1675 => to_signed(5239, LUT_AMPL_WIDTH),
		1676 => to_signed(5243, LUT_AMPL_WIDTH),
		1677 => to_signed(5246, LUT_AMPL_WIDTH),
		1678 => to_signed(5249, LUT_AMPL_WIDTH),
		1679 => to_signed(5252, LUT_AMPL_WIDTH),
		1680 => to_signed(5255, LUT_AMPL_WIDTH),
		1681 => to_signed(5258, LUT_AMPL_WIDTH),
		1682 => to_signed(5261, LUT_AMPL_WIDTH),
		1683 => to_signed(5264, LUT_AMPL_WIDTH),
		1684 => to_signed(5267, LUT_AMPL_WIDTH),
		1685 => to_signed(5270, LUT_AMPL_WIDTH),
		1686 => to_signed(5274, LUT_AMPL_WIDTH),
		1687 => to_signed(5277, LUT_AMPL_WIDTH),
		1688 => to_signed(5280, LUT_AMPL_WIDTH),
		1689 => to_signed(5283, LUT_AMPL_WIDTH),
		1690 => to_signed(5286, LUT_AMPL_WIDTH),
		1691 => to_signed(5289, LUT_AMPL_WIDTH),
		1692 => to_signed(5292, LUT_AMPL_WIDTH),
		1693 => to_signed(5295, LUT_AMPL_WIDTH),
		1694 => to_signed(5298, LUT_AMPL_WIDTH),
		1695 => to_signed(5301, LUT_AMPL_WIDTH),
		1696 => to_signed(5305, LUT_AMPL_WIDTH),
		1697 => to_signed(5308, LUT_AMPL_WIDTH),
		1698 => to_signed(5311, LUT_AMPL_WIDTH),
		1699 => to_signed(5314, LUT_AMPL_WIDTH),
		1700 => to_signed(5317, LUT_AMPL_WIDTH),
		1701 => to_signed(5320, LUT_AMPL_WIDTH),
		1702 => to_signed(5323, LUT_AMPL_WIDTH),
		1703 => to_signed(5326, LUT_AMPL_WIDTH),
		1704 => to_signed(5329, LUT_AMPL_WIDTH),
		1705 => to_signed(5332, LUT_AMPL_WIDTH),
		1706 => to_signed(5336, LUT_AMPL_WIDTH),
		1707 => to_signed(5339, LUT_AMPL_WIDTH),
		1708 => to_signed(5342, LUT_AMPL_WIDTH),
		1709 => to_signed(5345, LUT_AMPL_WIDTH),
		1710 => to_signed(5348, LUT_AMPL_WIDTH),
		1711 => to_signed(5351, LUT_AMPL_WIDTH),
		1712 => to_signed(5354, LUT_AMPL_WIDTH),
		1713 => to_signed(5357, LUT_AMPL_WIDTH),
		1714 => to_signed(5360, LUT_AMPL_WIDTH),
		1715 => to_signed(5363, LUT_AMPL_WIDTH),
		1716 => to_signed(5367, LUT_AMPL_WIDTH),
		1717 => to_signed(5370, LUT_AMPL_WIDTH),
		1718 => to_signed(5373, LUT_AMPL_WIDTH),
		1719 => to_signed(5376, LUT_AMPL_WIDTH),
		1720 => to_signed(5379, LUT_AMPL_WIDTH),
		1721 => to_signed(5382, LUT_AMPL_WIDTH),
		1722 => to_signed(5385, LUT_AMPL_WIDTH),
		1723 => to_signed(5388, LUT_AMPL_WIDTH),
		1724 => to_signed(5391, LUT_AMPL_WIDTH),
		1725 => to_signed(5394, LUT_AMPL_WIDTH),
		1726 => to_signed(5398, LUT_AMPL_WIDTH),
		1727 => to_signed(5401, LUT_AMPL_WIDTH),
		1728 => to_signed(5404, LUT_AMPL_WIDTH),
		1729 => to_signed(5407, LUT_AMPL_WIDTH),
		1730 => to_signed(5410, LUT_AMPL_WIDTH),
		1731 => to_signed(5413, LUT_AMPL_WIDTH),
		1732 => to_signed(5416, LUT_AMPL_WIDTH),
		1733 => to_signed(5419, LUT_AMPL_WIDTH),
		1734 => to_signed(5422, LUT_AMPL_WIDTH),
		1735 => to_signed(5425, LUT_AMPL_WIDTH),
		1736 => to_signed(5428, LUT_AMPL_WIDTH),
		1737 => to_signed(5432, LUT_AMPL_WIDTH),
		1738 => to_signed(5435, LUT_AMPL_WIDTH),
		1739 => to_signed(5438, LUT_AMPL_WIDTH),
		1740 => to_signed(5441, LUT_AMPL_WIDTH),
		1741 => to_signed(5444, LUT_AMPL_WIDTH),
		1742 => to_signed(5447, LUT_AMPL_WIDTH),
		1743 => to_signed(5450, LUT_AMPL_WIDTH),
		1744 => to_signed(5453, LUT_AMPL_WIDTH),
		1745 => to_signed(5456, LUT_AMPL_WIDTH),
		1746 => to_signed(5459, LUT_AMPL_WIDTH),
		1747 => to_signed(5463, LUT_AMPL_WIDTH),
		1748 => to_signed(5466, LUT_AMPL_WIDTH),
		1749 => to_signed(5469, LUT_AMPL_WIDTH),
		1750 => to_signed(5472, LUT_AMPL_WIDTH),
		1751 => to_signed(5475, LUT_AMPL_WIDTH),
		1752 => to_signed(5478, LUT_AMPL_WIDTH),
		1753 => to_signed(5481, LUT_AMPL_WIDTH),
		1754 => to_signed(5484, LUT_AMPL_WIDTH),
		1755 => to_signed(5487, LUT_AMPL_WIDTH),
		1756 => to_signed(5490, LUT_AMPL_WIDTH),
		1757 => to_signed(5494, LUT_AMPL_WIDTH),
		1758 => to_signed(5497, LUT_AMPL_WIDTH),
		1759 => to_signed(5500, LUT_AMPL_WIDTH),
		1760 => to_signed(5503, LUT_AMPL_WIDTH),
		1761 => to_signed(5506, LUT_AMPL_WIDTH),
		1762 => to_signed(5509, LUT_AMPL_WIDTH),
		1763 => to_signed(5512, LUT_AMPL_WIDTH),
		1764 => to_signed(5515, LUT_AMPL_WIDTH),
		1765 => to_signed(5518, LUT_AMPL_WIDTH),
		1766 => to_signed(5521, LUT_AMPL_WIDTH),
		1767 => to_signed(5525, LUT_AMPL_WIDTH),
		1768 => to_signed(5528, LUT_AMPL_WIDTH),
		1769 => to_signed(5531, LUT_AMPL_WIDTH),
		1770 => to_signed(5534, LUT_AMPL_WIDTH),
		1771 => to_signed(5537, LUT_AMPL_WIDTH),
		1772 => to_signed(5540, LUT_AMPL_WIDTH),
		1773 => to_signed(5543, LUT_AMPL_WIDTH),
		1774 => to_signed(5546, LUT_AMPL_WIDTH),
		1775 => to_signed(5549, LUT_AMPL_WIDTH),
		1776 => to_signed(5552, LUT_AMPL_WIDTH),
		1777 => to_signed(5555, LUT_AMPL_WIDTH),
		1778 => to_signed(5559, LUT_AMPL_WIDTH),
		1779 => to_signed(5562, LUT_AMPL_WIDTH),
		1780 => to_signed(5565, LUT_AMPL_WIDTH),
		1781 => to_signed(5568, LUT_AMPL_WIDTH),
		1782 => to_signed(5571, LUT_AMPL_WIDTH),
		1783 => to_signed(5574, LUT_AMPL_WIDTH),
		1784 => to_signed(5577, LUT_AMPL_WIDTH),
		1785 => to_signed(5580, LUT_AMPL_WIDTH),
		1786 => to_signed(5583, LUT_AMPL_WIDTH),
		1787 => to_signed(5586, LUT_AMPL_WIDTH),
		1788 => to_signed(5590, LUT_AMPL_WIDTH),
		1789 => to_signed(5593, LUT_AMPL_WIDTH),
		1790 => to_signed(5596, LUT_AMPL_WIDTH),
		1791 => to_signed(5599, LUT_AMPL_WIDTH),
		1792 => to_signed(5602, LUT_AMPL_WIDTH),
		1793 => to_signed(5605, LUT_AMPL_WIDTH),
		1794 => to_signed(5608, LUT_AMPL_WIDTH),
		1795 => to_signed(5611, LUT_AMPL_WIDTH),
		1796 => to_signed(5614, LUT_AMPL_WIDTH),
		1797 => to_signed(5617, LUT_AMPL_WIDTH),
		1798 => to_signed(5620, LUT_AMPL_WIDTH),
		1799 => to_signed(5624, LUT_AMPL_WIDTH),
		1800 => to_signed(5627, LUT_AMPL_WIDTH),
		1801 => to_signed(5630, LUT_AMPL_WIDTH),
		1802 => to_signed(5633, LUT_AMPL_WIDTH),
		1803 => to_signed(5636, LUT_AMPL_WIDTH),
		1804 => to_signed(5639, LUT_AMPL_WIDTH),
		1805 => to_signed(5642, LUT_AMPL_WIDTH),
		1806 => to_signed(5645, LUT_AMPL_WIDTH),
		1807 => to_signed(5648, LUT_AMPL_WIDTH),
		1808 => to_signed(5651, LUT_AMPL_WIDTH),
		1809 => to_signed(5655, LUT_AMPL_WIDTH),
		1810 => to_signed(5658, LUT_AMPL_WIDTH),
		1811 => to_signed(5661, LUT_AMPL_WIDTH),
		1812 => to_signed(5664, LUT_AMPL_WIDTH),
		1813 => to_signed(5667, LUT_AMPL_WIDTH),
		1814 => to_signed(5670, LUT_AMPL_WIDTH),
		1815 => to_signed(5673, LUT_AMPL_WIDTH),
		1816 => to_signed(5676, LUT_AMPL_WIDTH),
		1817 => to_signed(5679, LUT_AMPL_WIDTH),
		1818 => to_signed(5682, LUT_AMPL_WIDTH),
		1819 => to_signed(5685, LUT_AMPL_WIDTH),
		1820 => to_signed(5689, LUT_AMPL_WIDTH),
		1821 => to_signed(5692, LUT_AMPL_WIDTH),
		1822 => to_signed(5695, LUT_AMPL_WIDTH),
		1823 => to_signed(5698, LUT_AMPL_WIDTH),
		1824 => to_signed(5701, LUT_AMPL_WIDTH),
		1825 => to_signed(5704, LUT_AMPL_WIDTH),
		1826 => to_signed(5707, LUT_AMPL_WIDTH),
		1827 => to_signed(5710, LUT_AMPL_WIDTH),
		1828 => to_signed(5713, LUT_AMPL_WIDTH),
		1829 => to_signed(5716, LUT_AMPL_WIDTH),
		1830 => to_signed(5719, LUT_AMPL_WIDTH),
		1831 => to_signed(5723, LUT_AMPL_WIDTH),
		1832 => to_signed(5726, LUT_AMPL_WIDTH),
		1833 => to_signed(5729, LUT_AMPL_WIDTH),
		1834 => to_signed(5732, LUT_AMPL_WIDTH),
		1835 => to_signed(5735, LUT_AMPL_WIDTH),
		1836 => to_signed(5738, LUT_AMPL_WIDTH),
		1837 => to_signed(5741, LUT_AMPL_WIDTH),
		1838 => to_signed(5744, LUT_AMPL_WIDTH),
		1839 => to_signed(5747, LUT_AMPL_WIDTH),
		1840 => to_signed(5750, LUT_AMPL_WIDTH),
		1841 => to_signed(5754, LUT_AMPL_WIDTH),
		1842 => to_signed(5757, LUT_AMPL_WIDTH),
		1843 => to_signed(5760, LUT_AMPL_WIDTH),
		1844 => to_signed(5763, LUT_AMPL_WIDTH),
		1845 => to_signed(5766, LUT_AMPL_WIDTH),
		1846 => to_signed(5769, LUT_AMPL_WIDTH),
		1847 => to_signed(5772, LUT_AMPL_WIDTH),
		1848 => to_signed(5775, LUT_AMPL_WIDTH),
		1849 => to_signed(5778, LUT_AMPL_WIDTH),
		1850 => to_signed(5781, LUT_AMPL_WIDTH),
		1851 => to_signed(5784, LUT_AMPL_WIDTH),
		1852 => to_signed(5788, LUT_AMPL_WIDTH),
		1853 => to_signed(5791, LUT_AMPL_WIDTH),
		1854 => to_signed(5794, LUT_AMPL_WIDTH),
		1855 => to_signed(5797, LUT_AMPL_WIDTH),
		1856 => to_signed(5800, LUT_AMPL_WIDTH),
		1857 => to_signed(5803, LUT_AMPL_WIDTH),
		1858 => to_signed(5806, LUT_AMPL_WIDTH),
		1859 => to_signed(5809, LUT_AMPL_WIDTH),
		1860 => to_signed(5812, LUT_AMPL_WIDTH),
		1861 => to_signed(5815, LUT_AMPL_WIDTH),
		1862 => to_signed(5818, LUT_AMPL_WIDTH),
		1863 => to_signed(5822, LUT_AMPL_WIDTH),
		1864 => to_signed(5825, LUT_AMPL_WIDTH),
		1865 => to_signed(5828, LUT_AMPL_WIDTH),
		1866 => to_signed(5831, LUT_AMPL_WIDTH),
		1867 => to_signed(5834, LUT_AMPL_WIDTH),
		1868 => to_signed(5837, LUT_AMPL_WIDTH),
		1869 => to_signed(5840, LUT_AMPL_WIDTH),
		1870 => to_signed(5843, LUT_AMPL_WIDTH),
		1871 => to_signed(5846, LUT_AMPL_WIDTH),
		1872 => to_signed(5849, LUT_AMPL_WIDTH),
		1873 => to_signed(5852, LUT_AMPL_WIDTH),
		1874 => to_signed(5856, LUT_AMPL_WIDTH),
		1875 => to_signed(5859, LUT_AMPL_WIDTH),
		1876 => to_signed(5862, LUT_AMPL_WIDTH),
		1877 => to_signed(5865, LUT_AMPL_WIDTH),
		1878 => to_signed(5868, LUT_AMPL_WIDTH),
		1879 => to_signed(5871, LUT_AMPL_WIDTH),
		1880 => to_signed(5874, LUT_AMPL_WIDTH),
		1881 => to_signed(5877, LUT_AMPL_WIDTH),
		1882 => to_signed(5880, LUT_AMPL_WIDTH),
		1883 => to_signed(5883, LUT_AMPL_WIDTH),
		1884 => to_signed(5886, LUT_AMPL_WIDTH),
		1885 => to_signed(5890, LUT_AMPL_WIDTH),
		1886 => to_signed(5893, LUT_AMPL_WIDTH),
		1887 => to_signed(5896, LUT_AMPL_WIDTH),
		1888 => to_signed(5899, LUT_AMPL_WIDTH),
		1889 => to_signed(5902, LUT_AMPL_WIDTH),
		1890 => to_signed(5905, LUT_AMPL_WIDTH),
		1891 => to_signed(5908, LUT_AMPL_WIDTH),
		1892 => to_signed(5911, LUT_AMPL_WIDTH),
		1893 => to_signed(5914, LUT_AMPL_WIDTH),
		1894 => to_signed(5917, LUT_AMPL_WIDTH),
		1895 => to_signed(5920, LUT_AMPL_WIDTH),
		1896 => to_signed(5924, LUT_AMPL_WIDTH),
		1897 => to_signed(5927, LUT_AMPL_WIDTH),
		1898 => to_signed(5930, LUT_AMPL_WIDTH),
		1899 => to_signed(5933, LUT_AMPL_WIDTH),
		1900 => to_signed(5936, LUT_AMPL_WIDTH),
		1901 => to_signed(5939, LUT_AMPL_WIDTH),
		1902 => to_signed(5942, LUT_AMPL_WIDTH),
		1903 => to_signed(5945, LUT_AMPL_WIDTH),
		1904 => to_signed(5948, LUT_AMPL_WIDTH),
		1905 => to_signed(5951, LUT_AMPL_WIDTH),
		1906 => to_signed(5954, LUT_AMPL_WIDTH),
		1907 => to_signed(5958, LUT_AMPL_WIDTH),
		1908 => to_signed(5961, LUT_AMPL_WIDTH),
		1909 => to_signed(5964, LUT_AMPL_WIDTH),
		1910 => to_signed(5967, LUT_AMPL_WIDTH),
		1911 => to_signed(5970, LUT_AMPL_WIDTH),
		1912 => to_signed(5973, LUT_AMPL_WIDTH),
		1913 => to_signed(5976, LUT_AMPL_WIDTH),
		1914 => to_signed(5979, LUT_AMPL_WIDTH),
		1915 => to_signed(5982, LUT_AMPL_WIDTH),
		1916 => to_signed(5985, LUT_AMPL_WIDTH),
		1917 => to_signed(5988, LUT_AMPL_WIDTH),
		1918 => to_signed(5991, LUT_AMPL_WIDTH),
		1919 => to_signed(5995, LUT_AMPL_WIDTH),
		1920 => to_signed(5998, LUT_AMPL_WIDTH),
		1921 => to_signed(6001, LUT_AMPL_WIDTH),
		1922 => to_signed(6004, LUT_AMPL_WIDTH),
		1923 => to_signed(6007, LUT_AMPL_WIDTH),
		1924 => to_signed(6010, LUT_AMPL_WIDTH),
		1925 => to_signed(6013, LUT_AMPL_WIDTH),
		1926 => to_signed(6016, LUT_AMPL_WIDTH),
		1927 => to_signed(6019, LUT_AMPL_WIDTH),
		1928 => to_signed(6022, LUT_AMPL_WIDTH),
		1929 => to_signed(6025, LUT_AMPL_WIDTH),
		1930 => to_signed(6029, LUT_AMPL_WIDTH),
		1931 => to_signed(6032, LUT_AMPL_WIDTH),
		1932 => to_signed(6035, LUT_AMPL_WIDTH),
		1933 => to_signed(6038, LUT_AMPL_WIDTH),
		1934 => to_signed(6041, LUT_AMPL_WIDTH),
		1935 => to_signed(6044, LUT_AMPL_WIDTH),
		1936 => to_signed(6047, LUT_AMPL_WIDTH),
		1937 => to_signed(6050, LUT_AMPL_WIDTH),
		1938 => to_signed(6053, LUT_AMPL_WIDTH),
		1939 => to_signed(6056, LUT_AMPL_WIDTH),
		1940 => to_signed(6059, LUT_AMPL_WIDTH),
		1941 => to_signed(6063, LUT_AMPL_WIDTH),
		1942 => to_signed(6066, LUT_AMPL_WIDTH),
		1943 => to_signed(6069, LUT_AMPL_WIDTH),
		1944 => to_signed(6072, LUT_AMPL_WIDTH),
		1945 => to_signed(6075, LUT_AMPL_WIDTH),
		1946 => to_signed(6078, LUT_AMPL_WIDTH),
		1947 => to_signed(6081, LUT_AMPL_WIDTH),
		1948 => to_signed(6084, LUT_AMPL_WIDTH),
		1949 => to_signed(6087, LUT_AMPL_WIDTH),
		1950 => to_signed(6090, LUT_AMPL_WIDTH),
		1951 => to_signed(6093, LUT_AMPL_WIDTH),
		1952 => to_signed(6096, LUT_AMPL_WIDTH),
		1953 => to_signed(6100, LUT_AMPL_WIDTH),
		1954 => to_signed(6103, LUT_AMPL_WIDTH),
		1955 => to_signed(6106, LUT_AMPL_WIDTH),
		1956 => to_signed(6109, LUT_AMPL_WIDTH),
		1957 => to_signed(6112, LUT_AMPL_WIDTH),
		1958 => to_signed(6115, LUT_AMPL_WIDTH),
		1959 => to_signed(6118, LUT_AMPL_WIDTH),
		1960 => to_signed(6121, LUT_AMPL_WIDTH),
		1961 => to_signed(6124, LUT_AMPL_WIDTH),
		1962 => to_signed(6127, LUT_AMPL_WIDTH),
		1963 => to_signed(6130, LUT_AMPL_WIDTH),
		1964 => to_signed(6134, LUT_AMPL_WIDTH),
		1965 => to_signed(6137, LUT_AMPL_WIDTH),
		1966 => to_signed(6140, LUT_AMPL_WIDTH),
		1967 => to_signed(6143, LUT_AMPL_WIDTH),
		1968 => to_signed(6146, LUT_AMPL_WIDTH),
		1969 => to_signed(6149, LUT_AMPL_WIDTH),
		1970 => to_signed(6152, LUT_AMPL_WIDTH),
		1971 => to_signed(6155, LUT_AMPL_WIDTH),
		1972 => to_signed(6158, LUT_AMPL_WIDTH),
		1973 => to_signed(6161, LUT_AMPL_WIDTH),
		1974 => to_signed(6164, LUT_AMPL_WIDTH),
		1975 => to_signed(6167, LUT_AMPL_WIDTH),
		1976 => to_signed(6171, LUT_AMPL_WIDTH),
		1977 => to_signed(6174, LUT_AMPL_WIDTH),
		1978 => to_signed(6177, LUT_AMPL_WIDTH),
		1979 => to_signed(6180, LUT_AMPL_WIDTH),
		1980 => to_signed(6183, LUT_AMPL_WIDTH),
		1981 => to_signed(6186, LUT_AMPL_WIDTH),
		1982 => to_signed(6189, LUT_AMPL_WIDTH),
		1983 => to_signed(6192, LUT_AMPL_WIDTH),
		1984 => to_signed(6195, LUT_AMPL_WIDTH),
		1985 => to_signed(6198, LUT_AMPL_WIDTH),
		1986 => to_signed(6201, LUT_AMPL_WIDTH),
		1987 => to_signed(6204, LUT_AMPL_WIDTH),
		1988 => to_signed(6208, LUT_AMPL_WIDTH),
		1989 => to_signed(6211, LUT_AMPL_WIDTH),
		1990 => to_signed(6214, LUT_AMPL_WIDTH),
		1991 => to_signed(6217, LUT_AMPL_WIDTH),
		1992 => to_signed(6220, LUT_AMPL_WIDTH),
		1993 => to_signed(6223, LUT_AMPL_WIDTH),
		1994 => to_signed(6226, LUT_AMPL_WIDTH),
		1995 => to_signed(6229, LUT_AMPL_WIDTH),
		1996 => to_signed(6232, LUT_AMPL_WIDTH),
		1997 => to_signed(6235, LUT_AMPL_WIDTH),
		1998 => to_signed(6238, LUT_AMPL_WIDTH),
		1999 => to_signed(6241, LUT_AMPL_WIDTH),
		2000 => to_signed(6245, LUT_AMPL_WIDTH),
		2001 => to_signed(6248, LUT_AMPL_WIDTH),
		2002 => to_signed(6251, LUT_AMPL_WIDTH),
		2003 => to_signed(6254, LUT_AMPL_WIDTH),
		2004 => to_signed(6257, LUT_AMPL_WIDTH),
		2005 => to_signed(6260, LUT_AMPL_WIDTH),
		2006 => to_signed(6263, LUT_AMPL_WIDTH),
		2007 => to_signed(6266, LUT_AMPL_WIDTH),
		2008 => to_signed(6269, LUT_AMPL_WIDTH),
		2009 => to_signed(6272, LUT_AMPL_WIDTH),
		2010 => to_signed(6275, LUT_AMPL_WIDTH),
		2011 => to_signed(6278, LUT_AMPL_WIDTH),
		2012 => to_signed(6282, LUT_AMPL_WIDTH),
		2013 => to_signed(6285, LUT_AMPL_WIDTH),
		2014 => to_signed(6288, LUT_AMPL_WIDTH),
		2015 => to_signed(6291, LUT_AMPL_WIDTH),
		2016 => to_signed(6294, LUT_AMPL_WIDTH),
		2017 => to_signed(6297, LUT_AMPL_WIDTH),
		2018 => to_signed(6300, LUT_AMPL_WIDTH),
		2019 => to_signed(6303, LUT_AMPL_WIDTH),
		2020 => to_signed(6306, LUT_AMPL_WIDTH),
		2021 => to_signed(6309, LUT_AMPL_WIDTH),
		2022 => to_signed(6312, LUT_AMPL_WIDTH),
		2023 => to_signed(6315, LUT_AMPL_WIDTH),
		2024 => to_signed(6319, LUT_AMPL_WIDTH),
		2025 => to_signed(6322, LUT_AMPL_WIDTH),
		2026 => to_signed(6325, LUT_AMPL_WIDTH),
		2027 => to_signed(6328, LUT_AMPL_WIDTH),
		2028 => to_signed(6331, LUT_AMPL_WIDTH),
		2029 => to_signed(6334, LUT_AMPL_WIDTH),
		2030 => to_signed(6337, LUT_AMPL_WIDTH),
		2031 => to_signed(6340, LUT_AMPL_WIDTH),
		2032 => to_signed(6343, LUT_AMPL_WIDTH),
		2033 => to_signed(6346, LUT_AMPL_WIDTH),
		2034 => to_signed(6349, LUT_AMPL_WIDTH),
		2035 => to_signed(6352, LUT_AMPL_WIDTH),
		2036 => to_signed(6356, LUT_AMPL_WIDTH),
		2037 => to_signed(6359, LUT_AMPL_WIDTH),
		2038 => to_signed(6362, LUT_AMPL_WIDTH),
		2039 => to_signed(6365, LUT_AMPL_WIDTH),
		2040 => to_signed(6368, LUT_AMPL_WIDTH),
		2041 => to_signed(6371, LUT_AMPL_WIDTH),
		2042 => to_signed(6374, LUT_AMPL_WIDTH),
		2043 => to_signed(6377, LUT_AMPL_WIDTH),
		2044 => to_signed(6380, LUT_AMPL_WIDTH),
		2045 => to_signed(6383, LUT_AMPL_WIDTH),
		2046 => to_signed(6386, LUT_AMPL_WIDTH),
		2047 => to_signed(6389, LUT_AMPL_WIDTH),
		2048 => to_signed(6393, LUT_AMPL_WIDTH),
		2049 => to_signed(6396, LUT_AMPL_WIDTH),
		2050 => to_signed(6399, LUT_AMPL_WIDTH),
		2051 => to_signed(6402, LUT_AMPL_WIDTH),
		2052 => to_signed(6405, LUT_AMPL_WIDTH),
		2053 => to_signed(6408, LUT_AMPL_WIDTH),
		2054 => to_signed(6411, LUT_AMPL_WIDTH),
		2055 => to_signed(6414, LUT_AMPL_WIDTH),
		2056 => to_signed(6417, LUT_AMPL_WIDTH),
		2057 => to_signed(6420, LUT_AMPL_WIDTH),
		2058 => to_signed(6423, LUT_AMPL_WIDTH),
		2059 => to_signed(6426, LUT_AMPL_WIDTH),
		2060 => to_signed(6429, LUT_AMPL_WIDTH),
		2061 => to_signed(6433, LUT_AMPL_WIDTH),
		2062 => to_signed(6436, LUT_AMPL_WIDTH),
		2063 => to_signed(6439, LUT_AMPL_WIDTH),
		2064 => to_signed(6442, LUT_AMPL_WIDTH),
		2065 => to_signed(6445, LUT_AMPL_WIDTH),
		2066 => to_signed(6448, LUT_AMPL_WIDTH),
		2067 => to_signed(6451, LUT_AMPL_WIDTH),
		2068 => to_signed(6454, LUT_AMPL_WIDTH),
		2069 => to_signed(6457, LUT_AMPL_WIDTH),
		2070 => to_signed(6460, LUT_AMPL_WIDTH),
		2071 => to_signed(6463, LUT_AMPL_WIDTH),
		2072 => to_signed(6466, LUT_AMPL_WIDTH),
		2073 => to_signed(6470, LUT_AMPL_WIDTH),
		2074 => to_signed(6473, LUT_AMPL_WIDTH),
		2075 => to_signed(6476, LUT_AMPL_WIDTH),
		2076 => to_signed(6479, LUT_AMPL_WIDTH),
		2077 => to_signed(6482, LUT_AMPL_WIDTH),
		2078 => to_signed(6485, LUT_AMPL_WIDTH),
		2079 => to_signed(6488, LUT_AMPL_WIDTH),
		2080 => to_signed(6491, LUT_AMPL_WIDTH),
		2081 => to_signed(6494, LUT_AMPL_WIDTH),
		2082 => to_signed(6497, LUT_AMPL_WIDTH),
		2083 => to_signed(6500, LUT_AMPL_WIDTH),
		2084 => to_signed(6503, LUT_AMPL_WIDTH),
		2085 => to_signed(6506, LUT_AMPL_WIDTH),
		2086 => to_signed(6510, LUT_AMPL_WIDTH),
		2087 => to_signed(6513, LUT_AMPL_WIDTH),
		2088 => to_signed(6516, LUT_AMPL_WIDTH),
		2089 => to_signed(6519, LUT_AMPL_WIDTH),
		2090 => to_signed(6522, LUT_AMPL_WIDTH),
		2091 => to_signed(6525, LUT_AMPL_WIDTH),
		2092 => to_signed(6528, LUT_AMPL_WIDTH),
		2093 => to_signed(6531, LUT_AMPL_WIDTH),
		2094 => to_signed(6534, LUT_AMPL_WIDTH),
		2095 => to_signed(6537, LUT_AMPL_WIDTH),
		2096 => to_signed(6540, LUT_AMPL_WIDTH),
		2097 => to_signed(6543, LUT_AMPL_WIDTH),
		2098 => to_signed(6547, LUT_AMPL_WIDTH),
		2099 => to_signed(6550, LUT_AMPL_WIDTH),
		2100 => to_signed(6553, LUT_AMPL_WIDTH),
		2101 => to_signed(6556, LUT_AMPL_WIDTH),
		2102 => to_signed(6559, LUT_AMPL_WIDTH),
		2103 => to_signed(6562, LUT_AMPL_WIDTH),
		2104 => to_signed(6565, LUT_AMPL_WIDTH),
		2105 => to_signed(6568, LUT_AMPL_WIDTH),
		2106 => to_signed(6571, LUT_AMPL_WIDTH),
		2107 => to_signed(6574, LUT_AMPL_WIDTH),
		2108 => to_signed(6577, LUT_AMPL_WIDTH),
		2109 => to_signed(6580, LUT_AMPL_WIDTH),
		2110 => to_signed(6583, LUT_AMPL_WIDTH),
		2111 => to_signed(6587, LUT_AMPL_WIDTH),
		2112 => to_signed(6590, LUT_AMPL_WIDTH),
		2113 => to_signed(6593, LUT_AMPL_WIDTH),
		2114 => to_signed(6596, LUT_AMPL_WIDTH),
		2115 => to_signed(6599, LUT_AMPL_WIDTH),
		2116 => to_signed(6602, LUT_AMPL_WIDTH),
		2117 => to_signed(6605, LUT_AMPL_WIDTH),
		2118 => to_signed(6608, LUT_AMPL_WIDTH),
		2119 => to_signed(6611, LUT_AMPL_WIDTH),
		2120 => to_signed(6614, LUT_AMPL_WIDTH),
		2121 => to_signed(6617, LUT_AMPL_WIDTH),
		2122 => to_signed(6620, LUT_AMPL_WIDTH),
		2123 => to_signed(6623, LUT_AMPL_WIDTH),
		2124 => to_signed(6627, LUT_AMPL_WIDTH),
		2125 => to_signed(6630, LUT_AMPL_WIDTH),
		2126 => to_signed(6633, LUT_AMPL_WIDTH),
		2127 => to_signed(6636, LUT_AMPL_WIDTH),
		2128 => to_signed(6639, LUT_AMPL_WIDTH),
		2129 => to_signed(6642, LUT_AMPL_WIDTH),
		2130 => to_signed(6645, LUT_AMPL_WIDTH),
		2131 => to_signed(6648, LUT_AMPL_WIDTH),
		2132 => to_signed(6651, LUT_AMPL_WIDTH),
		2133 => to_signed(6654, LUT_AMPL_WIDTH),
		2134 => to_signed(6657, LUT_AMPL_WIDTH),
		2135 => to_signed(6660, LUT_AMPL_WIDTH),
		2136 => to_signed(6663, LUT_AMPL_WIDTH),
		2137 => to_signed(6667, LUT_AMPL_WIDTH),
		2138 => to_signed(6670, LUT_AMPL_WIDTH),
		2139 => to_signed(6673, LUT_AMPL_WIDTH),
		2140 => to_signed(6676, LUT_AMPL_WIDTH),
		2141 => to_signed(6679, LUT_AMPL_WIDTH),
		2142 => to_signed(6682, LUT_AMPL_WIDTH),
		2143 => to_signed(6685, LUT_AMPL_WIDTH),
		2144 => to_signed(6688, LUT_AMPL_WIDTH),
		2145 => to_signed(6691, LUT_AMPL_WIDTH),
		2146 => to_signed(6694, LUT_AMPL_WIDTH),
		2147 => to_signed(6697, LUT_AMPL_WIDTH),
		2148 => to_signed(6700, LUT_AMPL_WIDTH),
		2149 => to_signed(6703, LUT_AMPL_WIDTH),
		2150 => to_signed(6706, LUT_AMPL_WIDTH),
		2151 => to_signed(6710, LUT_AMPL_WIDTH),
		2152 => to_signed(6713, LUT_AMPL_WIDTH),
		2153 => to_signed(6716, LUT_AMPL_WIDTH),
		2154 => to_signed(6719, LUT_AMPL_WIDTH),
		2155 => to_signed(6722, LUT_AMPL_WIDTH),
		2156 => to_signed(6725, LUT_AMPL_WIDTH),
		2157 => to_signed(6728, LUT_AMPL_WIDTH),
		2158 => to_signed(6731, LUT_AMPL_WIDTH),
		2159 => to_signed(6734, LUT_AMPL_WIDTH),
		2160 => to_signed(6737, LUT_AMPL_WIDTH),
		2161 => to_signed(6740, LUT_AMPL_WIDTH),
		2162 => to_signed(6743, LUT_AMPL_WIDTH),
		2163 => to_signed(6746, LUT_AMPL_WIDTH),
		2164 => to_signed(6750, LUT_AMPL_WIDTH),
		2165 => to_signed(6753, LUT_AMPL_WIDTH),
		2166 => to_signed(6756, LUT_AMPL_WIDTH),
		2167 => to_signed(6759, LUT_AMPL_WIDTH),
		2168 => to_signed(6762, LUT_AMPL_WIDTH),
		2169 => to_signed(6765, LUT_AMPL_WIDTH),
		2170 => to_signed(6768, LUT_AMPL_WIDTH),
		2171 => to_signed(6771, LUT_AMPL_WIDTH),
		2172 => to_signed(6774, LUT_AMPL_WIDTH),
		2173 => to_signed(6777, LUT_AMPL_WIDTH),
		2174 => to_signed(6780, LUT_AMPL_WIDTH),
		2175 => to_signed(6783, LUT_AMPL_WIDTH),
		2176 => to_signed(6786, LUT_AMPL_WIDTH),
		2177 => to_signed(6789, LUT_AMPL_WIDTH),
		2178 => to_signed(6793, LUT_AMPL_WIDTH),
		2179 => to_signed(6796, LUT_AMPL_WIDTH),
		2180 => to_signed(6799, LUT_AMPL_WIDTH),
		2181 => to_signed(6802, LUT_AMPL_WIDTH),
		2182 => to_signed(6805, LUT_AMPL_WIDTH),
		2183 => to_signed(6808, LUT_AMPL_WIDTH),
		2184 => to_signed(6811, LUT_AMPL_WIDTH),
		2185 => to_signed(6814, LUT_AMPL_WIDTH),
		2186 => to_signed(6817, LUT_AMPL_WIDTH),
		2187 => to_signed(6820, LUT_AMPL_WIDTH),
		2188 => to_signed(6823, LUT_AMPL_WIDTH),
		2189 => to_signed(6826, LUT_AMPL_WIDTH),
		2190 => to_signed(6829, LUT_AMPL_WIDTH),
		2191 => to_signed(6833, LUT_AMPL_WIDTH),
		2192 => to_signed(6836, LUT_AMPL_WIDTH),
		2193 => to_signed(6839, LUT_AMPL_WIDTH),
		2194 => to_signed(6842, LUT_AMPL_WIDTH),
		2195 => to_signed(6845, LUT_AMPL_WIDTH),
		2196 => to_signed(6848, LUT_AMPL_WIDTH),
		2197 => to_signed(6851, LUT_AMPL_WIDTH),
		2198 => to_signed(6854, LUT_AMPL_WIDTH),
		2199 => to_signed(6857, LUT_AMPL_WIDTH),
		2200 => to_signed(6860, LUT_AMPL_WIDTH),
		2201 => to_signed(6863, LUT_AMPL_WIDTH),
		2202 => to_signed(6866, LUT_AMPL_WIDTH),
		2203 => to_signed(6869, LUT_AMPL_WIDTH),
		2204 => to_signed(6872, LUT_AMPL_WIDTH),
		2205 => to_signed(6876, LUT_AMPL_WIDTH),
		2206 => to_signed(6879, LUT_AMPL_WIDTH),
		2207 => to_signed(6882, LUT_AMPL_WIDTH),
		2208 => to_signed(6885, LUT_AMPL_WIDTH),
		2209 => to_signed(6888, LUT_AMPL_WIDTH),
		2210 => to_signed(6891, LUT_AMPL_WIDTH),
		2211 => to_signed(6894, LUT_AMPL_WIDTH),
		2212 => to_signed(6897, LUT_AMPL_WIDTH),
		2213 => to_signed(6900, LUT_AMPL_WIDTH),
		2214 => to_signed(6903, LUT_AMPL_WIDTH),
		2215 => to_signed(6906, LUT_AMPL_WIDTH),
		2216 => to_signed(6909, LUT_AMPL_WIDTH),
		2217 => to_signed(6912, LUT_AMPL_WIDTH),
		2218 => to_signed(6915, LUT_AMPL_WIDTH),
		2219 => to_signed(6919, LUT_AMPL_WIDTH),
		2220 => to_signed(6922, LUT_AMPL_WIDTH),
		2221 => to_signed(6925, LUT_AMPL_WIDTH),
		2222 => to_signed(6928, LUT_AMPL_WIDTH),
		2223 => to_signed(6931, LUT_AMPL_WIDTH),
		2224 => to_signed(6934, LUT_AMPL_WIDTH),
		2225 => to_signed(6937, LUT_AMPL_WIDTH),
		2226 => to_signed(6940, LUT_AMPL_WIDTH),
		2227 => to_signed(6943, LUT_AMPL_WIDTH),
		2228 => to_signed(6946, LUT_AMPL_WIDTH),
		2229 => to_signed(6949, LUT_AMPL_WIDTH),
		2230 => to_signed(6952, LUT_AMPL_WIDTH),
		2231 => to_signed(6955, LUT_AMPL_WIDTH),
		2232 => to_signed(6958, LUT_AMPL_WIDTH),
		2233 => to_signed(6961, LUT_AMPL_WIDTH),
		2234 => to_signed(6965, LUT_AMPL_WIDTH),
		2235 => to_signed(6968, LUT_AMPL_WIDTH),
		2236 => to_signed(6971, LUT_AMPL_WIDTH),
		2237 => to_signed(6974, LUT_AMPL_WIDTH),
		2238 => to_signed(6977, LUT_AMPL_WIDTH),
		2239 => to_signed(6980, LUT_AMPL_WIDTH),
		2240 => to_signed(6983, LUT_AMPL_WIDTH),
		2241 => to_signed(6986, LUT_AMPL_WIDTH),
		2242 => to_signed(6989, LUT_AMPL_WIDTH),
		2243 => to_signed(6992, LUT_AMPL_WIDTH),
		2244 => to_signed(6995, LUT_AMPL_WIDTH),
		2245 => to_signed(6998, LUT_AMPL_WIDTH),
		2246 => to_signed(7001, LUT_AMPL_WIDTH),
		2247 => to_signed(7004, LUT_AMPL_WIDTH),
		2248 => to_signed(7008, LUT_AMPL_WIDTH),
		2249 => to_signed(7011, LUT_AMPL_WIDTH),
		2250 => to_signed(7014, LUT_AMPL_WIDTH),
		2251 => to_signed(7017, LUT_AMPL_WIDTH),
		2252 => to_signed(7020, LUT_AMPL_WIDTH),
		2253 => to_signed(7023, LUT_AMPL_WIDTH),
		2254 => to_signed(7026, LUT_AMPL_WIDTH),
		2255 => to_signed(7029, LUT_AMPL_WIDTH),
		2256 => to_signed(7032, LUT_AMPL_WIDTH),
		2257 => to_signed(7035, LUT_AMPL_WIDTH),
		2258 => to_signed(7038, LUT_AMPL_WIDTH),
		2259 => to_signed(7041, LUT_AMPL_WIDTH),
		2260 => to_signed(7044, LUT_AMPL_WIDTH),
		2261 => to_signed(7047, LUT_AMPL_WIDTH),
		2262 => to_signed(7050, LUT_AMPL_WIDTH),
		2263 => to_signed(7054, LUT_AMPL_WIDTH),
		2264 => to_signed(7057, LUT_AMPL_WIDTH),
		2265 => to_signed(7060, LUT_AMPL_WIDTH),
		2266 => to_signed(7063, LUT_AMPL_WIDTH),
		2267 => to_signed(7066, LUT_AMPL_WIDTH),
		2268 => to_signed(7069, LUT_AMPL_WIDTH),
		2269 => to_signed(7072, LUT_AMPL_WIDTH),
		2270 => to_signed(7075, LUT_AMPL_WIDTH),
		2271 => to_signed(7078, LUT_AMPL_WIDTH),
		2272 => to_signed(7081, LUT_AMPL_WIDTH),
		2273 => to_signed(7084, LUT_AMPL_WIDTH),
		2274 => to_signed(7087, LUT_AMPL_WIDTH),
		2275 => to_signed(7090, LUT_AMPL_WIDTH),
		2276 => to_signed(7093, LUT_AMPL_WIDTH),
		2277 => to_signed(7097, LUT_AMPL_WIDTH),
		2278 => to_signed(7100, LUT_AMPL_WIDTH),
		2279 => to_signed(7103, LUT_AMPL_WIDTH),
		2280 => to_signed(7106, LUT_AMPL_WIDTH),
		2281 => to_signed(7109, LUT_AMPL_WIDTH),
		2282 => to_signed(7112, LUT_AMPL_WIDTH),
		2283 => to_signed(7115, LUT_AMPL_WIDTH),
		2284 => to_signed(7118, LUT_AMPL_WIDTH),
		2285 => to_signed(7121, LUT_AMPL_WIDTH),
		2286 => to_signed(7124, LUT_AMPL_WIDTH),
		2287 => to_signed(7127, LUT_AMPL_WIDTH),
		2288 => to_signed(7130, LUT_AMPL_WIDTH),
		2289 => to_signed(7133, LUT_AMPL_WIDTH),
		2290 => to_signed(7136, LUT_AMPL_WIDTH),
		2291 => to_signed(7139, LUT_AMPL_WIDTH),
		2292 => to_signed(7143, LUT_AMPL_WIDTH),
		2293 => to_signed(7146, LUT_AMPL_WIDTH),
		2294 => to_signed(7149, LUT_AMPL_WIDTH),
		2295 => to_signed(7152, LUT_AMPL_WIDTH),
		2296 => to_signed(7155, LUT_AMPL_WIDTH),
		2297 => to_signed(7158, LUT_AMPL_WIDTH),
		2298 => to_signed(7161, LUT_AMPL_WIDTH),
		2299 => to_signed(7164, LUT_AMPL_WIDTH),
		2300 => to_signed(7167, LUT_AMPL_WIDTH),
		2301 => to_signed(7170, LUT_AMPL_WIDTH),
		2302 => to_signed(7173, LUT_AMPL_WIDTH),
		2303 => to_signed(7176, LUT_AMPL_WIDTH),
		2304 => to_signed(7179, LUT_AMPL_WIDTH),
		2305 => to_signed(7182, LUT_AMPL_WIDTH),
		2306 => to_signed(7185, LUT_AMPL_WIDTH),
		2307 => to_signed(7188, LUT_AMPL_WIDTH),
		2308 => to_signed(7192, LUT_AMPL_WIDTH),
		2309 => to_signed(7195, LUT_AMPL_WIDTH),
		2310 => to_signed(7198, LUT_AMPL_WIDTH),
		2311 => to_signed(7201, LUT_AMPL_WIDTH),
		2312 => to_signed(7204, LUT_AMPL_WIDTH),
		2313 => to_signed(7207, LUT_AMPL_WIDTH),
		2314 => to_signed(7210, LUT_AMPL_WIDTH),
		2315 => to_signed(7213, LUT_AMPL_WIDTH),
		2316 => to_signed(7216, LUT_AMPL_WIDTH),
		2317 => to_signed(7219, LUT_AMPL_WIDTH),
		2318 => to_signed(7222, LUT_AMPL_WIDTH),
		2319 => to_signed(7225, LUT_AMPL_WIDTH),
		2320 => to_signed(7228, LUT_AMPL_WIDTH),
		2321 => to_signed(7231, LUT_AMPL_WIDTH),
		2322 => to_signed(7234, LUT_AMPL_WIDTH),
		2323 => to_signed(7238, LUT_AMPL_WIDTH),
		2324 => to_signed(7241, LUT_AMPL_WIDTH),
		2325 => to_signed(7244, LUT_AMPL_WIDTH),
		2326 => to_signed(7247, LUT_AMPL_WIDTH),
		2327 => to_signed(7250, LUT_AMPL_WIDTH),
		2328 => to_signed(7253, LUT_AMPL_WIDTH),
		2329 => to_signed(7256, LUT_AMPL_WIDTH),
		2330 => to_signed(7259, LUT_AMPL_WIDTH),
		2331 => to_signed(7262, LUT_AMPL_WIDTH),
		2332 => to_signed(7265, LUT_AMPL_WIDTH),
		2333 => to_signed(7268, LUT_AMPL_WIDTH),
		2334 => to_signed(7271, LUT_AMPL_WIDTH),
		2335 => to_signed(7274, LUT_AMPL_WIDTH),
		2336 => to_signed(7277, LUT_AMPL_WIDTH),
		2337 => to_signed(7280, LUT_AMPL_WIDTH),
		2338 => to_signed(7283, LUT_AMPL_WIDTH),
		2339 => to_signed(7287, LUT_AMPL_WIDTH),
		2340 => to_signed(7290, LUT_AMPL_WIDTH),
		2341 => to_signed(7293, LUT_AMPL_WIDTH),
		2342 => to_signed(7296, LUT_AMPL_WIDTH),
		2343 => to_signed(7299, LUT_AMPL_WIDTH),
		2344 => to_signed(7302, LUT_AMPL_WIDTH),
		2345 => to_signed(7305, LUT_AMPL_WIDTH),
		2346 => to_signed(7308, LUT_AMPL_WIDTH),
		2347 => to_signed(7311, LUT_AMPL_WIDTH),
		2348 => to_signed(7314, LUT_AMPL_WIDTH),
		2349 => to_signed(7317, LUT_AMPL_WIDTH),
		2350 => to_signed(7320, LUT_AMPL_WIDTH),
		2351 => to_signed(7323, LUT_AMPL_WIDTH),
		2352 => to_signed(7326, LUT_AMPL_WIDTH),
		2353 => to_signed(7329, LUT_AMPL_WIDTH),
		2354 => to_signed(7332, LUT_AMPL_WIDTH),
		2355 => to_signed(7336, LUT_AMPL_WIDTH),
		2356 => to_signed(7339, LUT_AMPL_WIDTH),
		2357 => to_signed(7342, LUT_AMPL_WIDTH),
		2358 => to_signed(7345, LUT_AMPL_WIDTH),
		2359 => to_signed(7348, LUT_AMPL_WIDTH),
		2360 => to_signed(7351, LUT_AMPL_WIDTH),
		2361 => to_signed(7354, LUT_AMPL_WIDTH),
		2362 => to_signed(7357, LUT_AMPL_WIDTH),
		2363 => to_signed(7360, LUT_AMPL_WIDTH),
		2364 => to_signed(7363, LUT_AMPL_WIDTH),
		2365 => to_signed(7366, LUT_AMPL_WIDTH),
		2366 => to_signed(7369, LUT_AMPL_WIDTH),
		2367 => to_signed(7372, LUT_AMPL_WIDTH),
		2368 => to_signed(7375, LUT_AMPL_WIDTH),
		2369 => to_signed(7378, LUT_AMPL_WIDTH),
		2370 => to_signed(7381, LUT_AMPL_WIDTH),
		2371 => to_signed(7385, LUT_AMPL_WIDTH),
		2372 => to_signed(7388, LUT_AMPL_WIDTH),
		2373 => to_signed(7391, LUT_AMPL_WIDTH),
		2374 => to_signed(7394, LUT_AMPL_WIDTH),
		2375 => to_signed(7397, LUT_AMPL_WIDTH),
		2376 => to_signed(7400, LUT_AMPL_WIDTH),
		2377 => to_signed(7403, LUT_AMPL_WIDTH),
		2378 => to_signed(7406, LUT_AMPL_WIDTH),
		2379 => to_signed(7409, LUT_AMPL_WIDTH),
		2380 => to_signed(7412, LUT_AMPL_WIDTH),
		2381 => to_signed(7415, LUT_AMPL_WIDTH),
		2382 => to_signed(7418, LUT_AMPL_WIDTH),
		2383 => to_signed(7421, LUT_AMPL_WIDTH),
		2384 => to_signed(7424, LUT_AMPL_WIDTH),
		2385 => to_signed(7427, LUT_AMPL_WIDTH),
		2386 => to_signed(7430, LUT_AMPL_WIDTH),
		2387 => to_signed(7433, LUT_AMPL_WIDTH),
		2388 => to_signed(7437, LUT_AMPL_WIDTH),
		2389 => to_signed(7440, LUT_AMPL_WIDTH),
		2390 => to_signed(7443, LUT_AMPL_WIDTH),
		2391 => to_signed(7446, LUT_AMPL_WIDTH),
		2392 => to_signed(7449, LUT_AMPL_WIDTH),
		2393 => to_signed(7452, LUT_AMPL_WIDTH),
		2394 => to_signed(7455, LUT_AMPL_WIDTH),
		2395 => to_signed(7458, LUT_AMPL_WIDTH),
		2396 => to_signed(7461, LUT_AMPL_WIDTH),
		2397 => to_signed(7464, LUT_AMPL_WIDTH),
		2398 => to_signed(7467, LUT_AMPL_WIDTH),
		2399 => to_signed(7470, LUT_AMPL_WIDTH),
		2400 => to_signed(7473, LUT_AMPL_WIDTH),
		2401 => to_signed(7476, LUT_AMPL_WIDTH),
		2402 => to_signed(7479, LUT_AMPL_WIDTH),
		2403 => to_signed(7482, LUT_AMPL_WIDTH),
		2404 => to_signed(7485, LUT_AMPL_WIDTH),
		2405 => to_signed(7489, LUT_AMPL_WIDTH),
		2406 => to_signed(7492, LUT_AMPL_WIDTH),
		2407 => to_signed(7495, LUT_AMPL_WIDTH),
		2408 => to_signed(7498, LUT_AMPL_WIDTH),
		2409 => to_signed(7501, LUT_AMPL_WIDTH),
		2410 => to_signed(7504, LUT_AMPL_WIDTH),
		2411 => to_signed(7507, LUT_AMPL_WIDTH),
		2412 => to_signed(7510, LUT_AMPL_WIDTH),
		2413 => to_signed(7513, LUT_AMPL_WIDTH),
		2414 => to_signed(7516, LUT_AMPL_WIDTH),
		2415 => to_signed(7519, LUT_AMPL_WIDTH),
		2416 => to_signed(7522, LUT_AMPL_WIDTH),
		2417 => to_signed(7525, LUT_AMPL_WIDTH),
		2418 => to_signed(7528, LUT_AMPL_WIDTH),
		2419 => to_signed(7531, LUT_AMPL_WIDTH),
		2420 => to_signed(7534, LUT_AMPL_WIDTH),
		2421 => to_signed(7537, LUT_AMPL_WIDTH),
		2422 => to_signed(7541, LUT_AMPL_WIDTH),
		2423 => to_signed(7544, LUT_AMPL_WIDTH),
		2424 => to_signed(7547, LUT_AMPL_WIDTH),
		2425 => to_signed(7550, LUT_AMPL_WIDTH),
		2426 => to_signed(7553, LUT_AMPL_WIDTH),
		2427 => to_signed(7556, LUT_AMPL_WIDTH),
		2428 => to_signed(7559, LUT_AMPL_WIDTH),
		2429 => to_signed(7562, LUT_AMPL_WIDTH),
		2430 => to_signed(7565, LUT_AMPL_WIDTH),
		2431 => to_signed(7568, LUT_AMPL_WIDTH),
		2432 => to_signed(7571, LUT_AMPL_WIDTH),
		2433 => to_signed(7574, LUT_AMPL_WIDTH),
		2434 => to_signed(7577, LUT_AMPL_WIDTH),
		2435 => to_signed(7580, LUT_AMPL_WIDTH),
		2436 => to_signed(7583, LUT_AMPL_WIDTH),
		2437 => to_signed(7586, LUT_AMPL_WIDTH),
		2438 => to_signed(7589, LUT_AMPL_WIDTH),
		2439 => to_signed(7592, LUT_AMPL_WIDTH),
		2440 => to_signed(7596, LUT_AMPL_WIDTH),
		2441 => to_signed(7599, LUT_AMPL_WIDTH),
		2442 => to_signed(7602, LUT_AMPL_WIDTH),
		2443 => to_signed(7605, LUT_AMPL_WIDTH),
		2444 => to_signed(7608, LUT_AMPL_WIDTH),
		2445 => to_signed(7611, LUT_AMPL_WIDTH),
		2446 => to_signed(7614, LUT_AMPL_WIDTH),
		2447 => to_signed(7617, LUT_AMPL_WIDTH),
		2448 => to_signed(7620, LUT_AMPL_WIDTH),
		2449 => to_signed(7623, LUT_AMPL_WIDTH),
		2450 => to_signed(7626, LUT_AMPL_WIDTH),
		2451 => to_signed(7629, LUT_AMPL_WIDTH),
		2452 => to_signed(7632, LUT_AMPL_WIDTH),
		2453 => to_signed(7635, LUT_AMPL_WIDTH),
		2454 => to_signed(7638, LUT_AMPL_WIDTH),
		2455 => to_signed(7641, LUT_AMPL_WIDTH),
		2456 => to_signed(7644, LUT_AMPL_WIDTH),
		2457 => to_signed(7647, LUT_AMPL_WIDTH),
		2458 => to_signed(7651, LUT_AMPL_WIDTH),
		2459 => to_signed(7654, LUT_AMPL_WIDTH),
		2460 => to_signed(7657, LUT_AMPL_WIDTH),
		2461 => to_signed(7660, LUT_AMPL_WIDTH),
		2462 => to_signed(7663, LUT_AMPL_WIDTH),
		2463 => to_signed(7666, LUT_AMPL_WIDTH),
		2464 => to_signed(7669, LUT_AMPL_WIDTH),
		2465 => to_signed(7672, LUT_AMPL_WIDTH),
		2466 => to_signed(7675, LUT_AMPL_WIDTH),
		2467 => to_signed(7678, LUT_AMPL_WIDTH),
		2468 => to_signed(7681, LUT_AMPL_WIDTH),
		2469 => to_signed(7684, LUT_AMPL_WIDTH),
		2470 => to_signed(7687, LUT_AMPL_WIDTH),
		2471 => to_signed(7690, LUT_AMPL_WIDTH),
		2472 => to_signed(7693, LUT_AMPL_WIDTH),
		2473 => to_signed(7696, LUT_AMPL_WIDTH),
		2474 => to_signed(7699, LUT_AMPL_WIDTH),
		2475 => to_signed(7702, LUT_AMPL_WIDTH),
		2476 => to_signed(7705, LUT_AMPL_WIDTH),
		2477 => to_signed(7709, LUT_AMPL_WIDTH),
		2478 => to_signed(7712, LUT_AMPL_WIDTH),
		2479 => to_signed(7715, LUT_AMPL_WIDTH),
		2480 => to_signed(7718, LUT_AMPL_WIDTH),
		2481 => to_signed(7721, LUT_AMPL_WIDTH),
		2482 => to_signed(7724, LUT_AMPL_WIDTH),
		2483 => to_signed(7727, LUT_AMPL_WIDTH),
		2484 => to_signed(7730, LUT_AMPL_WIDTH),
		2485 => to_signed(7733, LUT_AMPL_WIDTH),
		2486 => to_signed(7736, LUT_AMPL_WIDTH),
		2487 => to_signed(7739, LUT_AMPL_WIDTH),
		2488 => to_signed(7742, LUT_AMPL_WIDTH),
		2489 => to_signed(7745, LUT_AMPL_WIDTH),
		2490 => to_signed(7748, LUT_AMPL_WIDTH),
		2491 => to_signed(7751, LUT_AMPL_WIDTH),
		2492 => to_signed(7754, LUT_AMPL_WIDTH),
		2493 => to_signed(7757, LUT_AMPL_WIDTH),
		2494 => to_signed(7760, LUT_AMPL_WIDTH),
		2495 => to_signed(7764, LUT_AMPL_WIDTH),
		2496 => to_signed(7767, LUT_AMPL_WIDTH),
		2497 => to_signed(7770, LUT_AMPL_WIDTH),
		2498 => to_signed(7773, LUT_AMPL_WIDTH),
		2499 => to_signed(7776, LUT_AMPL_WIDTH),
		2500 => to_signed(7779, LUT_AMPL_WIDTH),
		2501 => to_signed(7782, LUT_AMPL_WIDTH),
		2502 => to_signed(7785, LUT_AMPL_WIDTH),
		2503 => to_signed(7788, LUT_AMPL_WIDTH),
		2504 => to_signed(7791, LUT_AMPL_WIDTH),
		2505 => to_signed(7794, LUT_AMPL_WIDTH),
		2506 => to_signed(7797, LUT_AMPL_WIDTH),
		2507 => to_signed(7800, LUT_AMPL_WIDTH),
		2508 => to_signed(7803, LUT_AMPL_WIDTH),
		2509 => to_signed(7806, LUT_AMPL_WIDTH),
		2510 => to_signed(7809, LUT_AMPL_WIDTH),
		2511 => to_signed(7812, LUT_AMPL_WIDTH),
		2512 => to_signed(7815, LUT_AMPL_WIDTH),
		2513 => to_signed(7818, LUT_AMPL_WIDTH),
		2514 => to_signed(7821, LUT_AMPL_WIDTH),
		2515 => to_signed(7825, LUT_AMPL_WIDTH),
		2516 => to_signed(7828, LUT_AMPL_WIDTH),
		2517 => to_signed(7831, LUT_AMPL_WIDTH),
		2518 => to_signed(7834, LUT_AMPL_WIDTH),
		2519 => to_signed(7837, LUT_AMPL_WIDTH),
		2520 => to_signed(7840, LUT_AMPL_WIDTH),
		2521 => to_signed(7843, LUT_AMPL_WIDTH),
		2522 => to_signed(7846, LUT_AMPL_WIDTH),
		2523 => to_signed(7849, LUT_AMPL_WIDTH),
		2524 => to_signed(7852, LUT_AMPL_WIDTH),
		2525 => to_signed(7855, LUT_AMPL_WIDTH),
		2526 => to_signed(7858, LUT_AMPL_WIDTH),
		2527 => to_signed(7861, LUT_AMPL_WIDTH),
		2528 => to_signed(7864, LUT_AMPL_WIDTH),
		2529 => to_signed(7867, LUT_AMPL_WIDTH),
		2530 => to_signed(7870, LUT_AMPL_WIDTH),
		2531 => to_signed(7873, LUT_AMPL_WIDTH),
		2532 => to_signed(7876, LUT_AMPL_WIDTH),
		2533 => to_signed(7879, LUT_AMPL_WIDTH),
		2534 => to_signed(7882, LUT_AMPL_WIDTH),
		2535 => to_signed(7886, LUT_AMPL_WIDTH),
		2536 => to_signed(7889, LUT_AMPL_WIDTH),
		2537 => to_signed(7892, LUT_AMPL_WIDTH),
		2538 => to_signed(7895, LUT_AMPL_WIDTH),
		2539 => to_signed(7898, LUT_AMPL_WIDTH),
		2540 => to_signed(7901, LUT_AMPL_WIDTH),
		2541 => to_signed(7904, LUT_AMPL_WIDTH),
		2542 => to_signed(7907, LUT_AMPL_WIDTH),
		2543 => to_signed(7910, LUT_AMPL_WIDTH),
		2544 => to_signed(7913, LUT_AMPL_WIDTH),
		2545 => to_signed(7916, LUT_AMPL_WIDTH),
		2546 => to_signed(7919, LUT_AMPL_WIDTH),
		2547 => to_signed(7922, LUT_AMPL_WIDTH),
		2548 => to_signed(7925, LUT_AMPL_WIDTH),
		2549 => to_signed(7928, LUT_AMPL_WIDTH),
		2550 => to_signed(7931, LUT_AMPL_WIDTH),
		2551 => to_signed(7934, LUT_AMPL_WIDTH),
		2552 => to_signed(7937, LUT_AMPL_WIDTH),
		2553 => to_signed(7940, LUT_AMPL_WIDTH),
		2554 => to_signed(7943, LUT_AMPL_WIDTH),
		2555 => to_signed(7946, LUT_AMPL_WIDTH),
		2556 => to_signed(7950, LUT_AMPL_WIDTH),
		2557 => to_signed(7953, LUT_AMPL_WIDTH),
		2558 => to_signed(7956, LUT_AMPL_WIDTH),
		2559 => to_signed(7959, LUT_AMPL_WIDTH),
		2560 => to_signed(7962, LUT_AMPL_WIDTH),
		2561 => to_signed(7965, LUT_AMPL_WIDTH),
		2562 => to_signed(7968, LUT_AMPL_WIDTH),
		2563 => to_signed(7971, LUT_AMPL_WIDTH),
		2564 => to_signed(7974, LUT_AMPL_WIDTH),
		2565 => to_signed(7977, LUT_AMPL_WIDTH),
		2566 => to_signed(7980, LUT_AMPL_WIDTH),
		2567 => to_signed(7983, LUT_AMPL_WIDTH),
		2568 => to_signed(7986, LUT_AMPL_WIDTH),
		2569 => to_signed(7989, LUT_AMPL_WIDTH),
		2570 => to_signed(7992, LUT_AMPL_WIDTH),
		2571 => to_signed(7995, LUT_AMPL_WIDTH),
		2572 => to_signed(7998, LUT_AMPL_WIDTH),
		2573 => to_signed(8001, LUT_AMPL_WIDTH),
		2574 => to_signed(8004, LUT_AMPL_WIDTH),
		2575 => to_signed(8007, LUT_AMPL_WIDTH),
		2576 => to_signed(8010, LUT_AMPL_WIDTH),
		2577 => to_signed(8014, LUT_AMPL_WIDTH),
		2578 => to_signed(8017, LUT_AMPL_WIDTH),
		2579 => to_signed(8020, LUT_AMPL_WIDTH),
		2580 => to_signed(8023, LUT_AMPL_WIDTH),
		2581 => to_signed(8026, LUT_AMPL_WIDTH),
		2582 => to_signed(8029, LUT_AMPL_WIDTH),
		2583 => to_signed(8032, LUT_AMPL_WIDTH),
		2584 => to_signed(8035, LUT_AMPL_WIDTH),
		2585 => to_signed(8038, LUT_AMPL_WIDTH),
		2586 => to_signed(8041, LUT_AMPL_WIDTH),
		2587 => to_signed(8044, LUT_AMPL_WIDTH),
		2588 => to_signed(8047, LUT_AMPL_WIDTH),
		2589 => to_signed(8050, LUT_AMPL_WIDTH),
		2590 => to_signed(8053, LUT_AMPL_WIDTH),
		2591 => to_signed(8056, LUT_AMPL_WIDTH),
		2592 => to_signed(8059, LUT_AMPL_WIDTH),
		2593 => to_signed(8062, LUT_AMPL_WIDTH),
		2594 => to_signed(8065, LUT_AMPL_WIDTH),
		2595 => to_signed(8068, LUT_AMPL_WIDTH),
		2596 => to_signed(8071, LUT_AMPL_WIDTH),
		2597 => to_signed(8074, LUT_AMPL_WIDTH),
		2598 => to_signed(8077, LUT_AMPL_WIDTH),
		2599 => to_signed(8081, LUT_AMPL_WIDTH),
		2600 => to_signed(8084, LUT_AMPL_WIDTH),
		2601 => to_signed(8087, LUT_AMPL_WIDTH),
		2602 => to_signed(8090, LUT_AMPL_WIDTH),
		2603 => to_signed(8093, LUT_AMPL_WIDTH),
		2604 => to_signed(8096, LUT_AMPL_WIDTH),
		2605 => to_signed(8099, LUT_AMPL_WIDTH),
		2606 => to_signed(8102, LUT_AMPL_WIDTH),
		2607 => to_signed(8105, LUT_AMPL_WIDTH),
		2608 => to_signed(8108, LUT_AMPL_WIDTH),
		2609 => to_signed(8111, LUT_AMPL_WIDTH),
		2610 => to_signed(8114, LUT_AMPL_WIDTH),
		2611 => to_signed(8117, LUT_AMPL_WIDTH),
		2612 => to_signed(8120, LUT_AMPL_WIDTH),
		2613 => to_signed(8123, LUT_AMPL_WIDTH),
		2614 => to_signed(8126, LUT_AMPL_WIDTH),
		2615 => to_signed(8129, LUT_AMPL_WIDTH),
		2616 => to_signed(8132, LUT_AMPL_WIDTH),
		2617 => to_signed(8135, LUT_AMPL_WIDTH),
		2618 => to_signed(8138, LUT_AMPL_WIDTH),
		2619 => to_signed(8141, LUT_AMPL_WIDTH),
		2620 => to_signed(8144, LUT_AMPL_WIDTH),
		2621 => to_signed(8147, LUT_AMPL_WIDTH),
		2622 => to_signed(8151, LUT_AMPL_WIDTH),
		2623 => to_signed(8154, LUT_AMPL_WIDTH),
		2624 => to_signed(8157, LUT_AMPL_WIDTH),
		2625 => to_signed(8160, LUT_AMPL_WIDTH),
		2626 => to_signed(8163, LUT_AMPL_WIDTH),
		2627 => to_signed(8166, LUT_AMPL_WIDTH),
		2628 => to_signed(8169, LUT_AMPL_WIDTH),
		2629 => to_signed(8172, LUT_AMPL_WIDTH),
		2630 => to_signed(8175, LUT_AMPL_WIDTH),
		2631 => to_signed(8178, LUT_AMPL_WIDTH),
		2632 => to_signed(8181, LUT_AMPL_WIDTH),
		2633 => to_signed(8184, LUT_AMPL_WIDTH),
		2634 => to_signed(8187, LUT_AMPL_WIDTH),
		2635 => to_signed(8190, LUT_AMPL_WIDTH),
		2636 => to_signed(8193, LUT_AMPL_WIDTH),
		2637 => to_signed(8196, LUT_AMPL_WIDTH),
		2638 => to_signed(8199, LUT_AMPL_WIDTH),
		2639 => to_signed(8202, LUT_AMPL_WIDTH),
		2640 => to_signed(8205, LUT_AMPL_WIDTH),
		2641 => to_signed(8208, LUT_AMPL_WIDTH),
		2642 => to_signed(8211, LUT_AMPL_WIDTH),
		2643 => to_signed(8214, LUT_AMPL_WIDTH),
		2644 => to_signed(8217, LUT_AMPL_WIDTH),
		2645 => to_signed(8220, LUT_AMPL_WIDTH),
		2646 => to_signed(8224, LUT_AMPL_WIDTH),
		2647 => to_signed(8227, LUT_AMPL_WIDTH),
		2648 => to_signed(8230, LUT_AMPL_WIDTH),
		2649 => to_signed(8233, LUT_AMPL_WIDTH),
		2650 => to_signed(8236, LUT_AMPL_WIDTH),
		2651 => to_signed(8239, LUT_AMPL_WIDTH),
		2652 => to_signed(8242, LUT_AMPL_WIDTH),
		2653 => to_signed(8245, LUT_AMPL_WIDTH),
		2654 => to_signed(8248, LUT_AMPL_WIDTH),
		2655 => to_signed(8251, LUT_AMPL_WIDTH),
		2656 => to_signed(8254, LUT_AMPL_WIDTH),
		2657 => to_signed(8257, LUT_AMPL_WIDTH),
		2658 => to_signed(8260, LUT_AMPL_WIDTH),
		2659 => to_signed(8263, LUT_AMPL_WIDTH),
		2660 => to_signed(8266, LUT_AMPL_WIDTH),
		2661 => to_signed(8269, LUT_AMPL_WIDTH),
		2662 => to_signed(8272, LUT_AMPL_WIDTH),
		2663 => to_signed(8275, LUT_AMPL_WIDTH),
		2664 => to_signed(8278, LUT_AMPL_WIDTH),
		2665 => to_signed(8281, LUT_AMPL_WIDTH),
		2666 => to_signed(8284, LUT_AMPL_WIDTH),
		2667 => to_signed(8287, LUT_AMPL_WIDTH),
		2668 => to_signed(8290, LUT_AMPL_WIDTH),
		2669 => to_signed(8293, LUT_AMPL_WIDTH),
		2670 => to_signed(8296, LUT_AMPL_WIDTH),
		2671 => to_signed(8300, LUT_AMPL_WIDTH),
		2672 => to_signed(8303, LUT_AMPL_WIDTH),
		2673 => to_signed(8306, LUT_AMPL_WIDTH),
		2674 => to_signed(8309, LUT_AMPL_WIDTH),
		2675 => to_signed(8312, LUT_AMPL_WIDTH),
		2676 => to_signed(8315, LUT_AMPL_WIDTH),
		2677 => to_signed(8318, LUT_AMPL_WIDTH),
		2678 => to_signed(8321, LUT_AMPL_WIDTH),
		2679 => to_signed(8324, LUT_AMPL_WIDTH),
		2680 => to_signed(8327, LUT_AMPL_WIDTH),
		2681 => to_signed(8330, LUT_AMPL_WIDTH),
		2682 => to_signed(8333, LUT_AMPL_WIDTH),
		2683 => to_signed(8336, LUT_AMPL_WIDTH),
		2684 => to_signed(8339, LUT_AMPL_WIDTH),
		2685 => to_signed(8342, LUT_AMPL_WIDTH),
		2686 => to_signed(8345, LUT_AMPL_WIDTH),
		2687 => to_signed(8348, LUT_AMPL_WIDTH),
		2688 => to_signed(8351, LUT_AMPL_WIDTH),
		2689 => to_signed(8354, LUT_AMPL_WIDTH),
		2690 => to_signed(8357, LUT_AMPL_WIDTH),
		2691 => to_signed(8360, LUT_AMPL_WIDTH),
		2692 => to_signed(8363, LUT_AMPL_WIDTH),
		2693 => to_signed(8366, LUT_AMPL_WIDTH),
		2694 => to_signed(8369, LUT_AMPL_WIDTH),
		2695 => to_signed(8372, LUT_AMPL_WIDTH),
		2696 => to_signed(8375, LUT_AMPL_WIDTH),
		2697 => to_signed(8379, LUT_AMPL_WIDTH),
		2698 => to_signed(8382, LUT_AMPL_WIDTH),
		2699 => to_signed(8385, LUT_AMPL_WIDTH),
		2700 => to_signed(8388, LUT_AMPL_WIDTH),
		2701 => to_signed(8391, LUT_AMPL_WIDTH),
		2702 => to_signed(8394, LUT_AMPL_WIDTH),
		2703 => to_signed(8397, LUT_AMPL_WIDTH),
		2704 => to_signed(8400, LUT_AMPL_WIDTH),
		2705 => to_signed(8403, LUT_AMPL_WIDTH),
		2706 => to_signed(8406, LUT_AMPL_WIDTH),
		2707 => to_signed(8409, LUT_AMPL_WIDTH),
		2708 => to_signed(8412, LUT_AMPL_WIDTH),
		2709 => to_signed(8415, LUT_AMPL_WIDTH),
		2710 => to_signed(8418, LUT_AMPL_WIDTH),
		2711 => to_signed(8421, LUT_AMPL_WIDTH),
		2712 => to_signed(8424, LUT_AMPL_WIDTH),
		2713 => to_signed(8427, LUT_AMPL_WIDTH),
		2714 => to_signed(8430, LUT_AMPL_WIDTH),
		2715 => to_signed(8433, LUT_AMPL_WIDTH),
		2716 => to_signed(8436, LUT_AMPL_WIDTH),
		2717 => to_signed(8439, LUT_AMPL_WIDTH),
		2718 => to_signed(8442, LUT_AMPL_WIDTH),
		2719 => to_signed(8445, LUT_AMPL_WIDTH),
		2720 => to_signed(8448, LUT_AMPL_WIDTH),
		2721 => to_signed(8451, LUT_AMPL_WIDTH),
		2722 => to_signed(8454, LUT_AMPL_WIDTH),
		2723 => to_signed(8457, LUT_AMPL_WIDTH),
		2724 => to_signed(8460, LUT_AMPL_WIDTH),
		2725 => to_signed(8464, LUT_AMPL_WIDTH),
		2726 => to_signed(8467, LUT_AMPL_WIDTH),
		2727 => to_signed(8470, LUT_AMPL_WIDTH),
		2728 => to_signed(8473, LUT_AMPL_WIDTH),
		2729 => to_signed(8476, LUT_AMPL_WIDTH),
		2730 => to_signed(8479, LUT_AMPL_WIDTH),
		2731 => to_signed(8482, LUT_AMPL_WIDTH),
		2732 => to_signed(8485, LUT_AMPL_WIDTH),
		2733 => to_signed(8488, LUT_AMPL_WIDTH),
		2734 => to_signed(8491, LUT_AMPL_WIDTH),
		2735 => to_signed(8494, LUT_AMPL_WIDTH),
		2736 => to_signed(8497, LUT_AMPL_WIDTH),
		2737 => to_signed(8500, LUT_AMPL_WIDTH),
		2738 => to_signed(8503, LUT_AMPL_WIDTH),
		2739 => to_signed(8506, LUT_AMPL_WIDTH),
		2740 => to_signed(8509, LUT_AMPL_WIDTH),
		2741 => to_signed(8512, LUT_AMPL_WIDTH),
		2742 => to_signed(8515, LUT_AMPL_WIDTH),
		2743 => to_signed(8518, LUT_AMPL_WIDTH),
		2744 => to_signed(8521, LUT_AMPL_WIDTH),
		2745 => to_signed(8524, LUT_AMPL_WIDTH),
		2746 => to_signed(8527, LUT_AMPL_WIDTH),
		2747 => to_signed(8530, LUT_AMPL_WIDTH),
		2748 => to_signed(8533, LUT_AMPL_WIDTH),
		2749 => to_signed(8536, LUT_AMPL_WIDTH),
		2750 => to_signed(8539, LUT_AMPL_WIDTH),
		2751 => to_signed(8542, LUT_AMPL_WIDTH),
		2752 => to_signed(8545, LUT_AMPL_WIDTH),
		2753 => to_signed(8548, LUT_AMPL_WIDTH),
		2754 => to_signed(8552, LUT_AMPL_WIDTH),
		2755 => to_signed(8555, LUT_AMPL_WIDTH),
		2756 => to_signed(8558, LUT_AMPL_WIDTH),
		2757 => to_signed(8561, LUT_AMPL_WIDTH),
		2758 => to_signed(8564, LUT_AMPL_WIDTH),
		2759 => to_signed(8567, LUT_AMPL_WIDTH),
		2760 => to_signed(8570, LUT_AMPL_WIDTH),
		2761 => to_signed(8573, LUT_AMPL_WIDTH),
		2762 => to_signed(8576, LUT_AMPL_WIDTH),
		2763 => to_signed(8579, LUT_AMPL_WIDTH),
		2764 => to_signed(8582, LUT_AMPL_WIDTH),
		2765 => to_signed(8585, LUT_AMPL_WIDTH),
		2766 => to_signed(8588, LUT_AMPL_WIDTH),
		2767 => to_signed(8591, LUT_AMPL_WIDTH),
		2768 => to_signed(8594, LUT_AMPL_WIDTH),
		2769 => to_signed(8597, LUT_AMPL_WIDTH),
		2770 => to_signed(8600, LUT_AMPL_WIDTH),
		2771 => to_signed(8603, LUT_AMPL_WIDTH),
		2772 => to_signed(8606, LUT_AMPL_WIDTH),
		2773 => to_signed(8609, LUT_AMPL_WIDTH),
		2774 => to_signed(8612, LUT_AMPL_WIDTH),
		2775 => to_signed(8615, LUT_AMPL_WIDTH),
		2776 => to_signed(8618, LUT_AMPL_WIDTH),
		2777 => to_signed(8621, LUT_AMPL_WIDTH),
		2778 => to_signed(8624, LUT_AMPL_WIDTH),
		2779 => to_signed(8627, LUT_AMPL_WIDTH),
		2780 => to_signed(8630, LUT_AMPL_WIDTH),
		2781 => to_signed(8633, LUT_AMPL_WIDTH),
		2782 => to_signed(8636, LUT_AMPL_WIDTH),
		2783 => to_signed(8639, LUT_AMPL_WIDTH),
		2784 => to_signed(8642, LUT_AMPL_WIDTH),
		2785 => to_signed(8645, LUT_AMPL_WIDTH),
		2786 => to_signed(8649, LUT_AMPL_WIDTH),
		2787 => to_signed(8652, LUT_AMPL_WIDTH),
		2788 => to_signed(8655, LUT_AMPL_WIDTH),
		2789 => to_signed(8658, LUT_AMPL_WIDTH),
		2790 => to_signed(8661, LUT_AMPL_WIDTH),
		2791 => to_signed(8664, LUT_AMPL_WIDTH),
		2792 => to_signed(8667, LUT_AMPL_WIDTH),
		2793 => to_signed(8670, LUT_AMPL_WIDTH),
		2794 => to_signed(8673, LUT_AMPL_WIDTH),
		2795 => to_signed(8676, LUT_AMPL_WIDTH),
		2796 => to_signed(8679, LUT_AMPL_WIDTH),
		2797 => to_signed(8682, LUT_AMPL_WIDTH),
		2798 => to_signed(8685, LUT_AMPL_WIDTH),
		2799 => to_signed(8688, LUT_AMPL_WIDTH),
		2800 => to_signed(8691, LUT_AMPL_WIDTH),
		2801 => to_signed(8694, LUT_AMPL_WIDTH),
		2802 => to_signed(8697, LUT_AMPL_WIDTH),
		2803 => to_signed(8700, LUT_AMPL_WIDTH),
		2804 => to_signed(8703, LUT_AMPL_WIDTH),
		2805 => to_signed(8706, LUT_AMPL_WIDTH),
		2806 => to_signed(8709, LUT_AMPL_WIDTH),
		2807 => to_signed(8712, LUT_AMPL_WIDTH),
		2808 => to_signed(8715, LUT_AMPL_WIDTH),
		2809 => to_signed(8718, LUT_AMPL_WIDTH),
		2810 => to_signed(8721, LUT_AMPL_WIDTH),
		2811 => to_signed(8724, LUT_AMPL_WIDTH),
		2812 => to_signed(8727, LUT_AMPL_WIDTH),
		2813 => to_signed(8730, LUT_AMPL_WIDTH),
		2814 => to_signed(8733, LUT_AMPL_WIDTH),
		2815 => to_signed(8736, LUT_AMPL_WIDTH),
		2816 => to_signed(8739, LUT_AMPL_WIDTH),
		2817 => to_signed(8742, LUT_AMPL_WIDTH),
		2818 => to_signed(8745, LUT_AMPL_WIDTH),
		2819 => to_signed(8748, LUT_AMPL_WIDTH),
		2820 => to_signed(8751, LUT_AMPL_WIDTH),
		2821 => to_signed(8755, LUT_AMPL_WIDTH),
		2822 => to_signed(8758, LUT_AMPL_WIDTH),
		2823 => to_signed(8761, LUT_AMPL_WIDTH),
		2824 => to_signed(8764, LUT_AMPL_WIDTH),
		2825 => to_signed(8767, LUT_AMPL_WIDTH),
		2826 => to_signed(8770, LUT_AMPL_WIDTH),
		2827 => to_signed(8773, LUT_AMPL_WIDTH),
		2828 => to_signed(8776, LUT_AMPL_WIDTH),
		2829 => to_signed(8779, LUT_AMPL_WIDTH),
		2830 => to_signed(8782, LUT_AMPL_WIDTH),
		2831 => to_signed(8785, LUT_AMPL_WIDTH),
		2832 => to_signed(8788, LUT_AMPL_WIDTH),
		2833 => to_signed(8791, LUT_AMPL_WIDTH),
		2834 => to_signed(8794, LUT_AMPL_WIDTH),
		2835 => to_signed(8797, LUT_AMPL_WIDTH),
		2836 => to_signed(8800, LUT_AMPL_WIDTH),
		2837 => to_signed(8803, LUT_AMPL_WIDTH),
		2838 => to_signed(8806, LUT_AMPL_WIDTH),
		2839 => to_signed(8809, LUT_AMPL_WIDTH),
		2840 => to_signed(8812, LUT_AMPL_WIDTH),
		2841 => to_signed(8815, LUT_AMPL_WIDTH),
		2842 => to_signed(8818, LUT_AMPL_WIDTH),
		2843 => to_signed(8821, LUT_AMPL_WIDTH),
		2844 => to_signed(8824, LUT_AMPL_WIDTH),
		2845 => to_signed(8827, LUT_AMPL_WIDTH),
		2846 => to_signed(8830, LUT_AMPL_WIDTH),
		2847 => to_signed(8833, LUT_AMPL_WIDTH),
		2848 => to_signed(8836, LUT_AMPL_WIDTH),
		2849 => to_signed(8839, LUT_AMPL_WIDTH),
		2850 => to_signed(8842, LUT_AMPL_WIDTH),
		2851 => to_signed(8845, LUT_AMPL_WIDTH),
		2852 => to_signed(8848, LUT_AMPL_WIDTH),
		2853 => to_signed(8851, LUT_AMPL_WIDTH),
		2854 => to_signed(8854, LUT_AMPL_WIDTH),
		2855 => to_signed(8857, LUT_AMPL_WIDTH),
		2856 => to_signed(8860, LUT_AMPL_WIDTH),
		2857 => to_signed(8863, LUT_AMPL_WIDTH),
		2858 => to_signed(8866, LUT_AMPL_WIDTH),
		2859 => to_signed(8869, LUT_AMPL_WIDTH),
		2860 => to_signed(8873, LUT_AMPL_WIDTH),
		2861 => to_signed(8876, LUT_AMPL_WIDTH),
		2862 => to_signed(8879, LUT_AMPL_WIDTH),
		2863 => to_signed(8882, LUT_AMPL_WIDTH),
		2864 => to_signed(8885, LUT_AMPL_WIDTH),
		2865 => to_signed(8888, LUT_AMPL_WIDTH),
		2866 => to_signed(8891, LUT_AMPL_WIDTH),
		2867 => to_signed(8894, LUT_AMPL_WIDTH),
		2868 => to_signed(8897, LUT_AMPL_WIDTH),
		2869 => to_signed(8900, LUT_AMPL_WIDTH),
		2870 => to_signed(8903, LUT_AMPL_WIDTH),
		2871 => to_signed(8906, LUT_AMPL_WIDTH),
		2872 => to_signed(8909, LUT_AMPL_WIDTH),
		2873 => to_signed(8912, LUT_AMPL_WIDTH),
		2874 => to_signed(8915, LUT_AMPL_WIDTH),
		2875 => to_signed(8918, LUT_AMPL_WIDTH),
		2876 => to_signed(8921, LUT_AMPL_WIDTH),
		2877 => to_signed(8924, LUT_AMPL_WIDTH),
		2878 => to_signed(8927, LUT_AMPL_WIDTH),
		2879 => to_signed(8930, LUT_AMPL_WIDTH),
		2880 => to_signed(8933, LUT_AMPL_WIDTH),
		2881 => to_signed(8936, LUT_AMPL_WIDTH),
		2882 => to_signed(8939, LUT_AMPL_WIDTH),
		2883 => to_signed(8942, LUT_AMPL_WIDTH),
		2884 => to_signed(8945, LUT_AMPL_WIDTH),
		2885 => to_signed(8948, LUT_AMPL_WIDTH),
		2886 => to_signed(8951, LUT_AMPL_WIDTH),
		2887 => to_signed(8954, LUT_AMPL_WIDTH),
		2888 => to_signed(8957, LUT_AMPL_WIDTH),
		2889 => to_signed(8960, LUT_AMPL_WIDTH),
		2890 => to_signed(8963, LUT_AMPL_WIDTH),
		2891 => to_signed(8966, LUT_AMPL_WIDTH),
		2892 => to_signed(8969, LUT_AMPL_WIDTH),
		2893 => to_signed(8972, LUT_AMPL_WIDTH),
		2894 => to_signed(8975, LUT_AMPL_WIDTH),
		2895 => to_signed(8978, LUT_AMPL_WIDTH),
		2896 => to_signed(8981, LUT_AMPL_WIDTH),
		2897 => to_signed(8984, LUT_AMPL_WIDTH),
		2898 => to_signed(8987, LUT_AMPL_WIDTH),
		2899 => to_signed(8990, LUT_AMPL_WIDTH),
		2900 => to_signed(8993, LUT_AMPL_WIDTH),
		2901 => to_signed(8996, LUT_AMPL_WIDTH),
		2902 => to_signed(8999, LUT_AMPL_WIDTH),
		2903 => to_signed(9002, LUT_AMPL_WIDTH),
		2904 => to_signed(9006, LUT_AMPL_WIDTH),
		2905 => to_signed(9009, LUT_AMPL_WIDTH),
		2906 => to_signed(9012, LUT_AMPL_WIDTH),
		2907 => to_signed(9015, LUT_AMPL_WIDTH),
		2908 => to_signed(9018, LUT_AMPL_WIDTH),
		2909 => to_signed(9021, LUT_AMPL_WIDTH),
		2910 => to_signed(9024, LUT_AMPL_WIDTH),
		2911 => to_signed(9027, LUT_AMPL_WIDTH),
		2912 => to_signed(9030, LUT_AMPL_WIDTH),
		2913 => to_signed(9033, LUT_AMPL_WIDTH),
		2914 => to_signed(9036, LUT_AMPL_WIDTH),
		2915 => to_signed(9039, LUT_AMPL_WIDTH),
		2916 => to_signed(9042, LUT_AMPL_WIDTH),
		2917 => to_signed(9045, LUT_AMPL_WIDTH),
		2918 => to_signed(9048, LUT_AMPL_WIDTH),
		2919 => to_signed(9051, LUT_AMPL_WIDTH),
		2920 => to_signed(9054, LUT_AMPL_WIDTH),
		2921 => to_signed(9057, LUT_AMPL_WIDTH),
		2922 => to_signed(9060, LUT_AMPL_WIDTH),
		2923 => to_signed(9063, LUT_AMPL_WIDTH),
		2924 => to_signed(9066, LUT_AMPL_WIDTH),
		2925 => to_signed(9069, LUT_AMPL_WIDTH),
		2926 => to_signed(9072, LUT_AMPL_WIDTH),
		2927 => to_signed(9075, LUT_AMPL_WIDTH),
		2928 => to_signed(9078, LUT_AMPL_WIDTH),
		2929 => to_signed(9081, LUT_AMPL_WIDTH),
		2930 => to_signed(9084, LUT_AMPL_WIDTH),
		2931 => to_signed(9087, LUT_AMPL_WIDTH),
		2932 => to_signed(9090, LUT_AMPL_WIDTH),
		2933 => to_signed(9093, LUT_AMPL_WIDTH),
		2934 => to_signed(9096, LUT_AMPL_WIDTH),
		2935 => to_signed(9099, LUT_AMPL_WIDTH),
		2936 => to_signed(9102, LUT_AMPL_WIDTH),
		2937 => to_signed(9105, LUT_AMPL_WIDTH),
		2938 => to_signed(9108, LUT_AMPL_WIDTH),
		2939 => to_signed(9111, LUT_AMPL_WIDTH),
		2940 => to_signed(9114, LUT_AMPL_WIDTH),
		2941 => to_signed(9117, LUT_AMPL_WIDTH),
		2942 => to_signed(9120, LUT_AMPL_WIDTH),
		2943 => to_signed(9123, LUT_AMPL_WIDTH),
		2944 => to_signed(9126, LUT_AMPL_WIDTH),
		2945 => to_signed(9129, LUT_AMPL_WIDTH),
		2946 => to_signed(9132, LUT_AMPL_WIDTH),
		2947 => to_signed(9135, LUT_AMPL_WIDTH),
		2948 => to_signed(9138, LUT_AMPL_WIDTH),
		2949 => to_signed(9141, LUT_AMPL_WIDTH),
		2950 => to_signed(9144, LUT_AMPL_WIDTH),
		2951 => to_signed(9147, LUT_AMPL_WIDTH),
		2952 => to_signed(9150, LUT_AMPL_WIDTH),
		2953 => to_signed(9153, LUT_AMPL_WIDTH),
		2954 => to_signed(9156, LUT_AMPL_WIDTH),
		2955 => to_signed(9159, LUT_AMPL_WIDTH),
		2956 => to_signed(9162, LUT_AMPL_WIDTH),
		2957 => to_signed(9165, LUT_AMPL_WIDTH),
		2958 => to_signed(9168, LUT_AMPL_WIDTH),
		2959 => to_signed(9172, LUT_AMPL_WIDTH),
		2960 => to_signed(9175, LUT_AMPL_WIDTH),
		2961 => to_signed(9178, LUT_AMPL_WIDTH),
		2962 => to_signed(9181, LUT_AMPL_WIDTH),
		2963 => to_signed(9184, LUT_AMPL_WIDTH),
		2964 => to_signed(9187, LUT_AMPL_WIDTH),
		2965 => to_signed(9190, LUT_AMPL_WIDTH),
		2966 => to_signed(9193, LUT_AMPL_WIDTH),
		2967 => to_signed(9196, LUT_AMPL_WIDTH),
		2968 => to_signed(9199, LUT_AMPL_WIDTH),
		2969 => to_signed(9202, LUT_AMPL_WIDTH),
		2970 => to_signed(9205, LUT_AMPL_WIDTH),
		2971 => to_signed(9208, LUT_AMPL_WIDTH),
		2972 => to_signed(9211, LUT_AMPL_WIDTH),
		2973 => to_signed(9214, LUT_AMPL_WIDTH),
		2974 => to_signed(9217, LUT_AMPL_WIDTH),
		2975 => to_signed(9220, LUT_AMPL_WIDTH),
		2976 => to_signed(9223, LUT_AMPL_WIDTH),
		2977 => to_signed(9226, LUT_AMPL_WIDTH),
		2978 => to_signed(9229, LUT_AMPL_WIDTH),
		2979 => to_signed(9232, LUT_AMPL_WIDTH),
		2980 => to_signed(9235, LUT_AMPL_WIDTH),
		2981 => to_signed(9238, LUT_AMPL_WIDTH),
		2982 => to_signed(9241, LUT_AMPL_WIDTH),
		2983 => to_signed(9244, LUT_AMPL_WIDTH),
		2984 => to_signed(9247, LUT_AMPL_WIDTH),
		2985 => to_signed(9250, LUT_AMPL_WIDTH),
		2986 => to_signed(9253, LUT_AMPL_WIDTH),
		2987 => to_signed(9256, LUT_AMPL_WIDTH),
		2988 => to_signed(9259, LUT_AMPL_WIDTH),
		2989 => to_signed(9262, LUT_AMPL_WIDTH),
		2990 => to_signed(9265, LUT_AMPL_WIDTH),
		2991 => to_signed(9268, LUT_AMPL_WIDTH),
		2992 => to_signed(9271, LUT_AMPL_WIDTH),
		2993 => to_signed(9274, LUT_AMPL_WIDTH),
		2994 => to_signed(9277, LUT_AMPL_WIDTH),
		2995 => to_signed(9280, LUT_AMPL_WIDTH),
		2996 => to_signed(9283, LUT_AMPL_WIDTH),
		2997 => to_signed(9286, LUT_AMPL_WIDTH),
		2998 => to_signed(9289, LUT_AMPL_WIDTH),
		2999 => to_signed(9292, LUT_AMPL_WIDTH),
		3000 => to_signed(9295, LUT_AMPL_WIDTH),
		3001 => to_signed(9298, LUT_AMPL_WIDTH),
		3002 => to_signed(9301, LUT_AMPL_WIDTH),
		3003 => to_signed(9304, LUT_AMPL_WIDTH),
		3004 => to_signed(9307, LUT_AMPL_WIDTH),
		3005 => to_signed(9310, LUT_AMPL_WIDTH),
		3006 => to_signed(9313, LUT_AMPL_WIDTH),
		3007 => to_signed(9316, LUT_AMPL_WIDTH),
		3008 => to_signed(9319, LUT_AMPL_WIDTH),
		3009 => to_signed(9322, LUT_AMPL_WIDTH),
		3010 => to_signed(9325, LUT_AMPL_WIDTH),
		3011 => to_signed(9328, LUT_AMPL_WIDTH),
		3012 => to_signed(9331, LUT_AMPL_WIDTH),
		3013 => to_signed(9334, LUT_AMPL_WIDTH),
		3014 => to_signed(9337, LUT_AMPL_WIDTH),
		3015 => to_signed(9340, LUT_AMPL_WIDTH),
		3016 => to_signed(9343, LUT_AMPL_WIDTH),
		3017 => to_signed(9346, LUT_AMPL_WIDTH),
		3018 => to_signed(9349, LUT_AMPL_WIDTH),
		3019 => to_signed(9352, LUT_AMPL_WIDTH),
		3020 => to_signed(9355, LUT_AMPL_WIDTH),
		3021 => to_signed(9358, LUT_AMPL_WIDTH),
		3022 => to_signed(9361, LUT_AMPL_WIDTH),
		3023 => to_signed(9364, LUT_AMPL_WIDTH),
		3024 => to_signed(9367, LUT_AMPL_WIDTH),
		3025 => to_signed(9370, LUT_AMPL_WIDTH),
		3026 => to_signed(9373, LUT_AMPL_WIDTH),
		3027 => to_signed(9376, LUT_AMPL_WIDTH),
		3028 => to_signed(9379, LUT_AMPL_WIDTH),
		3029 => to_signed(9382, LUT_AMPL_WIDTH),
		3030 => to_signed(9385, LUT_AMPL_WIDTH),
		3031 => to_signed(9388, LUT_AMPL_WIDTH),
		3032 => to_signed(9391, LUT_AMPL_WIDTH),
		3033 => to_signed(9394, LUT_AMPL_WIDTH),
		3034 => to_signed(9397, LUT_AMPL_WIDTH),
		3035 => to_signed(9400, LUT_AMPL_WIDTH),
		3036 => to_signed(9403, LUT_AMPL_WIDTH),
		3037 => to_signed(9406, LUT_AMPL_WIDTH),
		3038 => to_signed(9409, LUT_AMPL_WIDTH),
		3039 => to_signed(9413, LUT_AMPL_WIDTH),
		3040 => to_signed(9416, LUT_AMPL_WIDTH),
		3041 => to_signed(9419, LUT_AMPL_WIDTH),
		3042 => to_signed(9422, LUT_AMPL_WIDTH),
		3043 => to_signed(9425, LUT_AMPL_WIDTH),
		3044 => to_signed(9428, LUT_AMPL_WIDTH),
		3045 => to_signed(9431, LUT_AMPL_WIDTH),
		3046 => to_signed(9434, LUT_AMPL_WIDTH),
		3047 => to_signed(9437, LUT_AMPL_WIDTH),
		3048 => to_signed(9440, LUT_AMPL_WIDTH),
		3049 => to_signed(9443, LUT_AMPL_WIDTH),
		3050 => to_signed(9446, LUT_AMPL_WIDTH),
		3051 => to_signed(9449, LUT_AMPL_WIDTH),
		3052 => to_signed(9452, LUT_AMPL_WIDTH),
		3053 => to_signed(9455, LUT_AMPL_WIDTH),
		3054 => to_signed(9458, LUT_AMPL_WIDTH),
		3055 => to_signed(9461, LUT_AMPL_WIDTH),
		3056 => to_signed(9464, LUT_AMPL_WIDTH),
		3057 => to_signed(9467, LUT_AMPL_WIDTH),
		3058 => to_signed(9470, LUT_AMPL_WIDTH),
		3059 => to_signed(9473, LUT_AMPL_WIDTH),
		3060 => to_signed(9476, LUT_AMPL_WIDTH),
		3061 => to_signed(9479, LUT_AMPL_WIDTH),
		3062 => to_signed(9482, LUT_AMPL_WIDTH),
		3063 => to_signed(9485, LUT_AMPL_WIDTH),
		3064 => to_signed(9488, LUT_AMPL_WIDTH),
		3065 => to_signed(9491, LUT_AMPL_WIDTH),
		3066 => to_signed(9494, LUT_AMPL_WIDTH),
		3067 => to_signed(9497, LUT_AMPL_WIDTH),
		3068 => to_signed(9500, LUT_AMPL_WIDTH),
		3069 => to_signed(9503, LUT_AMPL_WIDTH),
		3070 => to_signed(9506, LUT_AMPL_WIDTH),
		3071 => to_signed(9509, LUT_AMPL_WIDTH),
		3072 => to_signed(9512, LUT_AMPL_WIDTH),
		3073 => to_signed(9515, LUT_AMPL_WIDTH),
		3074 => to_signed(9518, LUT_AMPL_WIDTH),
		3075 => to_signed(9521, LUT_AMPL_WIDTH),
		3076 => to_signed(9524, LUT_AMPL_WIDTH),
		3077 => to_signed(9527, LUT_AMPL_WIDTH),
		3078 => to_signed(9530, LUT_AMPL_WIDTH),
		3079 => to_signed(9533, LUT_AMPL_WIDTH),
		3080 => to_signed(9536, LUT_AMPL_WIDTH),
		3081 => to_signed(9539, LUT_AMPL_WIDTH),
		3082 => to_signed(9542, LUT_AMPL_WIDTH),
		3083 => to_signed(9545, LUT_AMPL_WIDTH),
		3084 => to_signed(9548, LUT_AMPL_WIDTH),
		3085 => to_signed(9551, LUT_AMPL_WIDTH),
		3086 => to_signed(9554, LUT_AMPL_WIDTH),
		3087 => to_signed(9557, LUT_AMPL_WIDTH),
		3088 => to_signed(9560, LUT_AMPL_WIDTH),
		3089 => to_signed(9563, LUT_AMPL_WIDTH),
		3090 => to_signed(9566, LUT_AMPL_WIDTH),
		3091 => to_signed(9569, LUT_AMPL_WIDTH),
		3092 => to_signed(9572, LUT_AMPL_WIDTH),
		3093 => to_signed(9575, LUT_AMPL_WIDTH),
		3094 => to_signed(9578, LUT_AMPL_WIDTH),
		3095 => to_signed(9581, LUT_AMPL_WIDTH),
		3096 => to_signed(9584, LUT_AMPL_WIDTH),
		3097 => to_signed(9587, LUT_AMPL_WIDTH),
		3098 => to_signed(9590, LUT_AMPL_WIDTH),
		3099 => to_signed(9593, LUT_AMPL_WIDTH),
		3100 => to_signed(9596, LUT_AMPL_WIDTH),
		3101 => to_signed(9599, LUT_AMPL_WIDTH),
		3102 => to_signed(9602, LUT_AMPL_WIDTH),
		3103 => to_signed(9605, LUT_AMPL_WIDTH),
		3104 => to_signed(9608, LUT_AMPL_WIDTH),
		3105 => to_signed(9611, LUT_AMPL_WIDTH),
		3106 => to_signed(9614, LUT_AMPL_WIDTH),
		3107 => to_signed(9617, LUT_AMPL_WIDTH),
		3108 => to_signed(9620, LUT_AMPL_WIDTH),
		3109 => to_signed(9623, LUT_AMPL_WIDTH),
		3110 => to_signed(9626, LUT_AMPL_WIDTH),
		3111 => to_signed(9629, LUT_AMPL_WIDTH),
		3112 => to_signed(9632, LUT_AMPL_WIDTH),
		3113 => to_signed(9635, LUT_AMPL_WIDTH),
		3114 => to_signed(9638, LUT_AMPL_WIDTH),
		3115 => to_signed(9641, LUT_AMPL_WIDTH),
		3116 => to_signed(9644, LUT_AMPL_WIDTH),
		3117 => to_signed(9647, LUT_AMPL_WIDTH),
		3118 => to_signed(9650, LUT_AMPL_WIDTH),
		3119 => to_signed(9653, LUT_AMPL_WIDTH),
		3120 => to_signed(9656, LUT_AMPL_WIDTH),
		3121 => to_signed(9659, LUT_AMPL_WIDTH),
		3122 => to_signed(9662, LUT_AMPL_WIDTH),
		3123 => to_signed(9665, LUT_AMPL_WIDTH),
		3124 => to_signed(9668, LUT_AMPL_WIDTH),
		3125 => to_signed(9671, LUT_AMPL_WIDTH),
		3126 => to_signed(9674, LUT_AMPL_WIDTH),
		3127 => to_signed(9677, LUT_AMPL_WIDTH),
		3128 => to_signed(9680, LUT_AMPL_WIDTH),
		3129 => to_signed(9683, LUT_AMPL_WIDTH),
		3130 => to_signed(9686, LUT_AMPL_WIDTH),
		3131 => to_signed(9689, LUT_AMPL_WIDTH),
		3132 => to_signed(9692, LUT_AMPL_WIDTH),
		3133 => to_signed(9695, LUT_AMPL_WIDTH),
		3134 => to_signed(9698, LUT_AMPL_WIDTH),
		3135 => to_signed(9701, LUT_AMPL_WIDTH),
		3136 => to_signed(9704, LUT_AMPL_WIDTH),
		3137 => to_signed(9707, LUT_AMPL_WIDTH),
		3138 => to_signed(9710, LUT_AMPL_WIDTH),
		3139 => to_signed(9713, LUT_AMPL_WIDTH),
		3140 => to_signed(9716, LUT_AMPL_WIDTH),
		3141 => to_signed(9719, LUT_AMPL_WIDTH),
		3142 => to_signed(9722, LUT_AMPL_WIDTH),
		3143 => to_signed(9725, LUT_AMPL_WIDTH),
		3144 => to_signed(9728, LUT_AMPL_WIDTH),
		3145 => to_signed(9731, LUT_AMPL_WIDTH),
		3146 => to_signed(9734, LUT_AMPL_WIDTH),
		3147 => to_signed(9737, LUT_AMPL_WIDTH),
		3148 => to_signed(9740, LUT_AMPL_WIDTH),
		3149 => to_signed(9743, LUT_AMPL_WIDTH),
		3150 => to_signed(9746, LUT_AMPL_WIDTH),
		3151 => to_signed(9749, LUT_AMPL_WIDTH),
		3152 => to_signed(9752, LUT_AMPL_WIDTH),
		3153 => to_signed(9755, LUT_AMPL_WIDTH),
		3154 => to_signed(9758, LUT_AMPL_WIDTH),
		3155 => to_signed(9761, LUT_AMPL_WIDTH),
		3156 => to_signed(9764, LUT_AMPL_WIDTH),
		3157 => to_signed(9767, LUT_AMPL_WIDTH),
		3158 => to_signed(9770, LUT_AMPL_WIDTH),
		3159 => to_signed(9773, LUT_AMPL_WIDTH),
		3160 => to_signed(9776, LUT_AMPL_WIDTH),
		3161 => to_signed(9779, LUT_AMPL_WIDTH),
		3162 => to_signed(9782, LUT_AMPL_WIDTH),
		3163 => to_signed(9785, LUT_AMPL_WIDTH),
		3164 => to_signed(9788, LUT_AMPL_WIDTH),
		3165 => to_signed(9791, LUT_AMPL_WIDTH),
		3166 => to_signed(9794, LUT_AMPL_WIDTH),
		3167 => to_signed(9797, LUT_AMPL_WIDTH),
		3168 => to_signed(9800, LUT_AMPL_WIDTH),
		3169 => to_signed(9803, LUT_AMPL_WIDTH),
		3170 => to_signed(9806, LUT_AMPL_WIDTH),
		3171 => to_signed(9809, LUT_AMPL_WIDTH),
		3172 => to_signed(9812, LUT_AMPL_WIDTH),
		3173 => to_signed(9815, LUT_AMPL_WIDTH),
		3174 => to_signed(9818, LUT_AMPL_WIDTH),
		3175 => to_signed(9821, LUT_AMPL_WIDTH),
		3176 => to_signed(9824, LUT_AMPL_WIDTH),
		3177 => to_signed(9827, LUT_AMPL_WIDTH),
		3178 => to_signed(9830, LUT_AMPL_WIDTH),
		3179 => to_signed(9833, LUT_AMPL_WIDTH),
		3180 => to_signed(9836, LUT_AMPL_WIDTH),
		3181 => to_signed(9839, LUT_AMPL_WIDTH),
		3182 => to_signed(9842, LUT_AMPL_WIDTH),
		3183 => to_signed(9845, LUT_AMPL_WIDTH),
		3184 => to_signed(9848, LUT_AMPL_WIDTH),
		3185 => to_signed(9851, LUT_AMPL_WIDTH),
		3186 => to_signed(9854, LUT_AMPL_WIDTH),
		3187 => to_signed(9857, LUT_AMPL_WIDTH),
		3188 => to_signed(9860, LUT_AMPL_WIDTH),
		3189 => to_signed(9863, LUT_AMPL_WIDTH),
		3190 => to_signed(9866, LUT_AMPL_WIDTH),
		3191 => to_signed(9869, LUT_AMPL_WIDTH),
		3192 => to_signed(9872, LUT_AMPL_WIDTH),
		3193 => to_signed(9875, LUT_AMPL_WIDTH),
		3194 => to_signed(9878, LUT_AMPL_WIDTH),
		3195 => to_signed(9881, LUT_AMPL_WIDTH),
		3196 => to_signed(9884, LUT_AMPL_WIDTH),
		3197 => to_signed(9887, LUT_AMPL_WIDTH),
		3198 => to_signed(9890, LUT_AMPL_WIDTH),
		3199 => to_signed(9893, LUT_AMPL_WIDTH),
		3200 => to_signed(9896, LUT_AMPL_WIDTH),
		3201 => to_signed(9899, LUT_AMPL_WIDTH),
		3202 => to_signed(9902, LUT_AMPL_WIDTH),
		3203 => to_signed(9905, LUT_AMPL_WIDTH),
		3204 => to_signed(9908, LUT_AMPL_WIDTH),
		3205 => to_signed(9911, LUT_AMPL_WIDTH),
		3206 => to_signed(9914, LUT_AMPL_WIDTH),
		3207 => to_signed(9917, LUT_AMPL_WIDTH),
		3208 => to_signed(9920, LUT_AMPL_WIDTH),
		3209 => to_signed(9923, LUT_AMPL_WIDTH),
		3210 => to_signed(9926, LUT_AMPL_WIDTH),
		3211 => to_signed(9929, LUT_AMPL_WIDTH),
		3212 => to_signed(9932, LUT_AMPL_WIDTH),
		3213 => to_signed(9935, LUT_AMPL_WIDTH),
		3214 => to_signed(9938, LUT_AMPL_WIDTH),
		3215 => to_signed(9941, LUT_AMPL_WIDTH),
		3216 => to_signed(9944, LUT_AMPL_WIDTH),
		3217 => to_signed(9947, LUT_AMPL_WIDTH),
		3218 => to_signed(9950, LUT_AMPL_WIDTH),
		3219 => to_signed(9953, LUT_AMPL_WIDTH),
		3220 => to_signed(9956, LUT_AMPL_WIDTH),
		3221 => to_signed(9959, LUT_AMPL_WIDTH),
		3222 => to_signed(9962, LUT_AMPL_WIDTH),
		3223 => to_signed(9965, LUT_AMPL_WIDTH),
		3224 => to_signed(9968, LUT_AMPL_WIDTH),
		3225 => to_signed(9971, LUT_AMPL_WIDTH),
		3226 => to_signed(9974, LUT_AMPL_WIDTH),
		3227 => to_signed(9977, LUT_AMPL_WIDTH),
		3228 => to_signed(9980, LUT_AMPL_WIDTH),
		3229 => to_signed(9983, LUT_AMPL_WIDTH),
		3230 => to_signed(9986, LUT_AMPL_WIDTH),
		3231 => to_signed(9989, LUT_AMPL_WIDTH),
		3232 => to_signed(9992, LUT_AMPL_WIDTH),
		3233 => to_signed(9995, LUT_AMPL_WIDTH),
		3234 => to_signed(9998, LUT_AMPL_WIDTH),
		3235 => to_signed(10001, LUT_AMPL_WIDTH),
		3236 => to_signed(10004, LUT_AMPL_WIDTH),
		3237 => to_signed(10007, LUT_AMPL_WIDTH),
		3238 => to_signed(10010, LUT_AMPL_WIDTH),
		3239 => to_signed(10013, LUT_AMPL_WIDTH),
		3240 => to_signed(10016, LUT_AMPL_WIDTH),
		3241 => to_signed(10019, LUT_AMPL_WIDTH),
		3242 => to_signed(10022, LUT_AMPL_WIDTH),
		3243 => to_signed(10025, LUT_AMPL_WIDTH),
		3244 => to_signed(10028, LUT_AMPL_WIDTH),
		3245 => to_signed(10031, LUT_AMPL_WIDTH),
		3246 => to_signed(10033, LUT_AMPL_WIDTH),
		3247 => to_signed(10036, LUT_AMPL_WIDTH),
		3248 => to_signed(10039, LUT_AMPL_WIDTH),
		3249 => to_signed(10042, LUT_AMPL_WIDTH),
		3250 => to_signed(10045, LUT_AMPL_WIDTH),
		3251 => to_signed(10048, LUT_AMPL_WIDTH),
		3252 => to_signed(10051, LUT_AMPL_WIDTH),
		3253 => to_signed(10054, LUT_AMPL_WIDTH),
		3254 => to_signed(10057, LUT_AMPL_WIDTH),
		3255 => to_signed(10060, LUT_AMPL_WIDTH),
		3256 => to_signed(10063, LUT_AMPL_WIDTH),
		3257 => to_signed(10066, LUT_AMPL_WIDTH),
		3258 => to_signed(10069, LUT_AMPL_WIDTH),
		3259 => to_signed(10072, LUT_AMPL_WIDTH),
		3260 => to_signed(10075, LUT_AMPL_WIDTH),
		3261 => to_signed(10078, LUT_AMPL_WIDTH),
		3262 => to_signed(10081, LUT_AMPL_WIDTH),
		3263 => to_signed(10084, LUT_AMPL_WIDTH),
		3264 => to_signed(10087, LUT_AMPL_WIDTH),
		3265 => to_signed(10090, LUT_AMPL_WIDTH),
		3266 => to_signed(10093, LUT_AMPL_WIDTH),
		3267 => to_signed(10096, LUT_AMPL_WIDTH),
		3268 => to_signed(10099, LUT_AMPL_WIDTH),
		3269 => to_signed(10102, LUT_AMPL_WIDTH),
		3270 => to_signed(10105, LUT_AMPL_WIDTH),
		3271 => to_signed(10108, LUT_AMPL_WIDTH),
		3272 => to_signed(10111, LUT_AMPL_WIDTH),
		3273 => to_signed(10114, LUT_AMPL_WIDTH),
		3274 => to_signed(10117, LUT_AMPL_WIDTH),
		3275 => to_signed(10120, LUT_AMPL_WIDTH),
		3276 => to_signed(10123, LUT_AMPL_WIDTH),
		3277 => to_signed(10126, LUT_AMPL_WIDTH),
		3278 => to_signed(10129, LUT_AMPL_WIDTH),
		3279 => to_signed(10132, LUT_AMPL_WIDTH),
		3280 => to_signed(10135, LUT_AMPL_WIDTH),
		3281 => to_signed(10138, LUT_AMPL_WIDTH),
		3282 => to_signed(10141, LUT_AMPL_WIDTH),
		3283 => to_signed(10144, LUT_AMPL_WIDTH),
		3284 => to_signed(10147, LUT_AMPL_WIDTH),
		3285 => to_signed(10150, LUT_AMPL_WIDTH),
		3286 => to_signed(10153, LUT_AMPL_WIDTH),
		3287 => to_signed(10156, LUT_AMPL_WIDTH),
		3288 => to_signed(10159, LUT_AMPL_WIDTH),
		3289 => to_signed(10162, LUT_AMPL_WIDTH),
		3290 => to_signed(10165, LUT_AMPL_WIDTH),
		3291 => to_signed(10168, LUT_AMPL_WIDTH),
		3292 => to_signed(10171, LUT_AMPL_WIDTH),
		3293 => to_signed(10174, LUT_AMPL_WIDTH),
		3294 => to_signed(10177, LUT_AMPL_WIDTH),
		3295 => to_signed(10180, LUT_AMPL_WIDTH),
		3296 => to_signed(10183, LUT_AMPL_WIDTH),
		3297 => to_signed(10186, LUT_AMPL_WIDTH),
		3298 => to_signed(10189, LUT_AMPL_WIDTH),
		3299 => to_signed(10192, LUT_AMPL_WIDTH),
		3300 => to_signed(10195, LUT_AMPL_WIDTH),
		3301 => to_signed(10198, LUT_AMPL_WIDTH),
		3302 => to_signed(10201, LUT_AMPL_WIDTH),
		3303 => to_signed(10204, LUT_AMPL_WIDTH),
		3304 => to_signed(10207, LUT_AMPL_WIDTH),
		3305 => to_signed(10210, LUT_AMPL_WIDTH),
		3306 => to_signed(10213, LUT_AMPL_WIDTH),
		3307 => to_signed(10216, LUT_AMPL_WIDTH),
		3308 => to_signed(10219, LUT_AMPL_WIDTH),
		3309 => to_signed(10222, LUT_AMPL_WIDTH),
		3310 => to_signed(10225, LUT_AMPL_WIDTH),
		3311 => to_signed(10228, LUT_AMPL_WIDTH),
		3312 => to_signed(10231, LUT_AMPL_WIDTH),
		3313 => to_signed(10234, LUT_AMPL_WIDTH),
		3314 => to_signed(10237, LUT_AMPL_WIDTH),
		3315 => to_signed(10240, LUT_AMPL_WIDTH),
		3316 => to_signed(10243, LUT_AMPL_WIDTH),
		3317 => to_signed(10246, LUT_AMPL_WIDTH),
		3318 => to_signed(10249, LUT_AMPL_WIDTH),
		3319 => to_signed(10252, LUT_AMPL_WIDTH),
		3320 => to_signed(10255, LUT_AMPL_WIDTH),
		3321 => to_signed(10258, LUT_AMPL_WIDTH),
		3322 => to_signed(10261, LUT_AMPL_WIDTH),
		3323 => to_signed(10263, LUT_AMPL_WIDTH),
		3324 => to_signed(10266, LUT_AMPL_WIDTH),
		3325 => to_signed(10269, LUT_AMPL_WIDTH),
		3326 => to_signed(10272, LUT_AMPL_WIDTH),
		3327 => to_signed(10275, LUT_AMPL_WIDTH),
		3328 => to_signed(10278, LUT_AMPL_WIDTH),
		3329 => to_signed(10281, LUT_AMPL_WIDTH),
		3330 => to_signed(10284, LUT_AMPL_WIDTH),
		3331 => to_signed(10287, LUT_AMPL_WIDTH),
		3332 => to_signed(10290, LUT_AMPL_WIDTH),
		3333 => to_signed(10293, LUT_AMPL_WIDTH),
		3334 => to_signed(10296, LUT_AMPL_WIDTH),
		3335 => to_signed(10299, LUT_AMPL_WIDTH),
		3336 => to_signed(10302, LUT_AMPL_WIDTH),
		3337 => to_signed(10305, LUT_AMPL_WIDTH),
		3338 => to_signed(10308, LUT_AMPL_WIDTH),
		3339 => to_signed(10311, LUT_AMPL_WIDTH),
		3340 => to_signed(10314, LUT_AMPL_WIDTH),
		3341 => to_signed(10317, LUT_AMPL_WIDTH),
		3342 => to_signed(10320, LUT_AMPL_WIDTH),
		3343 => to_signed(10323, LUT_AMPL_WIDTH),
		3344 => to_signed(10326, LUT_AMPL_WIDTH),
		3345 => to_signed(10329, LUT_AMPL_WIDTH),
		3346 => to_signed(10332, LUT_AMPL_WIDTH),
		3347 => to_signed(10335, LUT_AMPL_WIDTH),
		3348 => to_signed(10338, LUT_AMPL_WIDTH),
		3349 => to_signed(10341, LUT_AMPL_WIDTH),
		3350 => to_signed(10344, LUT_AMPL_WIDTH),
		3351 => to_signed(10347, LUT_AMPL_WIDTH),
		3352 => to_signed(10350, LUT_AMPL_WIDTH),
		3353 => to_signed(10353, LUT_AMPL_WIDTH),
		3354 => to_signed(10356, LUT_AMPL_WIDTH),
		3355 => to_signed(10359, LUT_AMPL_WIDTH),
		3356 => to_signed(10362, LUT_AMPL_WIDTH),
		3357 => to_signed(10365, LUT_AMPL_WIDTH),
		3358 => to_signed(10368, LUT_AMPL_WIDTH),
		3359 => to_signed(10371, LUT_AMPL_WIDTH),
		3360 => to_signed(10374, LUT_AMPL_WIDTH),
		3361 => to_signed(10377, LUT_AMPL_WIDTH),
		3362 => to_signed(10380, LUT_AMPL_WIDTH),
		3363 => to_signed(10383, LUT_AMPL_WIDTH),
		3364 => to_signed(10386, LUT_AMPL_WIDTH),
		3365 => to_signed(10389, LUT_AMPL_WIDTH),
		3366 => to_signed(10392, LUT_AMPL_WIDTH),
		3367 => to_signed(10395, LUT_AMPL_WIDTH),
		3368 => to_signed(10398, LUT_AMPL_WIDTH),
		3369 => to_signed(10401, LUT_AMPL_WIDTH),
		3370 => to_signed(10404, LUT_AMPL_WIDTH),
		3371 => to_signed(10407, LUT_AMPL_WIDTH),
		3372 => to_signed(10410, LUT_AMPL_WIDTH),
		3373 => to_signed(10413, LUT_AMPL_WIDTH),
		3374 => to_signed(10416, LUT_AMPL_WIDTH),
		3375 => to_signed(10419, LUT_AMPL_WIDTH),
		3376 => to_signed(10421, LUT_AMPL_WIDTH),
		3377 => to_signed(10424, LUT_AMPL_WIDTH),
		3378 => to_signed(10427, LUT_AMPL_WIDTH),
		3379 => to_signed(10430, LUT_AMPL_WIDTH),
		3380 => to_signed(10433, LUT_AMPL_WIDTH),
		3381 => to_signed(10436, LUT_AMPL_WIDTH),
		3382 => to_signed(10439, LUT_AMPL_WIDTH),
		3383 => to_signed(10442, LUT_AMPL_WIDTH),
		3384 => to_signed(10445, LUT_AMPL_WIDTH),
		3385 => to_signed(10448, LUT_AMPL_WIDTH),
		3386 => to_signed(10451, LUT_AMPL_WIDTH),
		3387 => to_signed(10454, LUT_AMPL_WIDTH),
		3388 => to_signed(10457, LUT_AMPL_WIDTH),
		3389 => to_signed(10460, LUT_AMPL_WIDTH),
		3390 => to_signed(10463, LUT_AMPL_WIDTH),
		3391 => to_signed(10466, LUT_AMPL_WIDTH),
		3392 => to_signed(10469, LUT_AMPL_WIDTH),
		3393 => to_signed(10472, LUT_AMPL_WIDTH),
		3394 => to_signed(10475, LUT_AMPL_WIDTH),
		3395 => to_signed(10478, LUT_AMPL_WIDTH),
		3396 => to_signed(10481, LUT_AMPL_WIDTH),
		3397 => to_signed(10484, LUT_AMPL_WIDTH),
		3398 => to_signed(10487, LUT_AMPL_WIDTH),
		3399 => to_signed(10490, LUT_AMPL_WIDTH),
		3400 => to_signed(10493, LUT_AMPL_WIDTH),
		3401 => to_signed(10496, LUT_AMPL_WIDTH),
		3402 => to_signed(10499, LUT_AMPL_WIDTH),
		3403 => to_signed(10502, LUT_AMPL_WIDTH),
		3404 => to_signed(10505, LUT_AMPL_WIDTH),
		3405 => to_signed(10508, LUT_AMPL_WIDTH),
		3406 => to_signed(10511, LUT_AMPL_WIDTH),
		3407 => to_signed(10514, LUT_AMPL_WIDTH),
		3408 => to_signed(10517, LUT_AMPL_WIDTH),
		3409 => to_signed(10520, LUT_AMPL_WIDTH),
		3410 => to_signed(10523, LUT_AMPL_WIDTH),
		3411 => to_signed(10526, LUT_AMPL_WIDTH),
		3412 => to_signed(10529, LUT_AMPL_WIDTH),
		3413 => to_signed(10532, LUT_AMPL_WIDTH),
		3414 => to_signed(10535, LUT_AMPL_WIDTH),
		3415 => to_signed(10538, LUT_AMPL_WIDTH),
		3416 => to_signed(10541, LUT_AMPL_WIDTH),
		3417 => to_signed(10544, LUT_AMPL_WIDTH),
		3418 => to_signed(10546, LUT_AMPL_WIDTH),
		3419 => to_signed(10549, LUT_AMPL_WIDTH),
		3420 => to_signed(10552, LUT_AMPL_WIDTH),
		3421 => to_signed(10555, LUT_AMPL_WIDTH),
		3422 => to_signed(10558, LUT_AMPL_WIDTH),
		3423 => to_signed(10561, LUT_AMPL_WIDTH),
		3424 => to_signed(10564, LUT_AMPL_WIDTH),
		3425 => to_signed(10567, LUT_AMPL_WIDTH),
		3426 => to_signed(10570, LUT_AMPL_WIDTH),
		3427 => to_signed(10573, LUT_AMPL_WIDTH),
		3428 => to_signed(10576, LUT_AMPL_WIDTH),
		3429 => to_signed(10579, LUT_AMPL_WIDTH),
		3430 => to_signed(10582, LUT_AMPL_WIDTH),
		3431 => to_signed(10585, LUT_AMPL_WIDTH),
		3432 => to_signed(10588, LUT_AMPL_WIDTH),
		3433 => to_signed(10591, LUT_AMPL_WIDTH),
		3434 => to_signed(10594, LUT_AMPL_WIDTH),
		3435 => to_signed(10597, LUT_AMPL_WIDTH),
		3436 => to_signed(10600, LUT_AMPL_WIDTH),
		3437 => to_signed(10603, LUT_AMPL_WIDTH),
		3438 => to_signed(10606, LUT_AMPL_WIDTH),
		3439 => to_signed(10609, LUT_AMPL_WIDTH),
		3440 => to_signed(10612, LUT_AMPL_WIDTH),
		3441 => to_signed(10615, LUT_AMPL_WIDTH),
		3442 => to_signed(10618, LUT_AMPL_WIDTH),
		3443 => to_signed(10621, LUT_AMPL_WIDTH),
		3444 => to_signed(10624, LUT_AMPL_WIDTH),
		3445 => to_signed(10627, LUT_AMPL_WIDTH),
		3446 => to_signed(10630, LUT_AMPL_WIDTH),
		3447 => to_signed(10633, LUT_AMPL_WIDTH),
		3448 => to_signed(10636, LUT_AMPL_WIDTH),
		3449 => to_signed(10639, LUT_AMPL_WIDTH),
		3450 => to_signed(10642, LUT_AMPL_WIDTH),
		3451 => to_signed(10645, LUT_AMPL_WIDTH),
		3452 => to_signed(10648, LUT_AMPL_WIDTH),
		3453 => to_signed(10651, LUT_AMPL_WIDTH),
		3454 => to_signed(10654, LUT_AMPL_WIDTH),
		3455 => to_signed(10656, LUT_AMPL_WIDTH),
		3456 => to_signed(10659, LUT_AMPL_WIDTH),
		3457 => to_signed(10662, LUT_AMPL_WIDTH),
		3458 => to_signed(10665, LUT_AMPL_WIDTH),
		3459 => to_signed(10668, LUT_AMPL_WIDTH),
		3460 => to_signed(10671, LUT_AMPL_WIDTH),
		3461 => to_signed(10674, LUT_AMPL_WIDTH),
		3462 => to_signed(10677, LUT_AMPL_WIDTH),
		3463 => to_signed(10680, LUT_AMPL_WIDTH),
		3464 => to_signed(10683, LUT_AMPL_WIDTH),
		3465 => to_signed(10686, LUT_AMPL_WIDTH),
		3466 => to_signed(10689, LUT_AMPL_WIDTH),
		3467 => to_signed(10692, LUT_AMPL_WIDTH),
		3468 => to_signed(10695, LUT_AMPL_WIDTH),
		3469 => to_signed(10698, LUT_AMPL_WIDTH),
		3470 => to_signed(10701, LUT_AMPL_WIDTH),
		3471 => to_signed(10704, LUT_AMPL_WIDTH),
		3472 => to_signed(10707, LUT_AMPL_WIDTH),
		3473 => to_signed(10710, LUT_AMPL_WIDTH),
		3474 => to_signed(10713, LUT_AMPL_WIDTH),
		3475 => to_signed(10716, LUT_AMPL_WIDTH),
		3476 => to_signed(10719, LUT_AMPL_WIDTH),
		3477 => to_signed(10722, LUT_AMPL_WIDTH),
		3478 => to_signed(10725, LUT_AMPL_WIDTH),
		3479 => to_signed(10728, LUT_AMPL_WIDTH),
		3480 => to_signed(10731, LUT_AMPL_WIDTH),
		3481 => to_signed(10734, LUT_AMPL_WIDTH),
		3482 => to_signed(10737, LUT_AMPL_WIDTH),
		3483 => to_signed(10740, LUT_AMPL_WIDTH),
		3484 => to_signed(10743, LUT_AMPL_WIDTH),
		3485 => to_signed(10746, LUT_AMPL_WIDTH),
		3486 => to_signed(10749, LUT_AMPL_WIDTH),
		3487 => to_signed(10751, LUT_AMPL_WIDTH),
		3488 => to_signed(10754, LUT_AMPL_WIDTH),
		3489 => to_signed(10757, LUT_AMPL_WIDTH),
		3490 => to_signed(10760, LUT_AMPL_WIDTH),
		3491 => to_signed(10763, LUT_AMPL_WIDTH),
		3492 => to_signed(10766, LUT_AMPL_WIDTH),
		3493 => to_signed(10769, LUT_AMPL_WIDTH),
		3494 => to_signed(10772, LUT_AMPL_WIDTH),
		3495 => to_signed(10775, LUT_AMPL_WIDTH),
		3496 => to_signed(10778, LUT_AMPL_WIDTH),
		3497 => to_signed(10781, LUT_AMPL_WIDTH),
		3498 => to_signed(10784, LUT_AMPL_WIDTH),
		3499 => to_signed(10787, LUT_AMPL_WIDTH),
		3500 => to_signed(10790, LUT_AMPL_WIDTH),
		3501 => to_signed(10793, LUT_AMPL_WIDTH),
		3502 => to_signed(10796, LUT_AMPL_WIDTH),
		3503 => to_signed(10799, LUT_AMPL_WIDTH),
		3504 => to_signed(10802, LUT_AMPL_WIDTH),
		3505 => to_signed(10805, LUT_AMPL_WIDTH),
		3506 => to_signed(10808, LUT_AMPL_WIDTH),
		3507 => to_signed(10811, LUT_AMPL_WIDTH),
		3508 => to_signed(10814, LUT_AMPL_WIDTH),
		3509 => to_signed(10817, LUT_AMPL_WIDTH),
		3510 => to_signed(10820, LUT_AMPL_WIDTH),
		3511 => to_signed(10823, LUT_AMPL_WIDTH),
		3512 => to_signed(10826, LUT_AMPL_WIDTH),
		3513 => to_signed(10829, LUT_AMPL_WIDTH),
		3514 => to_signed(10832, LUT_AMPL_WIDTH),
		3515 => to_signed(10835, LUT_AMPL_WIDTH),
		3516 => to_signed(10838, LUT_AMPL_WIDTH),
		3517 => to_signed(10840, LUT_AMPL_WIDTH),
		3518 => to_signed(10843, LUT_AMPL_WIDTH),
		3519 => to_signed(10846, LUT_AMPL_WIDTH),
		3520 => to_signed(10849, LUT_AMPL_WIDTH),
		3521 => to_signed(10852, LUT_AMPL_WIDTH),
		3522 => to_signed(10855, LUT_AMPL_WIDTH),
		3523 => to_signed(10858, LUT_AMPL_WIDTH),
		3524 => to_signed(10861, LUT_AMPL_WIDTH),
		3525 => to_signed(10864, LUT_AMPL_WIDTH),
		3526 => to_signed(10867, LUT_AMPL_WIDTH),
		3527 => to_signed(10870, LUT_AMPL_WIDTH),
		3528 => to_signed(10873, LUT_AMPL_WIDTH),
		3529 => to_signed(10876, LUT_AMPL_WIDTH),
		3530 => to_signed(10879, LUT_AMPL_WIDTH),
		3531 => to_signed(10882, LUT_AMPL_WIDTH),
		3532 => to_signed(10885, LUT_AMPL_WIDTH),
		3533 => to_signed(10888, LUT_AMPL_WIDTH),
		3534 => to_signed(10891, LUT_AMPL_WIDTH),
		3535 => to_signed(10894, LUT_AMPL_WIDTH),
		3536 => to_signed(10897, LUT_AMPL_WIDTH),
		3537 => to_signed(10900, LUT_AMPL_WIDTH),
		3538 => to_signed(10903, LUT_AMPL_WIDTH),
		3539 => to_signed(10906, LUT_AMPL_WIDTH),
		3540 => to_signed(10909, LUT_AMPL_WIDTH),
		3541 => to_signed(10912, LUT_AMPL_WIDTH),
		3542 => to_signed(10915, LUT_AMPL_WIDTH),
		3543 => to_signed(10918, LUT_AMPL_WIDTH),
		3544 => to_signed(10920, LUT_AMPL_WIDTH),
		3545 => to_signed(10923, LUT_AMPL_WIDTH),
		3546 => to_signed(10926, LUT_AMPL_WIDTH),
		3547 => to_signed(10929, LUT_AMPL_WIDTH),
		3548 => to_signed(10932, LUT_AMPL_WIDTH),
		3549 => to_signed(10935, LUT_AMPL_WIDTH),
		3550 => to_signed(10938, LUT_AMPL_WIDTH),
		3551 => to_signed(10941, LUT_AMPL_WIDTH),
		3552 => to_signed(10944, LUT_AMPL_WIDTH),
		3553 => to_signed(10947, LUT_AMPL_WIDTH),
		3554 => to_signed(10950, LUT_AMPL_WIDTH),
		3555 => to_signed(10953, LUT_AMPL_WIDTH),
		3556 => to_signed(10956, LUT_AMPL_WIDTH),
		3557 => to_signed(10959, LUT_AMPL_WIDTH),
		3558 => to_signed(10962, LUT_AMPL_WIDTH),
		3559 => to_signed(10965, LUT_AMPL_WIDTH),
		3560 => to_signed(10968, LUT_AMPL_WIDTH),
		3561 => to_signed(10971, LUT_AMPL_WIDTH),
		3562 => to_signed(10974, LUT_AMPL_WIDTH),
		3563 => to_signed(10977, LUT_AMPL_WIDTH),
		3564 => to_signed(10980, LUT_AMPL_WIDTH),
		3565 => to_signed(10983, LUT_AMPL_WIDTH),
		3566 => to_signed(10986, LUT_AMPL_WIDTH),
		3567 => to_signed(10989, LUT_AMPL_WIDTH),
		3568 => to_signed(10992, LUT_AMPL_WIDTH),
		3569 => to_signed(10994, LUT_AMPL_WIDTH),
		3570 => to_signed(10997, LUT_AMPL_WIDTH),
		3571 => to_signed(11000, LUT_AMPL_WIDTH),
		3572 => to_signed(11003, LUT_AMPL_WIDTH),
		3573 => to_signed(11006, LUT_AMPL_WIDTH),
		3574 => to_signed(11009, LUT_AMPL_WIDTH),
		3575 => to_signed(11012, LUT_AMPL_WIDTH),
		3576 => to_signed(11015, LUT_AMPL_WIDTH),
		3577 => to_signed(11018, LUT_AMPL_WIDTH),
		3578 => to_signed(11021, LUT_AMPL_WIDTH),
		3579 => to_signed(11024, LUT_AMPL_WIDTH),
		3580 => to_signed(11027, LUT_AMPL_WIDTH),
		3581 => to_signed(11030, LUT_AMPL_WIDTH),
		3582 => to_signed(11033, LUT_AMPL_WIDTH),
		3583 => to_signed(11036, LUT_AMPL_WIDTH),
		3584 => to_signed(11039, LUT_AMPL_WIDTH),
		3585 => to_signed(11042, LUT_AMPL_WIDTH),
		3586 => to_signed(11045, LUT_AMPL_WIDTH),
		3587 => to_signed(11048, LUT_AMPL_WIDTH),
		3588 => to_signed(11051, LUT_AMPL_WIDTH),
		3589 => to_signed(11054, LUT_AMPL_WIDTH),
		3590 => to_signed(11057, LUT_AMPL_WIDTH),
		3591 => to_signed(11060, LUT_AMPL_WIDTH),
		3592 => to_signed(11063, LUT_AMPL_WIDTH),
		3593 => to_signed(11065, LUT_AMPL_WIDTH),
		3594 => to_signed(11068, LUT_AMPL_WIDTH),
		3595 => to_signed(11071, LUT_AMPL_WIDTH),
		3596 => to_signed(11074, LUT_AMPL_WIDTH),
		3597 => to_signed(11077, LUT_AMPL_WIDTH),
		3598 => to_signed(11080, LUT_AMPL_WIDTH),
		3599 => to_signed(11083, LUT_AMPL_WIDTH),
		3600 => to_signed(11086, LUT_AMPL_WIDTH),
		3601 => to_signed(11089, LUT_AMPL_WIDTH),
		3602 => to_signed(11092, LUT_AMPL_WIDTH),
		3603 => to_signed(11095, LUT_AMPL_WIDTH),
		3604 => to_signed(11098, LUT_AMPL_WIDTH),
		3605 => to_signed(11101, LUT_AMPL_WIDTH),
		3606 => to_signed(11104, LUT_AMPL_WIDTH),
		3607 => to_signed(11107, LUT_AMPL_WIDTH),
		3608 => to_signed(11110, LUT_AMPL_WIDTH),
		3609 => to_signed(11113, LUT_AMPL_WIDTH),
		3610 => to_signed(11116, LUT_AMPL_WIDTH),
		3611 => to_signed(11119, LUT_AMPL_WIDTH),
		3612 => to_signed(11122, LUT_AMPL_WIDTH),
		3613 => to_signed(11125, LUT_AMPL_WIDTH),
		3614 => to_signed(11128, LUT_AMPL_WIDTH),
		3615 => to_signed(11131, LUT_AMPL_WIDTH),
		3616 => to_signed(11133, LUT_AMPL_WIDTH),
		3617 => to_signed(11136, LUT_AMPL_WIDTH),
		3618 => to_signed(11139, LUT_AMPL_WIDTH),
		3619 => to_signed(11142, LUT_AMPL_WIDTH),
		3620 => to_signed(11145, LUT_AMPL_WIDTH),
		3621 => to_signed(11148, LUT_AMPL_WIDTH),
		3622 => to_signed(11151, LUT_AMPL_WIDTH),
		3623 => to_signed(11154, LUT_AMPL_WIDTH),
		3624 => to_signed(11157, LUT_AMPL_WIDTH),
		3625 => to_signed(11160, LUT_AMPL_WIDTH),
		3626 => to_signed(11163, LUT_AMPL_WIDTH),
		3627 => to_signed(11166, LUT_AMPL_WIDTH),
		3628 => to_signed(11169, LUT_AMPL_WIDTH),
		3629 => to_signed(11172, LUT_AMPL_WIDTH),
		3630 => to_signed(11175, LUT_AMPL_WIDTH),
		3631 => to_signed(11178, LUT_AMPL_WIDTH),
		3632 => to_signed(11181, LUT_AMPL_WIDTH),
		3633 => to_signed(11184, LUT_AMPL_WIDTH),
		3634 => to_signed(11187, LUT_AMPL_WIDTH),
		3635 => to_signed(11190, LUT_AMPL_WIDTH),
		3636 => to_signed(11193, LUT_AMPL_WIDTH),
		3637 => to_signed(11195, LUT_AMPL_WIDTH),
		3638 => to_signed(11198, LUT_AMPL_WIDTH),
		3639 => to_signed(11201, LUT_AMPL_WIDTH),
		3640 => to_signed(11204, LUT_AMPL_WIDTH),
		3641 => to_signed(11207, LUT_AMPL_WIDTH),
		3642 => to_signed(11210, LUT_AMPL_WIDTH),
		3643 => to_signed(11213, LUT_AMPL_WIDTH),
		3644 => to_signed(11216, LUT_AMPL_WIDTH),
		3645 => to_signed(11219, LUT_AMPL_WIDTH),
		3646 => to_signed(11222, LUT_AMPL_WIDTH),
		3647 => to_signed(11225, LUT_AMPL_WIDTH),
		3648 => to_signed(11228, LUT_AMPL_WIDTH),
		3649 => to_signed(11231, LUT_AMPL_WIDTH),
		3650 => to_signed(11234, LUT_AMPL_WIDTH),
		3651 => to_signed(11237, LUT_AMPL_WIDTH),
		3652 => to_signed(11240, LUT_AMPL_WIDTH),
		3653 => to_signed(11243, LUT_AMPL_WIDTH),
		3654 => to_signed(11246, LUT_AMPL_WIDTH),
		3655 => to_signed(11249, LUT_AMPL_WIDTH),
		3656 => to_signed(11252, LUT_AMPL_WIDTH),
		3657 => to_signed(11255, LUT_AMPL_WIDTH),
		3658 => to_signed(11257, LUT_AMPL_WIDTH),
		3659 => to_signed(11260, LUT_AMPL_WIDTH),
		3660 => to_signed(11263, LUT_AMPL_WIDTH),
		3661 => to_signed(11266, LUT_AMPL_WIDTH),
		3662 => to_signed(11269, LUT_AMPL_WIDTH),
		3663 => to_signed(11272, LUT_AMPL_WIDTH),
		3664 => to_signed(11275, LUT_AMPL_WIDTH),
		3665 => to_signed(11278, LUT_AMPL_WIDTH),
		3666 => to_signed(11281, LUT_AMPL_WIDTH),
		3667 => to_signed(11284, LUT_AMPL_WIDTH),
		3668 => to_signed(11287, LUT_AMPL_WIDTH),
		3669 => to_signed(11290, LUT_AMPL_WIDTH),
		3670 => to_signed(11293, LUT_AMPL_WIDTH),
		3671 => to_signed(11296, LUT_AMPL_WIDTH),
		3672 => to_signed(11299, LUT_AMPL_WIDTH),
		3673 => to_signed(11302, LUT_AMPL_WIDTH),
		3674 => to_signed(11305, LUT_AMPL_WIDTH),
		3675 => to_signed(11308, LUT_AMPL_WIDTH),
		3676 => to_signed(11311, LUT_AMPL_WIDTH),
		3677 => to_signed(11314, LUT_AMPL_WIDTH),
		3678 => to_signed(11316, LUT_AMPL_WIDTH),
		3679 => to_signed(11319, LUT_AMPL_WIDTH),
		3680 => to_signed(11322, LUT_AMPL_WIDTH),
		3681 => to_signed(11325, LUT_AMPL_WIDTH),
		3682 => to_signed(11328, LUT_AMPL_WIDTH),
		3683 => to_signed(11331, LUT_AMPL_WIDTH),
		3684 => to_signed(11334, LUT_AMPL_WIDTH),
		3685 => to_signed(11337, LUT_AMPL_WIDTH),
		3686 => to_signed(11340, LUT_AMPL_WIDTH),
		3687 => to_signed(11343, LUT_AMPL_WIDTH),
		3688 => to_signed(11346, LUT_AMPL_WIDTH),
		3689 => to_signed(11349, LUT_AMPL_WIDTH),
		3690 => to_signed(11352, LUT_AMPL_WIDTH),
		3691 => to_signed(11355, LUT_AMPL_WIDTH),
		3692 => to_signed(11358, LUT_AMPL_WIDTH),
		3693 => to_signed(11361, LUT_AMPL_WIDTH),
		3694 => to_signed(11364, LUT_AMPL_WIDTH),
		3695 => to_signed(11367, LUT_AMPL_WIDTH),
		3696 => to_signed(11370, LUT_AMPL_WIDTH),
		3697 => to_signed(11372, LUT_AMPL_WIDTH),
		3698 => to_signed(11375, LUT_AMPL_WIDTH),
		3699 => to_signed(11378, LUT_AMPL_WIDTH),
		3700 => to_signed(11381, LUT_AMPL_WIDTH),
		3701 => to_signed(11384, LUT_AMPL_WIDTH),
		3702 => to_signed(11387, LUT_AMPL_WIDTH),
		3703 => to_signed(11390, LUT_AMPL_WIDTH),
		3704 => to_signed(11393, LUT_AMPL_WIDTH),
		3705 => to_signed(11396, LUT_AMPL_WIDTH),
		3706 => to_signed(11399, LUT_AMPL_WIDTH),
		3707 => to_signed(11402, LUT_AMPL_WIDTH),
		3708 => to_signed(11405, LUT_AMPL_WIDTH),
		3709 => to_signed(11408, LUT_AMPL_WIDTH),
		3710 => to_signed(11411, LUT_AMPL_WIDTH),
		3711 => to_signed(11414, LUT_AMPL_WIDTH),
		3712 => to_signed(11417, LUT_AMPL_WIDTH),
		3713 => to_signed(11420, LUT_AMPL_WIDTH),
		3714 => to_signed(11423, LUT_AMPL_WIDTH),
		3715 => to_signed(11425, LUT_AMPL_WIDTH),
		3716 => to_signed(11428, LUT_AMPL_WIDTH),
		3717 => to_signed(11431, LUT_AMPL_WIDTH),
		3718 => to_signed(11434, LUT_AMPL_WIDTH),
		3719 => to_signed(11437, LUT_AMPL_WIDTH),
		3720 => to_signed(11440, LUT_AMPL_WIDTH),
		3721 => to_signed(11443, LUT_AMPL_WIDTH),
		3722 => to_signed(11446, LUT_AMPL_WIDTH),
		3723 => to_signed(11449, LUT_AMPL_WIDTH),
		3724 => to_signed(11452, LUT_AMPL_WIDTH),
		3725 => to_signed(11455, LUT_AMPL_WIDTH),
		3726 => to_signed(11458, LUT_AMPL_WIDTH),
		3727 => to_signed(11461, LUT_AMPL_WIDTH),
		3728 => to_signed(11464, LUT_AMPL_WIDTH),
		3729 => to_signed(11467, LUT_AMPL_WIDTH),
		3730 => to_signed(11470, LUT_AMPL_WIDTH),
		3731 => to_signed(11473, LUT_AMPL_WIDTH),
		3732 => to_signed(11476, LUT_AMPL_WIDTH),
		3733 => to_signed(11478, LUT_AMPL_WIDTH),
		3734 => to_signed(11481, LUT_AMPL_WIDTH),
		3735 => to_signed(11484, LUT_AMPL_WIDTH),
		3736 => to_signed(11487, LUT_AMPL_WIDTH),
		3737 => to_signed(11490, LUT_AMPL_WIDTH),
		3738 => to_signed(11493, LUT_AMPL_WIDTH),
		3739 => to_signed(11496, LUT_AMPL_WIDTH),
		3740 => to_signed(11499, LUT_AMPL_WIDTH),
		3741 => to_signed(11502, LUT_AMPL_WIDTH),
		3742 => to_signed(11505, LUT_AMPL_WIDTH),
		3743 => to_signed(11508, LUT_AMPL_WIDTH),
		3744 => to_signed(11511, LUT_AMPL_WIDTH),
		3745 => to_signed(11514, LUT_AMPL_WIDTH),
		3746 => to_signed(11517, LUT_AMPL_WIDTH),
		3747 => to_signed(11520, LUT_AMPL_WIDTH),
		3748 => to_signed(11523, LUT_AMPL_WIDTH),
		3749 => to_signed(11526, LUT_AMPL_WIDTH),
		3750 => to_signed(11528, LUT_AMPL_WIDTH),
		3751 => to_signed(11531, LUT_AMPL_WIDTH),
		3752 => to_signed(11534, LUT_AMPL_WIDTH),
		3753 => to_signed(11537, LUT_AMPL_WIDTH),
		3754 => to_signed(11540, LUT_AMPL_WIDTH),
		3755 => to_signed(11543, LUT_AMPL_WIDTH),
		3756 => to_signed(11546, LUT_AMPL_WIDTH),
		3757 => to_signed(11549, LUT_AMPL_WIDTH),
		3758 => to_signed(11552, LUT_AMPL_WIDTH),
		3759 => to_signed(11555, LUT_AMPL_WIDTH),
		3760 => to_signed(11558, LUT_AMPL_WIDTH),
		3761 => to_signed(11561, LUT_AMPL_WIDTH),
		3762 => to_signed(11564, LUT_AMPL_WIDTH),
		3763 => to_signed(11567, LUT_AMPL_WIDTH),
		3764 => to_signed(11570, LUT_AMPL_WIDTH),
		3765 => to_signed(11573, LUT_AMPL_WIDTH),
		3766 => to_signed(11575, LUT_AMPL_WIDTH),
		3767 => to_signed(11578, LUT_AMPL_WIDTH),
		3768 => to_signed(11581, LUT_AMPL_WIDTH),
		3769 => to_signed(11584, LUT_AMPL_WIDTH),
		3770 => to_signed(11587, LUT_AMPL_WIDTH),
		3771 => to_signed(11590, LUT_AMPL_WIDTH),
		3772 => to_signed(11593, LUT_AMPL_WIDTH),
		3773 => to_signed(11596, LUT_AMPL_WIDTH),
		3774 => to_signed(11599, LUT_AMPL_WIDTH),
		3775 => to_signed(11602, LUT_AMPL_WIDTH),
		3776 => to_signed(11605, LUT_AMPL_WIDTH),
		3777 => to_signed(11608, LUT_AMPL_WIDTH),
		3778 => to_signed(11611, LUT_AMPL_WIDTH),
		3779 => to_signed(11614, LUT_AMPL_WIDTH),
		3780 => to_signed(11617, LUT_AMPL_WIDTH),
		3781 => to_signed(11620, LUT_AMPL_WIDTH),
		3782 => to_signed(11623, LUT_AMPL_WIDTH),
		3783 => to_signed(11625, LUT_AMPL_WIDTH),
		3784 => to_signed(11628, LUT_AMPL_WIDTH),
		3785 => to_signed(11631, LUT_AMPL_WIDTH),
		3786 => to_signed(11634, LUT_AMPL_WIDTH),
		3787 => to_signed(11637, LUT_AMPL_WIDTH),
		3788 => to_signed(11640, LUT_AMPL_WIDTH),
		3789 => to_signed(11643, LUT_AMPL_WIDTH),
		3790 => to_signed(11646, LUT_AMPL_WIDTH),
		3791 => to_signed(11649, LUT_AMPL_WIDTH),
		3792 => to_signed(11652, LUT_AMPL_WIDTH),
		3793 => to_signed(11655, LUT_AMPL_WIDTH),
		3794 => to_signed(11658, LUT_AMPL_WIDTH),
		3795 => to_signed(11661, LUT_AMPL_WIDTH),
		3796 => to_signed(11664, LUT_AMPL_WIDTH),
		3797 => to_signed(11667, LUT_AMPL_WIDTH),
		3798 => to_signed(11669, LUT_AMPL_WIDTH),
		3799 => to_signed(11672, LUT_AMPL_WIDTH),
		3800 => to_signed(11675, LUT_AMPL_WIDTH),
		3801 => to_signed(11678, LUT_AMPL_WIDTH),
		3802 => to_signed(11681, LUT_AMPL_WIDTH),
		3803 => to_signed(11684, LUT_AMPL_WIDTH),
		3804 => to_signed(11687, LUT_AMPL_WIDTH),
		3805 => to_signed(11690, LUT_AMPL_WIDTH),
		3806 => to_signed(11693, LUT_AMPL_WIDTH),
		3807 => to_signed(11696, LUT_AMPL_WIDTH),
		3808 => to_signed(11699, LUT_AMPL_WIDTH),
		3809 => to_signed(11702, LUT_AMPL_WIDTH),
		3810 => to_signed(11705, LUT_AMPL_WIDTH),
		3811 => to_signed(11708, LUT_AMPL_WIDTH),
		3812 => to_signed(11711, LUT_AMPL_WIDTH),
		3813 => to_signed(11714, LUT_AMPL_WIDTH),
		3814 => to_signed(11716, LUT_AMPL_WIDTH),
		3815 => to_signed(11719, LUT_AMPL_WIDTH),
		3816 => to_signed(11722, LUT_AMPL_WIDTH),
		3817 => to_signed(11725, LUT_AMPL_WIDTH),
		3818 => to_signed(11728, LUT_AMPL_WIDTH),
		3819 => to_signed(11731, LUT_AMPL_WIDTH),
		3820 => to_signed(11734, LUT_AMPL_WIDTH),
		3821 => to_signed(11737, LUT_AMPL_WIDTH),
		3822 => to_signed(11740, LUT_AMPL_WIDTH),
		3823 => to_signed(11743, LUT_AMPL_WIDTH),
		3824 => to_signed(11746, LUT_AMPL_WIDTH),
		3825 => to_signed(11749, LUT_AMPL_WIDTH),
		3826 => to_signed(11752, LUT_AMPL_WIDTH),
		3827 => to_signed(11755, LUT_AMPL_WIDTH),
		3828 => to_signed(11758, LUT_AMPL_WIDTH),
		3829 => to_signed(11760, LUT_AMPL_WIDTH),
		3830 => to_signed(11763, LUT_AMPL_WIDTH),
		3831 => to_signed(11766, LUT_AMPL_WIDTH),
		3832 => to_signed(11769, LUT_AMPL_WIDTH),
		3833 => to_signed(11772, LUT_AMPL_WIDTH),
		3834 => to_signed(11775, LUT_AMPL_WIDTH),
		3835 => to_signed(11778, LUT_AMPL_WIDTH),
		3836 => to_signed(11781, LUT_AMPL_WIDTH),
		3837 => to_signed(11784, LUT_AMPL_WIDTH),
		3838 => to_signed(11787, LUT_AMPL_WIDTH),
		3839 => to_signed(11790, LUT_AMPL_WIDTH),
		3840 => to_signed(11793, LUT_AMPL_WIDTH),
		3841 => to_signed(11796, LUT_AMPL_WIDTH),
		3842 => to_signed(11799, LUT_AMPL_WIDTH),
		3843 => to_signed(11801, LUT_AMPL_WIDTH),
		3844 => to_signed(11804, LUT_AMPL_WIDTH),
		3845 => to_signed(11807, LUT_AMPL_WIDTH),
		3846 => to_signed(11810, LUT_AMPL_WIDTH),
		3847 => to_signed(11813, LUT_AMPL_WIDTH),
		3848 => to_signed(11816, LUT_AMPL_WIDTH),
		3849 => to_signed(11819, LUT_AMPL_WIDTH),
		3850 => to_signed(11822, LUT_AMPL_WIDTH),
		3851 => to_signed(11825, LUT_AMPL_WIDTH),
		3852 => to_signed(11828, LUT_AMPL_WIDTH),
		3853 => to_signed(11831, LUT_AMPL_WIDTH),
		3854 => to_signed(11834, LUT_AMPL_WIDTH),
		3855 => to_signed(11837, LUT_AMPL_WIDTH),
		3856 => to_signed(11840, LUT_AMPL_WIDTH),
		3857 => to_signed(11842, LUT_AMPL_WIDTH),
		3858 => to_signed(11845, LUT_AMPL_WIDTH),
		3859 => to_signed(11848, LUT_AMPL_WIDTH),
		3860 => to_signed(11851, LUT_AMPL_WIDTH),
		3861 => to_signed(11854, LUT_AMPL_WIDTH),
		3862 => to_signed(11857, LUT_AMPL_WIDTH),
		3863 => to_signed(11860, LUT_AMPL_WIDTH),
		3864 => to_signed(11863, LUT_AMPL_WIDTH),
		3865 => to_signed(11866, LUT_AMPL_WIDTH),
		3866 => to_signed(11869, LUT_AMPL_WIDTH),
		3867 => to_signed(11872, LUT_AMPL_WIDTH),
		3868 => to_signed(11875, LUT_AMPL_WIDTH),
		3869 => to_signed(11878, LUT_AMPL_WIDTH),
		3870 => to_signed(11881, LUT_AMPL_WIDTH),
		3871 => to_signed(11883, LUT_AMPL_WIDTH),
		3872 => to_signed(11886, LUT_AMPL_WIDTH),
		3873 => to_signed(11889, LUT_AMPL_WIDTH),
		3874 => to_signed(11892, LUT_AMPL_WIDTH),
		3875 => to_signed(11895, LUT_AMPL_WIDTH),
		3876 => to_signed(11898, LUT_AMPL_WIDTH),
		3877 => to_signed(11901, LUT_AMPL_WIDTH),
		3878 => to_signed(11904, LUT_AMPL_WIDTH),
		3879 => to_signed(11907, LUT_AMPL_WIDTH),
		3880 => to_signed(11910, LUT_AMPL_WIDTH),
		3881 => to_signed(11913, LUT_AMPL_WIDTH),
		3882 => to_signed(11916, LUT_AMPL_WIDTH),
		3883 => to_signed(11919, LUT_AMPL_WIDTH),
		3884 => to_signed(11922, LUT_AMPL_WIDTH),
		3885 => to_signed(11924, LUT_AMPL_WIDTH),
		3886 => to_signed(11927, LUT_AMPL_WIDTH),
		3887 => to_signed(11930, LUT_AMPL_WIDTH),
		3888 => to_signed(11933, LUT_AMPL_WIDTH),
		3889 => to_signed(11936, LUT_AMPL_WIDTH),
		3890 => to_signed(11939, LUT_AMPL_WIDTH),
		3891 => to_signed(11942, LUT_AMPL_WIDTH),
		3892 => to_signed(11945, LUT_AMPL_WIDTH),
		3893 => to_signed(11948, LUT_AMPL_WIDTH),
		3894 => to_signed(11951, LUT_AMPL_WIDTH),
		3895 => to_signed(11954, LUT_AMPL_WIDTH),
		3896 => to_signed(11957, LUT_AMPL_WIDTH),
		3897 => to_signed(11960, LUT_AMPL_WIDTH),
		3898 => to_signed(11962, LUT_AMPL_WIDTH),
		3899 => to_signed(11965, LUT_AMPL_WIDTH),
		3900 => to_signed(11968, LUT_AMPL_WIDTH),
		3901 => to_signed(11971, LUT_AMPL_WIDTH),
		3902 => to_signed(11974, LUT_AMPL_WIDTH),
		3903 => to_signed(11977, LUT_AMPL_WIDTH),
		3904 => to_signed(11980, LUT_AMPL_WIDTH),
		3905 => to_signed(11983, LUT_AMPL_WIDTH),
		3906 => to_signed(11986, LUT_AMPL_WIDTH),
		3907 => to_signed(11989, LUT_AMPL_WIDTH),
		3908 => to_signed(11992, LUT_AMPL_WIDTH),
		3909 => to_signed(11995, LUT_AMPL_WIDTH),
		3910 => to_signed(11998, LUT_AMPL_WIDTH),
		3911 => to_signed(12001, LUT_AMPL_WIDTH),
		3912 => to_signed(12003, LUT_AMPL_WIDTH),
		3913 => to_signed(12006, LUT_AMPL_WIDTH),
		3914 => to_signed(12009, LUT_AMPL_WIDTH),
		3915 => to_signed(12012, LUT_AMPL_WIDTH),
		3916 => to_signed(12015, LUT_AMPL_WIDTH),
		3917 => to_signed(12018, LUT_AMPL_WIDTH),
		3918 => to_signed(12021, LUT_AMPL_WIDTH),
		3919 => to_signed(12024, LUT_AMPL_WIDTH),
		3920 => to_signed(12027, LUT_AMPL_WIDTH),
		3921 => to_signed(12030, LUT_AMPL_WIDTH),
		3922 => to_signed(12033, LUT_AMPL_WIDTH),
		3923 => to_signed(12036, LUT_AMPL_WIDTH),
		3924 => to_signed(12038, LUT_AMPL_WIDTH),
		3925 => to_signed(12041, LUT_AMPL_WIDTH),
		3926 => to_signed(12044, LUT_AMPL_WIDTH),
		3927 => to_signed(12047, LUT_AMPL_WIDTH),
		3928 => to_signed(12050, LUT_AMPL_WIDTH),
		3929 => to_signed(12053, LUT_AMPL_WIDTH),
		3930 => to_signed(12056, LUT_AMPL_WIDTH),
		3931 => to_signed(12059, LUT_AMPL_WIDTH),
		3932 => to_signed(12062, LUT_AMPL_WIDTH),
		3933 => to_signed(12065, LUT_AMPL_WIDTH),
		3934 => to_signed(12068, LUT_AMPL_WIDTH),
		3935 => to_signed(12071, LUT_AMPL_WIDTH),
		3936 => to_signed(12074, LUT_AMPL_WIDTH),
		3937 => to_signed(12076, LUT_AMPL_WIDTH),
		3938 => to_signed(12079, LUT_AMPL_WIDTH),
		3939 => to_signed(12082, LUT_AMPL_WIDTH),
		3940 => to_signed(12085, LUT_AMPL_WIDTH),
		3941 => to_signed(12088, LUT_AMPL_WIDTH),
		3942 => to_signed(12091, LUT_AMPL_WIDTH),
		3943 => to_signed(12094, LUT_AMPL_WIDTH),
		3944 => to_signed(12097, LUT_AMPL_WIDTH),
		3945 => to_signed(12100, LUT_AMPL_WIDTH),
		3946 => to_signed(12103, LUT_AMPL_WIDTH),
		3947 => to_signed(12106, LUT_AMPL_WIDTH),
		3948 => to_signed(12109, LUT_AMPL_WIDTH),
		3949 => to_signed(12112, LUT_AMPL_WIDTH),
		3950 => to_signed(12114, LUT_AMPL_WIDTH),
		3951 => to_signed(12117, LUT_AMPL_WIDTH),
		3952 => to_signed(12120, LUT_AMPL_WIDTH),
		3953 => to_signed(12123, LUT_AMPL_WIDTH),
		3954 => to_signed(12126, LUT_AMPL_WIDTH),
		3955 => to_signed(12129, LUT_AMPL_WIDTH),
		3956 => to_signed(12132, LUT_AMPL_WIDTH),
		3957 => to_signed(12135, LUT_AMPL_WIDTH),
		3958 => to_signed(12138, LUT_AMPL_WIDTH),
		3959 => to_signed(12141, LUT_AMPL_WIDTH),
		3960 => to_signed(12144, LUT_AMPL_WIDTH),
		3961 => to_signed(12147, LUT_AMPL_WIDTH),
		3962 => to_signed(12149, LUT_AMPL_WIDTH),
		3963 => to_signed(12152, LUT_AMPL_WIDTH),
		3964 => to_signed(12155, LUT_AMPL_WIDTH),
		3965 => to_signed(12158, LUT_AMPL_WIDTH),
		3966 => to_signed(12161, LUT_AMPL_WIDTH),
		3967 => to_signed(12164, LUT_AMPL_WIDTH),
		3968 => to_signed(12167, LUT_AMPL_WIDTH),
		3969 => to_signed(12170, LUT_AMPL_WIDTH),
		3970 => to_signed(12173, LUT_AMPL_WIDTH),
		3971 => to_signed(12176, LUT_AMPL_WIDTH),
		3972 => to_signed(12179, LUT_AMPL_WIDTH),
		3973 => to_signed(12182, LUT_AMPL_WIDTH),
		3974 => to_signed(12184, LUT_AMPL_WIDTH),
		3975 => to_signed(12187, LUT_AMPL_WIDTH),
		3976 => to_signed(12190, LUT_AMPL_WIDTH),
		3977 => to_signed(12193, LUT_AMPL_WIDTH),
		3978 => to_signed(12196, LUT_AMPL_WIDTH),
		3979 => to_signed(12199, LUT_AMPL_WIDTH),
		3980 => to_signed(12202, LUT_AMPL_WIDTH),
		3981 => to_signed(12205, LUT_AMPL_WIDTH),
		3982 => to_signed(12208, LUT_AMPL_WIDTH),
		3983 => to_signed(12211, LUT_AMPL_WIDTH),
		3984 => to_signed(12214, LUT_AMPL_WIDTH),
		3985 => to_signed(12217, LUT_AMPL_WIDTH),
		3986 => to_signed(12219, LUT_AMPL_WIDTH),
		3987 => to_signed(12222, LUT_AMPL_WIDTH),
		3988 => to_signed(12225, LUT_AMPL_WIDTH),
		3989 => to_signed(12228, LUT_AMPL_WIDTH),
		3990 => to_signed(12231, LUT_AMPL_WIDTH),
		3991 => to_signed(12234, LUT_AMPL_WIDTH),
		3992 => to_signed(12237, LUT_AMPL_WIDTH),
		3993 => to_signed(12240, LUT_AMPL_WIDTH),
		3994 => to_signed(12243, LUT_AMPL_WIDTH),
		3995 => to_signed(12246, LUT_AMPL_WIDTH),
		3996 => to_signed(12249, LUT_AMPL_WIDTH),
		3997 => to_signed(12251, LUT_AMPL_WIDTH),
		3998 => to_signed(12254, LUT_AMPL_WIDTH),
		3999 => to_signed(12257, LUT_AMPL_WIDTH),
		4000 => to_signed(12260, LUT_AMPL_WIDTH),
		4001 => to_signed(12263, LUT_AMPL_WIDTH),
		4002 => to_signed(12266, LUT_AMPL_WIDTH),
		4003 => to_signed(12269, LUT_AMPL_WIDTH),
		4004 => to_signed(12272, LUT_AMPL_WIDTH),
		4005 => to_signed(12275, LUT_AMPL_WIDTH),
		4006 => to_signed(12278, LUT_AMPL_WIDTH),
		4007 => to_signed(12281, LUT_AMPL_WIDTH),
		4008 => to_signed(12284, LUT_AMPL_WIDTH),
		4009 => to_signed(12286, LUT_AMPL_WIDTH),
		4010 => to_signed(12289, LUT_AMPL_WIDTH),
		4011 => to_signed(12292, LUT_AMPL_WIDTH),
		4012 => to_signed(12295, LUT_AMPL_WIDTH),
		4013 => to_signed(12298, LUT_AMPL_WIDTH),
		4014 => to_signed(12301, LUT_AMPL_WIDTH),
		4015 => to_signed(12304, LUT_AMPL_WIDTH),
		4016 => to_signed(12307, LUT_AMPL_WIDTH),
		4017 => to_signed(12310, LUT_AMPL_WIDTH),
		4018 => to_signed(12313, LUT_AMPL_WIDTH),
		4019 => to_signed(12316, LUT_AMPL_WIDTH),
		4020 => to_signed(12318, LUT_AMPL_WIDTH),
		4021 => to_signed(12321, LUT_AMPL_WIDTH),
		4022 => to_signed(12324, LUT_AMPL_WIDTH),
		4023 => to_signed(12327, LUT_AMPL_WIDTH),
		4024 => to_signed(12330, LUT_AMPL_WIDTH),
		4025 => to_signed(12333, LUT_AMPL_WIDTH),
		4026 => to_signed(12336, LUT_AMPL_WIDTH),
		4027 => to_signed(12339, LUT_AMPL_WIDTH),
		4028 => to_signed(12342, LUT_AMPL_WIDTH),
		4029 => to_signed(12345, LUT_AMPL_WIDTH),
		4030 => to_signed(12348, LUT_AMPL_WIDTH),
		4031 => to_signed(12350, LUT_AMPL_WIDTH),
		4032 => to_signed(12353, LUT_AMPL_WIDTH),
		4033 => to_signed(12356, LUT_AMPL_WIDTH),
		4034 => to_signed(12359, LUT_AMPL_WIDTH),
		4035 => to_signed(12362, LUT_AMPL_WIDTH),
		4036 => to_signed(12365, LUT_AMPL_WIDTH),
		4037 => to_signed(12368, LUT_AMPL_WIDTH),
		4038 => to_signed(12371, LUT_AMPL_WIDTH),
		4039 => to_signed(12374, LUT_AMPL_WIDTH),
		4040 => to_signed(12377, LUT_AMPL_WIDTH),
		4041 => to_signed(12380, LUT_AMPL_WIDTH),
		4042 => to_signed(12382, LUT_AMPL_WIDTH),
		4043 => to_signed(12385, LUT_AMPL_WIDTH),
		4044 => to_signed(12388, LUT_AMPL_WIDTH),
		4045 => to_signed(12391, LUT_AMPL_WIDTH),
		4046 => to_signed(12394, LUT_AMPL_WIDTH),
		4047 => to_signed(12397, LUT_AMPL_WIDTH),
		4048 => to_signed(12400, LUT_AMPL_WIDTH),
		4049 => to_signed(12403, LUT_AMPL_WIDTH),
		4050 => to_signed(12406, LUT_AMPL_WIDTH),
		4051 => to_signed(12409, LUT_AMPL_WIDTH),
		4052 => to_signed(12412, LUT_AMPL_WIDTH),
		4053 => to_signed(12414, LUT_AMPL_WIDTH),
		4054 => to_signed(12417, LUT_AMPL_WIDTH),
		4055 => to_signed(12420, LUT_AMPL_WIDTH),
		4056 => to_signed(12423, LUT_AMPL_WIDTH),
		4057 => to_signed(12426, LUT_AMPL_WIDTH),
		4058 => to_signed(12429, LUT_AMPL_WIDTH),
		4059 => to_signed(12432, LUT_AMPL_WIDTH),
		4060 => to_signed(12435, LUT_AMPL_WIDTH),
		4061 => to_signed(12438, LUT_AMPL_WIDTH),
		4062 => to_signed(12441, LUT_AMPL_WIDTH),
		4063 => to_signed(12444, LUT_AMPL_WIDTH),
		4064 => to_signed(12446, LUT_AMPL_WIDTH),
		4065 => to_signed(12449, LUT_AMPL_WIDTH),
		4066 => to_signed(12452, LUT_AMPL_WIDTH),
		4067 => to_signed(12455, LUT_AMPL_WIDTH),
		4068 => to_signed(12458, LUT_AMPL_WIDTH),
		4069 => to_signed(12461, LUT_AMPL_WIDTH),
		4070 => to_signed(12464, LUT_AMPL_WIDTH),
		4071 => to_signed(12467, LUT_AMPL_WIDTH),
		4072 => to_signed(12470, LUT_AMPL_WIDTH),
		4073 => to_signed(12473, LUT_AMPL_WIDTH),
		4074 => to_signed(12476, LUT_AMPL_WIDTH),
		4075 => to_signed(12478, LUT_AMPL_WIDTH),
		4076 => to_signed(12481, LUT_AMPL_WIDTH),
		4077 => to_signed(12484, LUT_AMPL_WIDTH),
		4078 => to_signed(12487, LUT_AMPL_WIDTH),
		4079 => to_signed(12490, LUT_AMPL_WIDTH),
		4080 => to_signed(12493, LUT_AMPL_WIDTH),
		4081 => to_signed(12496, LUT_AMPL_WIDTH),
		4082 => to_signed(12499, LUT_AMPL_WIDTH),
		4083 => to_signed(12502, LUT_AMPL_WIDTH),
		4084 => to_signed(12505, LUT_AMPL_WIDTH),
		4085 => to_signed(12507, LUT_AMPL_WIDTH),
		4086 => to_signed(12510, LUT_AMPL_WIDTH),
		4087 => to_signed(12513, LUT_AMPL_WIDTH),
		4088 => to_signed(12516, LUT_AMPL_WIDTH),
		4089 => to_signed(12519, LUT_AMPL_WIDTH),
		4090 => to_signed(12522, LUT_AMPL_WIDTH),
		4091 => to_signed(12525, LUT_AMPL_WIDTH),
		4092 => to_signed(12528, LUT_AMPL_WIDTH),
		4093 => to_signed(12531, LUT_AMPL_WIDTH),
		4094 => to_signed(12534, LUT_AMPL_WIDTH),
		4095 => to_signed(12536, LUT_AMPL_WIDTH),
		4096 => to_signed(12539, LUT_AMPL_WIDTH),
		4097 => to_signed(12542, LUT_AMPL_WIDTH),
		4098 => to_signed(12545, LUT_AMPL_WIDTH),
		4099 => to_signed(12548, LUT_AMPL_WIDTH),
		4100 => to_signed(12551, LUT_AMPL_WIDTH),
		4101 => to_signed(12554, LUT_AMPL_WIDTH),
		4102 => to_signed(12557, LUT_AMPL_WIDTH),
		4103 => to_signed(12560, LUT_AMPL_WIDTH),
		4104 => to_signed(12563, LUT_AMPL_WIDTH),
		4105 => to_signed(12566, LUT_AMPL_WIDTH),
		4106 => to_signed(12568, LUT_AMPL_WIDTH),
		4107 => to_signed(12571, LUT_AMPL_WIDTH),
		4108 => to_signed(12574, LUT_AMPL_WIDTH),
		4109 => to_signed(12577, LUT_AMPL_WIDTH),
		4110 => to_signed(12580, LUT_AMPL_WIDTH),
		4111 => to_signed(12583, LUT_AMPL_WIDTH),
		4112 => to_signed(12586, LUT_AMPL_WIDTH),
		4113 => to_signed(12589, LUT_AMPL_WIDTH),
		4114 => to_signed(12592, LUT_AMPL_WIDTH),
		4115 => to_signed(12595, LUT_AMPL_WIDTH),
		4116 => to_signed(12597, LUT_AMPL_WIDTH),
		4117 => to_signed(12600, LUT_AMPL_WIDTH),
		4118 => to_signed(12603, LUT_AMPL_WIDTH),
		4119 => to_signed(12606, LUT_AMPL_WIDTH),
		4120 => to_signed(12609, LUT_AMPL_WIDTH),
		4121 => to_signed(12612, LUT_AMPL_WIDTH),
		4122 => to_signed(12615, LUT_AMPL_WIDTH),
		4123 => to_signed(12618, LUT_AMPL_WIDTH),
		4124 => to_signed(12621, LUT_AMPL_WIDTH),
		4125 => to_signed(12624, LUT_AMPL_WIDTH),
		4126 => to_signed(12626, LUT_AMPL_WIDTH),
		4127 => to_signed(12629, LUT_AMPL_WIDTH),
		4128 => to_signed(12632, LUT_AMPL_WIDTH),
		4129 => to_signed(12635, LUT_AMPL_WIDTH),
		4130 => to_signed(12638, LUT_AMPL_WIDTH),
		4131 => to_signed(12641, LUT_AMPL_WIDTH),
		4132 => to_signed(12644, LUT_AMPL_WIDTH),
		4133 => to_signed(12647, LUT_AMPL_WIDTH),
		4134 => to_signed(12650, LUT_AMPL_WIDTH),
		4135 => to_signed(12652, LUT_AMPL_WIDTH),
		4136 => to_signed(12655, LUT_AMPL_WIDTH),
		4137 => to_signed(12658, LUT_AMPL_WIDTH),
		4138 => to_signed(12661, LUT_AMPL_WIDTH),
		4139 => to_signed(12664, LUT_AMPL_WIDTH),
		4140 => to_signed(12667, LUT_AMPL_WIDTH),
		4141 => to_signed(12670, LUT_AMPL_WIDTH),
		4142 => to_signed(12673, LUT_AMPL_WIDTH),
		4143 => to_signed(12676, LUT_AMPL_WIDTH),
		4144 => to_signed(12679, LUT_AMPL_WIDTH),
		4145 => to_signed(12681, LUT_AMPL_WIDTH),
		4146 => to_signed(12684, LUT_AMPL_WIDTH),
		4147 => to_signed(12687, LUT_AMPL_WIDTH),
		4148 => to_signed(12690, LUT_AMPL_WIDTH),
		4149 => to_signed(12693, LUT_AMPL_WIDTH),
		4150 => to_signed(12696, LUT_AMPL_WIDTH),
		4151 => to_signed(12699, LUT_AMPL_WIDTH),
		4152 => to_signed(12702, LUT_AMPL_WIDTH),
		4153 => to_signed(12705, LUT_AMPL_WIDTH),
		4154 => to_signed(12708, LUT_AMPL_WIDTH),
		4155 => to_signed(12710, LUT_AMPL_WIDTH),
		4156 => to_signed(12713, LUT_AMPL_WIDTH),
		4157 => to_signed(12716, LUT_AMPL_WIDTH),
		4158 => to_signed(12719, LUT_AMPL_WIDTH),
		4159 => to_signed(12722, LUT_AMPL_WIDTH),
		4160 => to_signed(12725, LUT_AMPL_WIDTH),
		4161 => to_signed(12728, LUT_AMPL_WIDTH),
		4162 => to_signed(12731, LUT_AMPL_WIDTH),
		4163 => to_signed(12734, LUT_AMPL_WIDTH),
		4164 => to_signed(12736, LUT_AMPL_WIDTH),
		4165 => to_signed(12739, LUT_AMPL_WIDTH),
		4166 => to_signed(12742, LUT_AMPL_WIDTH),
		4167 => to_signed(12745, LUT_AMPL_WIDTH),
		4168 => to_signed(12748, LUT_AMPL_WIDTH),
		4169 => to_signed(12751, LUT_AMPL_WIDTH),
		4170 => to_signed(12754, LUT_AMPL_WIDTH),
		4171 => to_signed(12757, LUT_AMPL_WIDTH),
		4172 => to_signed(12760, LUT_AMPL_WIDTH),
		4173 => to_signed(12763, LUT_AMPL_WIDTH),
		4174 => to_signed(12765, LUT_AMPL_WIDTH),
		4175 => to_signed(12768, LUT_AMPL_WIDTH),
		4176 => to_signed(12771, LUT_AMPL_WIDTH),
		4177 => to_signed(12774, LUT_AMPL_WIDTH),
		4178 => to_signed(12777, LUT_AMPL_WIDTH),
		4179 => to_signed(12780, LUT_AMPL_WIDTH),
		4180 => to_signed(12783, LUT_AMPL_WIDTH),
		4181 => to_signed(12786, LUT_AMPL_WIDTH),
		4182 => to_signed(12789, LUT_AMPL_WIDTH),
		4183 => to_signed(12791, LUT_AMPL_WIDTH),
		4184 => to_signed(12794, LUT_AMPL_WIDTH),
		4185 => to_signed(12797, LUT_AMPL_WIDTH),
		4186 => to_signed(12800, LUT_AMPL_WIDTH),
		4187 => to_signed(12803, LUT_AMPL_WIDTH),
		4188 => to_signed(12806, LUT_AMPL_WIDTH),
		4189 => to_signed(12809, LUT_AMPL_WIDTH),
		4190 => to_signed(12812, LUT_AMPL_WIDTH),
		4191 => to_signed(12815, LUT_AMPL_WIDTH),
		4192 => to_signed(12817, LUT_AMPL_WIDTH),
		4193 => to_signed(12820, LUT_AMPL_WIDTH),
		4194 => to_signed(12823, LUT_AMPL_WIDTH),
		4195 => to_signed(12826, LUT_AMPL_WIDTH),
		4196 => to_signed(12829, LUT_AMPL_WIDTH),
		4197 => to_signed(12832, LUT_AMPL_WIDTH),
		4198 => to_signed(12835, LUT_AMPL_WIDTH),
		4199 => to_signed(12838, LUT_AMPL_WIDTH),
		4200 => to_signed(12841, LUT_AMPL_WIDTH),
		4201 => to_signed(12843, LUT_AMPL_WIDTH),
		4202 => to_signed(12846, LUT_AMPL_WIDTH),
		4203 => to_signed(12849, LUT_AMPL_WIDTH),
		4204 => to_signed(12852, LUT_AMPL_WIDTH),
		4205 => to_signed(12855, LUT_AMPL_WIDTH),
		4206 => to_signed(12858, LUT_AMPL_WIDTH),
		4207 => to_signed(12861, LUT_AMPL_WIDTH),
		4208 => to_signed(12864, LUT_AMPL_WIDTH),
		4209 => to_signed(12867, LUT_AMPL_WIDTH),
		4210 => to_signed(12870, LUT_AMPL_WIDTH),
		4211 => to_signed(12872, LUT_AMPL_WIDTH),
		4212 => to_signed(12875, LUT_AMPL_WIDTH),
		4213 => to_signed(12878, LUT_AMPL_WIDTH),
		4214 => to_signed(12881, LUT_AMPL_WIDTH),
		4215 => to_signed(12884, LUT_AMPL_WIDTH),
		4216 => to_signed(12887, LUT_AMPL_WIDTH),
		4217 => to_signed(12890, LUT_AMPL_WIDTH),
		4218 => to_signed(12893, LUT_AMPL_WIDTH),
		4219 => to_signed(12895, LUT_AMPL_WIDTH),
		4220 => to_signed(12898, LUT_AMPL_WIDTH),
		4221 => to_signed(12901, LUT_AMPL_WIDTH),
		4222 => to_signed(12904, LUT_AMPL_WIDTH),
		4223 => to_signed(12907, LUT_AMPL_WIDTH),
		4224 => to_signed(12910, LUT_AMPL_WIDTH),
		4225 => to_signed(12913, LUT_AMPL_WIDTH),
		4226 => to_signed(12916, LUT_AMPL_WIDTH),
		4227 => to_signed(12919, LUT_AMPL_WIDTH),
		4228 => to_signed(12921, LUT_AMPL_WIDTH),
		4229 => to_signed(12924, LUT_AMPL_WIDTH),
		4230 => to_signed(12927, LUT_AMPL_WIDTH),
		4231 => to_signed(12930, LUT_AMPL_WIDTH),
		4232 => to_signed(12933, LUT_AMPL_WIDTH),
		4233 => to_signed(12936, LUT_AMPL_WIDTH),
		4234 => to_signed(12939, LUT_AMPL_WIDTH),
		4235 => to_signed(12942, LUT_AMPL_WIDTH),
		4236 => to_signed(12945, LUT_AMPL_WIDTH),
		4237 => to_signed(12947, LUT_AMPL_WIDTH),
		4238 => to_signed(12950, LUT_AMPL_WIDTH),
		4239 => to_signed(12953, LUT_AMPL_WIDTH),
		4240 => to_signed(12956, LUT_AMPL_WIDTH),
		4241 => to_signed(12959, LUT_AMPL_WIDTH),
		4242 => to_signed(12962, LUT_AMPL_WIDTH),
		4243 => to_signed(12965, LUT_AMPL_WIDTH),
		4244 => to_signed(12968, LUT_AMPL_WIDTH),
		4245 => to_signed(12971, LUT_AMPL_WIDTH),
		4246 => to_signed(12973, LUT_AMPL_WIDTH),
		4247 => to_signed(12976, LUT_AMPL_WIDTH),
		4248 => to_signed(12979, LUT_AMPL_WIDTH),
		4249 => to_signed(12982, LUT_AMPL_WIDTH),
		4250 => to_signed(12985, LUT_AMPL_WIDTH),
		4251 => to_signed(12988, LUT_AMPL_WIDTH),
		4252 => to_signed(12991, LUT_AMPL_WIDTH),
		4253 => to_signed(12994, LUT_AMPL_WIDTH),
		4254 => to_signed(12997, LUT_AMPL_WIDTH),
		4255 => to_signed(12999, LUT_AMPL_WIDTH),
		4256 => to_signed(13002, LUT_AMPL_WIDTH),
		4257 => to_signed(13005, LUT_AMPL_WIDTH),
		4258 => to_signed(13008, LUT_AMPL_WIDTH),
		4259 => to_signed(13011, LUT_AMPL_WIDTH),
		4260 => to_signed(13014, LUT_AMPL_WIDTH),
		4261 => to_signed(13017, LUT_AMPL_WIDTH),
		4262 => to_signed(13020, LUT_AMPL_WIDTH),
		4263 => to_signed(13022, LUT_AMPL_WIDTH),
		4264 => to_signed(13025, LUT_AMPL_WIDTH),
		4265 => to_signed(13028, LUT_AMPL_WIDTH),
		4266 => to_signed(13031, LUT_AMPL_WIDTH),
		4267 => to_signed(13034, LUT_AMPL_WIDTH),
		4268 => to_signed(13037, LUT_AMPL_WIDTH),
		4269 => to_signed(13040, LUT_AMPL_WIDTH),
		4270 => to_signed(13043, LUT_AMPL_WIDTH),
		4271 => to_signed(13046, LUT_AMPL_WIDTH),
		4272 => to_signed(13048, LUT_AMPL_WIDTH),
		4273 => to_signed(13051, LUT_AMPL_WIDTH),
		4274 => to_signed(13054, LUT_AMPL_WIDTH),
		4275 => to_signed(13057, LUT_AMPL_WIDTH),
		4276 => to_signed(13060, LUT_AMPL_WIDTH),
		4277 => to_signed(13063, LUT_AMPL_WIDTH),
		4278 => to_signed(13066, LUT_AMPL_WIDTH),
		4279 => to_signed(13069, LUT_AMPL_WIDTH),
		4280 => to_signed(13071, LUT_AMPL_WIDTH),
		4281 => to_signed(13074, LUT_AMPL_WIDTH),
		4282 => to_signed(13077, LUT_AMPL_WIDTH),
		4283 => to_signed(13080, LUT_AMPL_WIDTH),
		4284 => to_signed(13083, LUT_AMPL_WIDTH),
		4285 => to_signed(13086, LUT_AMPL_WIDTH),
		4286 => to_signed(13089, LUT_AMPL_WIDTH),
		4287 => to_signed(13092, LUT_AMPL_WIDTH),
		4288 => to_signed(13094, LUT_AMPL_WIDTH),
		4289 => to_signed(13097, LUT_AMPL_WIDTH),
		4290 => to_signed(13100, LUT_AMPL_WIDTH),
		4291 => to_signed(13103, LUT_AMPL_WIDTH),
		4292 => to_signed(13106, LUT_AMPL_WIDTH),
		4293 => to_signed(13109, LUT_AMPL_WIDTH),
		4294 => to_signed(13112, LUT_AMPL_WIDTH),
		4295 => to_signed(13115, LUT_AMPL_WIDTH),
		4296 => to_signed(13118, LUT_AMPL_WIDTH),
		4297 => to_signed(13120, LUT_AMPL_WIDTH),
		4298 => to_signed(13123, LUT_AMPL_WIDTH),
		4299 => to_signed(13126, LUT_AMPL_WIDTH),
		4300 => to_signed(13129, LUT_AMPL_WIDTH),
		4301 => to_signed(13132, LUT_AMPL_WIDTH),
		4302 => to_signed(13135, LUT_AMPL_WIDTH),
		4303 => to_signed(13138, LUT_AMPL_WIDTH),
		4304 => to_signed(13141, LUT_AMPL_WIDTH),
		4305 => to_signed(13143, LUT_AMPL_WIDTH),
		4306 => to_signed(13146, LUT_AMPL_WIDTH),
		4307 => to_signed(13149, LUT_AMPL_WIDTH),
		4308 => to_signed(13152, LUT_AMPL_WIDTH),
		4309 => to_signed(13155, LUT_AMPL_WIDTH),
		4310 => to_signed(13158, LUT_AMPL_WIDTH),
		4311 => to_signed(13161, LUT_AMPL_WIDTH),
		4312 => to_signed(13164, LUT_AMPL_WIDTH),
		4313 => to_signed(13166, LUT_AMPL_WIDTH),
		4314 => to_signed(13169, LUT_AMPL_WIDTH),
		4315 => to_signed(13172, LUT_AMPL_WIDTH),
		4316 => to_signed(13175, LUT_AMPL_WIDTH),
		4317 => to_signed(13178, LUT_AMPL_WIDTH),
		4318 => to_signed(13181, LUT_AMPL_WIDTH),
		4319 => to_signed(13184, LUT_AMPL_WIDTH),
		4320 => to_signed(13187, LUT_AMPL_WIDTH),
		4321 => to_signed(13189, LUT_AMPL_WIDTH),
		4322 => to_signed(13192, LUT_AMPL_WIDTH),
		4323 => to_signed(13195, LUT_AMPL_WIDTH),
		4324 => to_signed(13198, LUT_AMPL_WIDTH),
		4325 => to_signed(13201, LUT_AMPL_WIDTH),
		4326 => to_signed(13204, LUT_AMPL_WIDTH),
		4327 => to_signed(13207, LUT_AMPL_WIDTH),
		4328 => to_signed(13210, LUT_AMPL_WIDTH),
		4329 => to_signed(13212, LUT_AMPL_WIDTH),
		4330 => to_signed(13215, LUT_AMPL_WIDTH),
		4331 => to_signed(13218, LUT_AMPL_WIDTH),
		4332 => to_signed(13221, LUT_AMPL_WIDTH),
		4333 => to_signed(13224, LUT_AMPL_WIDTH),
		4334 => to_signed(13227, LUT_AMPL_WIDTH),
		4335 => to_signed(13230, LUT_AMPL_WIDTH),
		4336 => to_signed(13233, LUT_AMPL_WIDTH),
		4337 => to_signed(13235, LUT_AMPL_WIDTH),
		4338 => to_signed(13238, LUT_AMPL_WIDTH),
		4339 => to_signed(13241, LUT_AMPL_WIDTH),
		4340 => to_signed(13244, LUT_AMPL_WIDTH),
		4341 => to_signed(13247, LUT_AMPL_WIDTH),
		4342 => to_signed(13250, LUT_AMPL_WIDTH),
		4343 => to_signed(13253, LUT_AMPL_WIDTH),
		4344 => to_signed(13256, LUT_AMPL_WIDTH),
		4345 => to_signed(13258, LUT_AMPL_WIDTH),
		4346 => to_signed(13261, LUT_AMPL_WIDTH),
		4347 => to_signed(13264, LUT_AMPL_WIDTH),
		4348 => to_signed(13267, LUT_AMPL_WIDTH),
		4349 => to_signed(13270, LUT_AMPL_WIDTH),
		4350 => to_signed(13273, LUT_AMPL_WIDTH),
		4351 => to_signed(13276, LUT_AMPL_WIDTH),
		4352 => to_signed(13279, LUT_AMPL_WIDTH),
		4353 => to_signed(13281, LUT_AMPL_WIDTH),
		4354 => to_signed(13284, LUT_AMPL_WIDTH),
		4355 => to_signed(13287, LUT_AMPL_WIDTH),
		4356 => to_signed(13290, LUT_AMPL_WIDTH),
		4357 => to_signed(13293, LUT_AMPL_WIDTH),
		4358 => to_signed(13296, LUT_AMPL_WIDTH),
		4359 => to_signed(13299, LUT_AMPL_WIDTH),
		4360 => to_signed(13302, LUT_AMPL_WIDTH),
		4361 => to_signed(13304, LUT_AMPL_WIDTH),
		4362 => to_signed(13307, LUT_AMPL_WIDTH),
		4363 => to_signed(13310, LUT_AMPL_WIDTH),
		4364 => to_signed(13313, LUT_AMPL_WIDTH),
		4365 => to_signed(13316, LUT_AMPL_WIDTH),
		4366 => to_signed(13319, LUT_AMPL_WIDTH),
		4367 => to_signed(13322, LUT_AMPL_WIDTH),
		4368 => to_signed(13324, LUT_AMPL_WIDTH),
		4369 => to_signed(13327, LUT_AMPL_WIDTH),
		4370 => to_signed(13330, LUT_AMPL_WIDTH),
		4371 => to_signed(13333, LUT_AMPL_WIDTH),
		4372 => to_signed(13336, LUT_AMPL_WIDTH),
		4373 => to_signed(13339, LUT_AMPL_WIDTH),
		4374 => to_signed(13342, LUT_AMPL_WIDTH),
		4375 => to_signed(13345, LUT_AMPL_WIDTH),
		4376 => to_signed(13347, LUT_AMPL_WIDTH),
		4377 => to_signed(13350, LUT_AMPL_WIDTH),
		4378 => to_signed(13353, LUT_AMPL_WIDTH),
		4379 => to_signed(13356, LUT_AMPL_WIDTH),
		4380 => to_signed(13359, LUT_AMPL_WIDTH),
		4381 => to_signed(13362, LUT_AMPL_WIDTH),
		4382 => to_signed(13365, LUT_AMPL_WIDTH),
		4383 => to_signed(13368, LUT_AMPL_WIDTH),
		4384 => to_signed(13370, LUT_AMPL_WIDTH),
		4385 => to_signed(13373, LUT_AMPL_WIDTH),
		4386 => to_signed(13376, LUT_AMPL_WIDTH),
		4387 => to_signed(13379, LUT_AMPL_WIDTH),
		4388 => to_signed(13382, LUT_AMPL_WIDTH),
		4389 => to_signed(13385, LUT_AMPL_WIDTH),
		4390 => to_signed(13388, LUT_AMPL_WIDTH),
		4391 => to_signed(13390, LUT_AMPL_WIDTH),
		4392 => to_signed(13393, LUT_AMPL_WIDTH),
		4393 => to_signed(13396, LUT_AMPL_WIDTH),
		4394 => to_signed(13399, LUT_AMPL_WIDTH),
		4395 => to_signed(13402, LUT_AMPL_WIDTH),
		4396 => to_signed(13405, LUT_AMPL_WIDTH),
		4397 => to_signed(13408, LUT_AMPL_WIDTH),
		4398 => to_signed(13411, LUT_AMPL_WIDTH),
		4399 => to_signed(13413, LUT_AMPL_WIDTH),
		4400 => to_signed(13416, LUT_AMPL_WIDTH),
		4401 => to_signed(13419, LUT_AMPL_WIDTH),
		4402 => to_signed(13422, LUT_AMPL_WIDTH),
		4403 => to_signed(13425, LUT_AMPL_WIDTH),
		4404 => to_signed(13428, LUT_AMPL_WIDTH),
		4405 => to_signed(13431, LUT_AMPL_WIDTH),
		4406 => to_signed(13433, LUT_AMPL_WIDTH),
		4407 => to_signed(13436, LUT_AMPL_WIDTH),
		4408 => to_signed(13439, LUT_AMPL_WIDTH),
		4409 => to_signed(13442, LUT_AMPL_WIDTH),
		4410 => to_signed(13445, LUT_AMPL_WIDTH),
		4411 => to_signed(13448, LUT_AMPL_WIDTH),
		4412 => to_signed(13451, LUT_AMPL_WIDTH),
		4413 => to_signed(13454, LUT_AMPL_WIDTH),
		4414 => to_signed(13456, LUT_AMPL_WIDTH),
		4415 => to_signed(13459, LUT_AMPL_WIDTH),
		4416 => to_signed(13462, LUT_AMPL_WIDTH),
		4417 => to_signed(13465, LUT_AMPL_WIDTH),
		4418 => to_signed(13468, LUT_AMPL_WIDTH),
		4419 => to_signed(13471, LUT_AMPL_WIDTH),
		4420 => to_signed(13474, LUT_AMPL_WIDTH),
		4421 => to_signed(13476, LUT_AMPL_WIDTH),
		4422 => to_signed(13479, LUT_AMPL_WIDTH),
		4423 => to_signed(13482, LUT_AMPL_WIDTH),
		4424 => to_signed(13485, LUT_AMPL_WIDTH),
		4425 => to_signed(13488, LUT_AMPL_WIDTH),
		4426 => to_signed(13491, LUT_AMPL_WIDTH),
		4427 => to_signed(13494, LUT_AMPL_WIDTH),
		4428 => to_signed(13496, LUT_AMPL_WIDTH),
		4429 => to_signed(13499, LUT_AMPL_WIDTH),
		4430 => to_signed(13502, LUT_AMPL_WIDTH),
		4431 => to_signed(13505, LUT_AMPL_WIDTH),
		4432 => to_signed(13508, LUT_AMPL_WIDTH),
		4433 => to_signed(13511, LUT_AMPL_WIDTH),
		4434 => to_signed(13514, LUT_AMPL_WIDTH),
		4435 => to_signed(13516, LUT_AMPL_WIDTH),
		4436 => to_signed(13519, LUT_AMPL_WIDTH),
		4437 => to_signed(13522, LUT_AMPL_WIDTH),
		4438 => to_signed(13525, LUT_AMPL_WIDTH),
		4439 => to_signed(13528, LUT_AMPL_WIDTH),
		4440 => to_signed(13531, LUT_AMPL_WIDTH),
		4441 => to_signed(13534, LUT_AMPL_WIDTH),
		4442 => to_signed(13537, LUT_AMPL_WIDTH),
		4443 => to_signed(13539, LUT_AMPL_WIDTH),
		4444 => to_signed(13542, LUT_AMPL_WIDTH),
		4445 => to_signed(13545, LUT_AMPL_WIDTH),
		4446 => to_signed(13548, LUT_AMPL_WIDTH),
		4447 => to_signed(13551, LUT_AMPL_WIDTH),
		4448 => to_signed(13554, LUT_AMPL_WIDTH),
		4449 => to_signed(13557, LUT_AMPL_WIDTH),
		4450 => to_signed(13559, LUT_AMPL_WIDTH),
		4451 => to_signed(13562, LUT_AMPL_WIDTH),
		4452 => to_signed(13565, LUT_AMPL_WIDTH),
		4453 => to_signed(13568, LUT_AMPL_WIDTH),
		4454 => to_signed(13571, LUT_AMPL_WIDTH),
		4455 => to_signed(13574, LUT_AMPL_WIDTH),
		4456 => to_signed(13577, LUT_AMPL_WIDTH),
		4457 => to_signed(13579, LUT_AMPL_WIDTH),
		4458 => to_signed(13582, LUT_AMPL_WIDTH),
		4459 => to_signed(13585, LUT_AMPL_WIDTH),
		4460 => to_signed(13588, LUT_AMPL_WIDTH),
		4461 => to_signed(13591, LUT_AMPL_WIDTH),
		4462 => to_signed(13594, LUT_AMPL_WIDTH),
		4463 => to_signed(13597, LUT_AMPL_WIDTH),
		4464 => to_signed(13599, LUT_AMPL_WIDTH),
		4465 => to_signed(13602, LUT_AMPL_WIDTH),
		4466 => to_signed(13605, LUT_AMPL_WIDTH),
		4467 => to_signed(13608, LUT_AMPL_WIDTH),
		4468 => to_signed(13611, LUT_AMPL_WIDTH),
		4469 => to_signed(13614, LUT_AMPL_WIDTH),
		4470 => to_signed(13617, LUT_AMPL_WIDTH),
		4471 => to_signed(13619, LUT_AMPL_WIDTH),
		4472 => to_signed(13622, LUT_AMPL_WIDTH),
		4473 => to_signed(13625, LUT_AMPL_WIDTH),
		4474 => to_signed(13628, LUT_AMPL_WIDTH),
		4475 => to_signed(13631, LUT_AMPL_WIDTH),
		4476 => to_signed(13634, LUT_AMPL_WIDTH),
		4477 => to_signed(13637, LUT_AMPL_WIDTH),
		4478 => to_signed(13639, LUT_AMPL_WIDTH),
		4479 => to_signed(13642, LUT_AMPL_WIDTH),
		4480 => to_signed(13645, LUT_AMPL_WIDTH),
		4481 => to_signed(13648, LUT_AMPL_WIDTH),
		4482 => to_signed(13651, LUT_AMPL_WIDTH),
		4483 => to_signed(13654, LUT_AMPL_WIDTH),
		4484 => to_signed(13657, LUT_AMPL_WIDTH),
		4485 => to_signed(13659, LUT_AMPL_WIDTH),
		4486 => to_signed(13662, LUT_AMPL_WIDTH),
		4487 => to_signed(13665, LUT_AMPL_WIDTH),
		4488 => to_signed(13668, LUT_AMPL_WIDTH),
		4489 => to_signed(13671, LUT_AMPL_WIDTH),
		4490 => to_signed(13674, LUT_AMPL_WIDTH),
		4491 => to_signed(13677, LUT_AMPL_WIDTH),
		4492 => to_signed(13679, LUT_AMPL_WIDTH),
		4493 => to_signed(13682, LUT_AMPL_WIDTH),
		4494 => to_signed(13685, LUT_AMPL_WIDTH),
		4495 => to_signed(13688, LUT_AMPL_WIDTH),
		4496 => to_signed(13691, LUT_AMPL_WIDTH),
		4497 => to_signed(13694, LUT_AMPL_WIDTH),
		4498 => to_signed(13697, LUT_AMPL_WIDTH),
		4499 => to_signed(13699, LUT_AMPL_WIDTH),
		4500 => to_signed(13702, LUT_AMPL_WIDTH),
		4501 => to_signed(13705, LUT_AMPL_WIDTH),
		4502 => to_signed(13708, LUT_AMPL_WIDTH),
		4503 => to_signed(13711, LUT_AMPL_WIDTH),
		4504 => to_signed(13714, LUT_AMPL_WIDTH),
		4505 => to_signed(13717, LUT_AMPL_WIDTH),
		4506 => to_signed(13719, LUT_AMPL_WIDTH),
		4507 => to_signed(13722, LUT_AMPL_WIDTH),
		4508 => to_signed(13725, LUT_AMPL_WIDTH),
		4509 => to_signed(13728, LUT_AMPL_WIDTH),
		4510 => to_signed(13731, LUT_AMPL_WIDTH),
		4511 => to_signed(13734, LUT_AMPL_WIDTH),
		4512 => to_signed(13736, LUT_AMPL_WIDTH),
		4513 => to_signed(13739, LUT_AMPL_WIDTH),
		4514 => to_signed(13742, LUT_AMPL_WIDTH),
		4515 => to_signed(13745, LUT_AMPL_WIDTH),
		4516 => to_signed(13748, LUT_AMPL_WIDTH),
		4517 => to_signed(13751, LUT_AMPL_WIDTH),
		4518 => to_signed(13754, LUT_AMPL_WIDTH),
		4519 => to_signed(13756, LUT_AMPL_WIDTH),
		4520 => to_signed(13759, LUT_AMPL_WIDTH),
		4521 => to_signed(13762, LUT_AMPL_WIDTH),
		4522 => to_signed(13765, LUT_AMPL_WIDTH),
		4523 => to_signed(13768, LUT_AMPL_WIDTH),
		4524 => to_signed(13771, LUT_AMPL_WIDTH),
		4525 => to_signed(13774, LUT_AMPL_WIDTH),
		4526 => to_signed(13776, LUT_AMPL_WIDTH),
		4527 => to_signed(13779, LUT_AMPL_WIDTH),
		4528 => to_signed(13782, LUT_AMPL_WIDTH),
		4529 => to_signed(13785, LUT_AMPL_WIDTH),
		4530 => to_signed(13788, LUT_AMPL_WIDTH),
		4531 => to_signed(13791, LUT_AMPL_WIDTH),
		4532 => to_signed(13793, LUT_AMPL_WIDTH),
		4533 => to_signed(13796, LUT_AMPL_WIDTH),
		4534 => to_signed(13799, LUT_AMPL_WIDTH),
		4535 => to_signed(13802, LUT_AMPL_WIDTH),
		4536 => to_signed(13805, LUT_AMPL_WIDTH),
		4537 => to_signed(13808, LUT_AMPL_WIDTH),
		4538 => to_signed(13811, LUT_AMPL_WIDTH),
		4539 => to_signed(13813, LUT_AMPL_WIDTH),
		4540 => to_signed(13816, LUT_AMPL_WIDTH),
		4541 => to_signed(13819, LUT_AMPL_WIDTH),
		4542 => to_signed(13822, LUT_AMPL_WIDTH),
		4543 => to_signed(13825, LUT_AMPL_WIDTH),
		4544 => to_signed(13828, LUT_AMPL_WIDTH),
		4545 => to_signed(13831, LUT_AMPL_WIDTH),
		4546 => to_signed(13833, LUT_AMPL_WIDTH),
		4547 => to_signed(13836, LUT_AMPL_WIDTH),
		4548 => to_signed(13839, LUT_AMPL_WIDTH),
		4549 => to_signed(13842, LUT_AMPL_WIDTH),
		4550 => to_signed(13845, LUT_AMPL_WIDTH),
		4551 => to_signed(13848, LUT_AMPL_WIDTH),
		4552 => to_signed(13850, LUT_AMPL_WIDTH),
		4553 => to_signed(13853, LUT_AMPL_WIDTH),
		4554 => to_signed(13856, LUT_AMPL_WIDTH),
		4555 => to_signed(13859, LUT_AMPL_WIDTH),
		4556 => to_signed(13862, LUT_AMPL_WIDTH),
		4557 => to_signed(13865, LUT_AMPL_WIDTH),
		4558 => to_signed(13868, LUT_AMPL_WIDTH),
		4559 => to_signed(13870, LUT_AMPL_WIDTH),
		4560 => to_signed(13873, LUT_AMPL_WIDTH),
		4561 => to_signed(13876, LUT_AMPL_WIDTH),
		4562 => to_signed(13879, LUT_AMPL_WIDTH),
		4563 => to_signed(13882, LUT_AMPL_WIDTH),
		4564 => to_signed(13885, LUT_AMPL_WIDTH),
		4565 => to_signed(13887, LUT_AMPL_WIDTH),
		4566 => to_signed(13890, LUT_AMPL_WIDTH),
		4567 => to_signed(13893, LUT_AMPL_WIDTH),
		4568 => to_signed(13896, LUT_AMPL_WIDTH),
		4569 => to_signed(13899, LUT_AMPL_WIDTH),
		4570 => to_signed(13902, LUT_AMPL_WIDTH),
		4571 => to_signed(13905, LUT_AMPL_WIDTH),
		4572 => to_signed(13907, LUT_AMPL_WIDTH),
		4573 => to_signed(13910, LUT_AMPL_WIDTH),
		4574 => to_signed(13913, LUT_AMPL_WIDTH),
		4575 => to_signed(13916, LUT_AMPL_WIDTH),
		4576 => to_signed(13919, LUT_AMPL_WIDTH),
		4577 => to_signed(13922, LUT_AMPL_WIDTH),
		4578 => to_signed(13924, LUT_AMPL_WIDTH),
		4579 => to_signed(13927, LUT_AMPL_WIDTH),
		4580 => to_signed(13930, LUT_AMPL_WIDTH),
		4581 => to_signed(13933, LUT_AMPL_WIDTH),
		4582 => to_signed(13936, LUT_AMPL_WIDTH),
		4583 => to_signed(13939, LUT_AMPL_WIDTH),
		4584 => to_signed(13942, LUT_AMPL_WIDTH),
		4585 => to_signed(13944, LUT_AMPL_WIDTH),
		4586 => to_signed(13947, LUT_AMPL_WIDTH),
		4587 => to_signed(13950, LUT_AMPL_WIDTH),
		4588 => to_signed(13953, LUT_AMPL_WIDTH),
		4589 => to_signed(13956, LUT_AMPL_WIDTH),
		4590 => to_signed(13959, LUT_AMPL_WIDTH),
		4591 => to_signed(13961, LUT_AMPL_WIDTH),
		4592 => to_signed(13964, LUT_AMPL_WIDTH),
		4593 => to_signed(13967, LUT_AMPL_WIDTH),
		4594 => to_signed(13970, LUT_AMPL_WIDTH),
		4595 => to_signed(13973, LUT_AMPL_WIDTH),
		4596 => to_signed(13976, LUT_AMPL_WIDTH),
		4597 => to_signed(13978, LUT_AMPL_WIDTH),
		4598 => to_signed(13981, LUT_AMPL_WIDTH),
		4599 => to_signed(13984, LUT_AMPL_WIDTH),
		4600 => to_signed(13987, LUT_AMPL_WIDTH),
		4601 => to_signed(13990, LUT_AMPL_WIDTH),
		4602 => to_signed(13993, LUT_AMPL_WIDTH),
		4603 => to_signed(13995, LUT_AMPL_WIDTH),
		4604 => to_signed(13998, LUT_AMPL_WIDTH),
		4605 => to_signed(14001, LUT_AMPL_WIDTH),
		4606 => to_signed(14004, LUT_AMPL_WIDTH),
		4607 => to_signed(14007, LUT_AMPL_WIDTH),
		4608 => to_signed(14010, LUT_AMPL_WIDTH),
		4609 => to_signed(14013, LUT_AMPL_WIDTH),
		4610 => to_signed(14015, LUT_AMPL_WIDTH),
		4611 => to_signed(14018, LUT_AMPL_WIDTH),
		4612 => to_signed(14021, LUT_AMPL_WIDTH),
		4613 => to_signed(14024, LUT_AMPL_WIDTH),
		4614 => to_signed(14027, LUT_AMPL_WIDTH),
		4615 => to_signed(14030, LUT_AMPL_WIDTH),
		4616 => to_signed(14032, LUT_AMPL_WIDTH),
		4617 => to_signed(14035, LUT_AMPL_WIDTH),
		4618 => to_signed(14038, LUT_AMPL_WIDTH),
		4619 => to_signed(14041, LUT_AMPL_WIDTH),
		4620 => to_signed(14044, LUT_AMPL_WIDTH),
		4621 => to_signed(14047, LUT_AMPL_WIDTH),
		4622 => to_signed(14049, LUT_AMPL_WIDTH),
		4623 => to_signed(14052, LUT_AMPL_WIDTH),
		4624 => to_signed(14055, LUT_AMPL_WIDTH),
		4625 => to_signed(14058, LUT_AMPL_WIDTH),
		4626 => to_signed(14061, LUT_AMPL_WIDTH),
		4627 => to_signed(14064, LUT_AMPL_WIDTH),
		4628 => to_signed(14066, LUT_AMPL_WIDTH),
		4629 => to_signed(14069, LUT_AMPL_WIDTH),
		4630 => to_signed(14072, LUT_AMPL_WIDTH),
		4631 => to_signed(14075, LUT_AMPL_WIDTH),
		4632 => to_signed(14078, LUT_AMPL_WIDTH),
		4633 => to_signed(14081, LUT_AMPL_WIDTH),
		4634 => to_signed(14083, LUT_AMPL_WIDTH),
		4635 => to_signed(14086, LUT_AMPL_WIDTH),
		4636 => to_signed(14089, LUT_AMPL_WIDTH),
		4637 => to_signed(14092, LUT_AMPL_WIDTH),
		4638 => to_signed(14095, LUT_AMPL_WIDTH),
		4639 => to_signed(14098, LUT_AMPL_WIDTH),
		4640 => to_signed(14101, LUT_AMPL_WIDTH),
		4641 => to_signed(14103, LUT_AMPL_WIDTH),
		4642 => to_signed(14106, LUT_AMPL_WIDTH),
		4643 => to_signed(14109, LUT_AMPL_WIDTH),
		4644 => to_signed(14112, LUT_AMPL_WIDTH),
		4645 => to_signed(14115, LUT_AMPL_WIDTH),
		4646 => to_signed(14118, LUT_AMPL_WIDTH),
		4647 => to_signed(14120, LUT_AMPL_WIDTH),
		4648 => to_signed(14123, LUT_AMPL_WIDTH),
		4649 => to_signed(14126, LUT_AMPL_WIDTH),
		4650 => to_signed(14129, LUT_AMPL_WIDTH),
		4651 => to_signed(14132, LUT_AMPL_WIDTH),
		4652 => to_signed(14135, LUT_AMPL_WIDTH),
		4653 => to_signed(14137, LUT_AMPL_WIDTH),
		4654 => to_signed(14140, LUT_AMPL_WIDTH),
		4655 => to_signed(14143, LUT_AMPL_WIDTH),
		4656 => to_signed(14146, LUT_AMPL_WIDTH),
		4657 => to_signed(14149, LUT_AMPL_WIDTH),
		4658 => to_signed(14152, LUT_AMPL_WIDTH),
		4659 => to_signed(14154, LUT_AMPL_WIDTH),
		4660 => to_signed(14157, LUT_AMPL_WIDTH),
		4661 => to_signed(14160, LUT_AMPL_WIDTH),
		4662 => to_signed(14163, LUT_AMPL_WIDTH),
		4663 => to_signed(14166, LUT_AMPL_WIDTH),
		4664 => to_signed(14169, LUT_AMPL_WIDTH),
		4665 => to_signed(14171, LUT_AMPL_WIDTH),
		4666 => to_signed(14174, LUT_AMPL_WIDTH),
		4667 => to_signed(14177, LUT_AMPL_WIDTH),
		4668 => to_signed(14180, LUT_AMPL_WIDTH),
		4669 => to_signed(14183, LUT_AMPL_WIDTH),
		4670 => to_signed(14186, LUT_AMPL_WIDTH),
		4671 => to_signed(14188, LUT_AMPL_WIDTH),
		4672 => to_signed(14191, LUT_AMPL_WIDTH),
		4673 => to_signed(14194, LUT_AMPL_WIDTH),
		4674 => to_signed(14197, LUT_AMPL_WIDTH),
		4675 => to_signed(14200, LUT_AMPL_WIDTH),
		4676 => to_signed(14203, LUT_AMPL_WIDTH),
		4677 => to_signed(14205, LUT_AMPL_WIDTH),
		4678 => to_signed(14208, LUT_AMPL_WIDTH),
		4679 => to_signed(14211, LUT_AMPL_WIDTH),
		4680 => to_signed(14214, LUT_AMPL_WIDTH),
		4681 => to_signed(14217, LUT_AMPL_WIDTH),
		4682 => to_signed(14219, LUT_AMPL_WIDTH),
		4683 => to_signed(14222, LUT_AMPL_WIDTH),
		4684 => to_signed(14225, LUT_AMPL_WIDTH),
		4685 => to_signed(14228, LUT_AMPL_WIDTH),
		4686 => to_signed(14231, LUT_AMPL_WIDTH),
		4687 => to_signed(14234, LUT_AMPL_WIDTH),
		4688 => to_signed(14236, LUT_AMPL_WIDTH),
		4689 => to_signed(14239, LUT_AMPL_WIDTH),
		4690 => to_signed(14242, LUT_AMPL_WIDTH),
		4691 => to_signed(14245, LUT_AMPL_WIDTH),
		4692 => to_signed(14248, LUT_AMPL_WIDTH),
		4693 => to_signed(14251, LUT_AMPL_WIDTH),
		4694 => to_signed(14253, LUT_AMPL_WIDTH),
		4695 => to_signed(14256, LUT_AMPL_WIDTH),
		4696 => to_signed(14259, LUT_AMPL_WIDTH),
		4697 => to_signed(14262, LUT_AMPL_WIDTH),
		4698 => to_signed(14265, LUT_AMPL_WIDTH),
		4699 => to_signed(14268, LUT_AMPL_WIDTH),
		4700 => to_signed(14270, LUT_AMPL_WIDTH),
		4701 => to_signed(14273, LUT_AMPL_WIDTH),
		4702 => to_signed(14276, LUT_AMPL_WIDTH),
		4703 => to_signed(14279, LUT_AMPL_WIDTH),
		4704 => to_signed(14282, LUT_AMPL_WIDTH),
		4705 => to_signed(14285, LUT_AMPL_WIDTH),
		4706 => to_signed(14287, LUT_AMPL_WIDTH),
		4707 => to_signed(14290, LUT_AMPL_WIDTH),
		4708 => to_signed(14293, LUT_AMPL_WIDTH),
		4709 => to_signed(14296, LUT_AMPL_WIDTH),
		4710 => to_signed(14299, LUT_AMPL_WIDTH),
		4711 => to_signed(14302, LUT_AMPL_WIDTH),
		4712 => to_signed(14304, LUT_AMPL_WIDTH),
		4713 => to_signed(14307, LUT_AMPL_WIDTH),
		4714 => to_signed(14310, LUT_AMPL_WIDTH),
		4715 => to_signed(14313, LUT_AMPL_WIDTH),
		4716 => to_signed(14316, LUT_AMPL_WIDTH),
		4717 => to_signed(14318, LUT_AMPL_WIDTH),
		4718 => to_signed(14321, LUT_AMPL_WIDTH),
		4719 => to_signed(14324, LUT_AMPL_WIDTH),
		4720 => to_signed(14327, LUT_AMPL_WIDTH),
		4721 => to_signed(14330, LUT_AMPL_WIDTH),
		4722 => to_signed(14333, LUT_AMPL_WIDTH),
		4723 => to_signed(14335, LUT_AMPL_WIDTH),
		4724 => to_signed(14338, LUT_AMPL_WIDTH),
		4725 => to_signed(14341, LUT_AMPL_WIDTH),
		4726 => to_signed(14344, LUT_AMPL_WIDTH),
		4727 => to_signed(14347, LUT_AMPL_WIDTH),
		4728 => to_signed(14350, LUT_AMPL_WIDTH),
		4729 => to_signed(14352, LUT_AMPL_WIDTH),
		4730 => to_signed(14355, LUT_AMPL_WIDTH),
		4731 => to_signed(14358, LUT_AMPL_WIDTH),
		4732 => to_signed(14361, LUT_AMPL_WIDTH),
		4733 => to_signed(14364, LUT_AMPL_WIDTH),
		4734 => to_signed(14366, LUT_AMPL_WIDTH),
		4735 => to_signed(14369, LUT_AMPL_WIDTH),
		4736 => to_signed(14372, LUT_AMPL_WIDTH),
		4737 => to_signed(14375, LUT_AMPL_WIDTH),
		4738 => to_signed(14378, LUT_AMPL_WIDTH),
		4739 => to_signed(14381, LUT_AMPL_WIDTH),
		4740 => to_signed(14383, LUT_AMPL_WIDTH),
		4741 => to_signed(14386, LUT_AMPL_WIDTH),
		4742 => to_signed(14389, LUT_AMPL_WIDTH),
		4743 => to_signed(14392, LUT_AMPL_WIDTH),
		4744 => to_signed(14395, LUT_AMPL_WIDTH),
		4745 => to_signed(14398, LUT_AMPL_WIDTH),
		4746 => to_signed(14400, LUT_AMPL_WIDTH),
		4747 => to_signed(14403, LUT_AMPL_WIDTH),
		4748 => to_signed(14406, LUT_AMPL_WIDTH),
		4749 => to_signed(14409, LUT_AMPL_WIDTH),
		4750 => to_signed(14412, LUT_AMPL_WIDTH),
		4751 => to_signed(14414, LUT_AMPL_WIDTH),
		4752 => to_signed(14417, LUT_AMPL_WIDTH),
		4753 => to_signed(14420, LUT_AMPL_WIDTH),
		4754 => to_signed(14423, LUT_AMPL_WIDTH),
		4755 => to_signed(14426, LUT_AMPL_WIDTH),
		4756 => to_signed(14429, LUT_AMPL_WIDTH),
		4757 => to_signed(14431, LUT_AMPL_WIDTH),
		4758 => to_signed(14434, LUT_AMPL_WIDTH),
		4759 => to_signed(14437, LUT_AMPL_WIDTH),
		4760 => to_signed(14440, LUT_AMPL_WIDTH),
		4761 => to_signed(14443, LUT_AMPL_WIDTH),
		4762 => to_signed(14445, LUT_AMPL_WIDTH),
		4763 => to_signed(14448, LUT_AMPL_WIDTH),
		4764 => to_signed(14451, LUT_AMPL_WIDTH),
		4765 => to_signed(14454, LUT_AMPL_WIDTH),
		4766 => to_signed(14457, LUT_AMPL_WIDTH),
		4767 => to_signed(14460, LUT_AMPL_WIDTH),
		4768 => to_signed(14462, LUT_AMPL_WIDTH),
		4769 => to_signed(14465, LUT_AMPL_WIDTH),
		4770 => to_signed(14468, LUT_AMPL_WIDTH),
		4771 => to_signed(14471, LUT_AMPL_WIDTH),
		4772 => to_signed(14474, LUT_AMPL_WIDTH),
		4773 => to_signed(14477, LUT_AMPL_WIDTH),
		4774 => to_signed(14479, LUT_AMPL_WIDTH),
		4775 => to_signed(14482, LUT_AMPL_WIDTH),
		4776 => to_signed(14485, LUT_AMPL_WIDTH),
		4777 => to_signed(14488, LUT_AMPL_WIDTH),
		4778 => to_signed(14491, LUT_AMPL_WIDTH),
		4779 => to_signed(14493, LUT_AMPL_WIDTH),
		4780 => to_signed(14496, LUT_AMPL_WIDTH),
		4781 => to_signed(14499, LUT_AMPL_WIDTH),
		4782 => to_signed(14502, LUT_AMPL_WIDTH),
		4783 => to_signed(14505, LUT_AMPL_WIDTH),
		4784 => to_signed(14507, LUT_AMPL_WIDTH),
		4785 => to_signed(14510, LUT_AMPL_WIDTH),
		4786 => to_signed(14513, LUT_AMPL_WIDTH),
		4787 => to_signed(14516, LUT_AMPL_WIDTH),
		4788 => to_signed(14519, LUT_AMPL_WIDTH),
		4789 => to_signed(14522, LUT_AMPL_WIDTH),
		4790 => to_signed(14524, LUT_AMPL_WIDTH),
		4791 => to_signed(14527, LUT_AMPL_WIDTH),
		4792 => to_signed(14530, LUT_AMPL_WIDTH),
		4793 => to_signed(14533, LUT_AMPL_WIDTH),
		4794 => to_signed(14536, LUT_AMPL_WIDTH),
		4795 => to_signed(14538, LUT_AMPL_WIDTH),
		4796 => to_signed(14541, LUT_AMPL_WIDTH),
		4797 => to_signed(14544, LUT_AMPL_WIDTH),
		4798 => to_signed(14547, LUT_AMPL_WIDTH),
		4799 => to_signed(14550, LUT_AMPL_WIDTH),
		4800 => to_signed(14553, LUT_AMPL_WIDTH),
		4801 => to_signed(14555, LUT_AMPL_WIDTH),
		4802 => to_signed(14558, LUT_AMPL_WIDTH),
		4803 => to_signed(14561, LUT_AMPL_WIDTH),
		4804 => to_signed(14564, LUT_AMPL_WIDTH),
		4805 => to_signed(14567, LUT_AMPL_WIDTH),
		4806 => to_signed(14569, LUT_AMPL_WIDTH),
		4807 => to_signed(14572, LUT_AMPL_WIDTH),
		4808 => to_signed(14575, LUT_AMPL_WIDTH),
		4809 => to_signed(14578, LUT_AMPL_WIDTH),
		4810 => to_signed(14581, LUT_AMPL_WIDTH),
		4811 => to_signed(14584, LUT_AMPL_WIDTH),
		4812 => to_signed(14586, LUT_AMPL_WIDTH),
		4813 => to_signed(14589, LUT_AMPL_WIDTH),
		4814 => to_signed(14592, LUT_AMPL_WIDTH),
		4815 => to_signed(14595, LUT_AMPL_WIDTH),
		4816 => to_signed(14598, LUT_AMPL_WIDTH),
		4817 => to_signed(14600, LUT_AMPL_WIDTH),
		4818 => to_signed(14603, LUT_AMPL_WIDTH),
		4819 => to_signed(14606, LUT_AMPL_WIDTH),
		4820 => to_signed(14609, LUT_AMPL_WIDTH),
		4821 => to_signed(14612, LUT_AMPL_WIDTH),
		4822 => to_signed(14614, LUT_AMPL_WIDTH),
		4823 => to_signed(14617, LUT_AMPL_WIDTH),
		4824 => to_signed(14620, LUT_AMPL_WIDTH),
		4825 => to_signed(14623, LUT_AMPL_WIDTH),
		4826 => to_signed(14626, LUT_AMPL_WIDTH),
		4827 => to_signed(14628, LUT_AMPL_WIDTH),
		4828 => to_signed(14631, LUT_AMPL_WIDTH),
		4829 => to_signed(14634, LUT_AMPL_WIDTH),
		4830 => to_signed(14637, LUT_AMPL_WIDTH),
		4831 => to_signed(14640, LUT_AMPL_WIDTH),
		4832 => to_signed(14643, LUT_AMPL_WIDTH),
		4833 => to_signed(14645, LUT_AMPL_WIDTH),
		4834 => to_signed(14648, LUT_AMPL_WIDTH),
		4835 => to_signed(14651, LUT_AMPL_WIDTH),
		4836 => to_signed(14654, LUT_AMPL_WIDTH),
		4837 => to_signed(14657, LUT_AMPL_WIDTH),
		4838 => to_signed(14659, LUT_AMPL_WIDTH),
		4839 => to_signed(14662, LUT_AMPL_WIDTH),
		4840 => to_signed(14665, LUT_AMPL_WIDTH),
		4841 => to_signed(14668, LUT_AMPL_WIDTH),
		4842 => to_signed(14671, LUT_AMPL_WIDTH),
		4843 => to_signed(14673, LUT_AMPL_WIDTH),
		4844 => to_signed(14676, LUT_AMPL_WIDTH),
		4845 => to_signed(14679, LUT_AMPL_WIDTH),
		4846 => to_signed(14682, LUT_AMPL_WIDTH),
		4847 => to_signed(14685, LUT_AMPL_WIDTH),
		4848 => to_signed(14688, LUT_AMPL_WIDTH),
		4849 => to_signed(14690, LUT_AMPL_WIDTH),
		4850 => to_signed(14693, LUT_AMPL_WIDTH),
		4851 => to_signed(14696, LUT_AMPL_WIDTH),
		4852 => to_signed(14699, LUT_AMPL_WIDTH),
		4853 => to_signed(14702, LUT_AMPL_WIDTH),
		4854 => to_signed(14704, LUT_AMPL_WIDTH),
		4855 => to_signed(14707, LUT_AMPL_WIDTH),
		4856 => to_signed(14710, LUT_AMPL_WIDTH),
		4857 => to_signed(14713, LUT_AMPL_WIDTH),
		4858 => to_signed(14716, LUT_AMPL_WIDTH),
		4859 => to_signed(14718, LUT_AMPL_WIDTH),
		4860 => to_signed(14721, LUT_AMPL_WIDTH),
		4861 => to_signed(14724, LUT_AMPL_WIDTH),
		4862 => to_signed(14727, LUT_AMPL_WIDTH),
		4863 => to_signed(14730, LUT_AMPL_WIDTH),
		4864 => to_signed(14732, LUT_AMPL_WIDTH),
		4865 => to_signed(14735, LUT_AMPL_WIDTH),
		4866 => to_signed(14738, LUT_AMPL_WIDTH),
		4867 => to_signed(14741, LUT_AMPL_WIDTH),
		4868 => to_signed(14744, LUT_AMPL_WIDTH),
		4869 => to_signed(14746, LUT_AMPL_WIDTH),
		4870 => to_signed(14749, LUT_AMPL_WIDTH),
		4871 => to_signed(14752, LUT_AMPL_WIDTH),
		4872 => to_signed(14755, LUT_AMPL_WIDTH),
		4873 => to_signed(14758, LUT_AMPL_WIDTH),
		4874 => to_signed(14760, LUT_AMPL_WIDTH),
		4875 => to_signed(14763, LUT_AMPL_WIDTH),
		4876 => to_signed(14766, LUT_AMPL_WIDTH),
		4877 => to_signed(14769, LUT_AMPL_WIDTH),
		4878 => to_signed(14772, LUT_AMPL_WIDTH),
		4879 => to_signed(14774, LUT_AMPL_WIDTH),
		4880 => to_signed(14777, LUT_AMPL_WIDTH),
		4881 => to_signed(14780, LUT_AMPL_WIDTH),
		4882 => to_signed(14783, LUT_AMPL_WIDTH),
		4883 => to_signed(14786, LUT_AMPL_WIDTH),
		4884 => to_signed(14789, LUT_AMPL_WIDTH),
		4885 => to_signed(14791, LUT_AMPL_WIDTH),
		4886 => to_signed(14794, LUT_AMPL_WIDTH),
		4887 => to_signed(14797, LUT_AMPL_WIDTH),
		4888 => to_signed(14800, LUT_AMPL_WIDTH),
		4889 => to_signed(14803, LUT_AMPL_WIDTH),
		4890 => to_signed(14805, LUT_AMPL_WIDTH),
		4891 => to_signed(14808, LUT_AMPL_WIDTH),
		4892 => to_signed(14811, LUT_AMPL_WIDTH),
		4893 => to_signed(14814, LUT_AMPL_WIDTH),
		4894 => to_signed(14817, LUT_AMPL_WIDTH),
		4895 => to_signed(14819, LUT_AMPL_WIDTH),
		4896 => to_signed(14822, LUT_AMPL_WIDTH),
		4897 => to_signed(14825, LUT_AMPL_WIDTH),
		4898 => to_signed(14828, LUT_AMPL_WIDTH),
		4899 => to_signed(14831, LUT_AMPL_WIDTH),
		4900 => to_signed(14833, LUT_AMPL_WIDTH),
		4901 => to_signed(14836, LUT_AMPL_WIDTH),
		4902 => to_signed(14839, LUT_AMPL_WIDTH),
		4903 => to_signed(14842, LUT_AMPL_WIDTH),
		4904 => to_signed(14845, LUT_AMPL_WIDTH),
		4905 => to_signed(14847, LUT_AMPL_WIDTH),
		4906 => to_signed(14850, LUT_AMPL_WIDTH),
		4907 => to_signed(14853, LUT_AMPL_WIDTH),
		4908 => to_signed(14856, LUT_AMPL_WIDTH),
		4909 => to_signed(14859, LUT_AMPL_WIDTH),
		4910 => to_signed(14861, LUT_AMPL_WIDTH),
		4911 => to_signed(14864, LUT_AMPL_WIDTH),
		4912 => to_signed(14867, LUT_AMPL_WIDTH),
		4913 => to_signed(14870, LUT_AMPL_WIDTH),
		4914 => to_signed(14873, LUT_AMPL_WIDTH),
		4915 => to_signed(14875, LUT_AMPL_WIDTH),
		4916 => to_signed(14878, LUT_AMPL_WIDTH),
		4917 => to_signed(14881, LUT_AMPL_WIDTH),
		4918 => to_signed(14884, LUT_AMPL_WIDTH),
		4919 => to_signed(14887, LUT_AMPL_WIDTH),
		4920 => to_signed(14889, LUT_AMPL_WIDTH),
		4921 => to_signed(14892, LUT_AMPL_WIDTH),
		4922 => to_signed(14895, LUT_AMPL_WIDTH),
		4923 => to_signed(14898, LUT_AMPL_WIDTH),
		4924 => to_signed(14901, LUT_AMPL_WIDTH),
		4925 => to_signed(14903, LUT_AMPL_WIDTH),
		4926 => to_signed(14906, LUT_AMPL_WIDTH),
		4927 => to_signed(14909, LUT_AMPL_WIDTH),
		4928 => to_signed(14912, LUT_AMPL_WIDTH),
		4929 => to_signed(14915, LUT_AMPL_WIDTH),
		4930 => to_signed(14917, LUT_AMPL_WIDTH),
		4931 => to_signed(14920, LUT_AMPL_WIDTH),
		4932 => to_signed(14923, LUT_AMPL_WIDTH),
		4933 => to_signed(14926, LUT_AMPL_WIDTH),
		4934 => to_signed(14929, LUT_AMPL_WIDTH),
		4935 => to_signed(14931, LUT_AMPL_WIDTH),
		4936 => to_signed(14934, LUT_AMPL_WIDTH),
		4937 => to_signed(14937, LUT_AMPL_WIDTH),
		4938 => to_signed(14940, LUT_AMPL_WIDTH),
		4939 => to_signed(14942, LUT_AMPL_WIDTH),
		4940 => to_signed(14945, LUT_AMPL_WIDTH),
		4941 => to_signed(14948, LUT_AMPL_WIDTH),
		4942 => to_signed(14951, LUT_AMPL_WIDTH),
		4943 => to_signed(14954, LUT_AMPL_WIDTH),
		4944 => to_signed(14956, LUT_AMPL_WIDTH),
		4945 => to_signed(14959, LUT_AMPL_WIDTH),
		4946 => to_signed(14962, LUT_AMPL_WIDTH),
		4947 => to_signed(14965, LUT_AMPL_WIDTH),
		4948 => to_signed(14968, LUT_AMPL_WIDTH),
		4949 => to_signed(14970, LUT_AMPL_WIDTH),
		4950 => to_signed(14973, LUT_AMPL_WIDTH),
		4951 => to_signed(14976, LUT_AMPL_WIDTH),
		4952 => to_signed(14979, LUT_AMPL_WIDTH),
		4953 => to_signed(14982, LUT_AMPL_WIDTH),
		4954 => to_signed(14984, LUT_AMPL_WIDTH),
		4955 => to_signed(14987, LUT_AMPL_WIDTH),
		4956 => to_signed(14990, LUT_AMPL_WIDTH),
		4957 => to_signed(14993, LUT_AMPL_WIDTH),
		4958 => to_signed(14996, LUT_AMPL_WIDTH),
		4959 => to_signed(14998, LUT_AMPL_WIDTH),
		4960 => to_signed(15001, LUT_AMPL_WIDTH),
		4961 => to_signed(15004, LUT_AMPL_WIDTH),
		4962 => to_signed(15007, LUT_AMPL_WIDTH),
		4963 => to_signed(15010, LUT_AMPL_WIDTH),
		4964 => to_signed(15012, LUT_AMPL_WIDTH),
		4965 => to_signed(15015, LUT_AMPL_WIDTH),
		4966 => to_signed(15018, LUT_AMPL_WIDTH),
		4967 => to_signed(15021, LUT_AMPL_WIDTH),
		4968 => to_signed(15024, LUT_AMPL_WIDTH),
		4969 => to_signed(15026, LUT_AMPL_WIDTH),
		4970 => to_signed(15029, LUT_AMPL_WIDTH),
		4971 => to_signed(15032, LUT_AMPL_WIDTH),
		4972 => to_signed(15035, LUT_AMPL_WIDTH),
		4973 => to_signed(15037, LUT_AMPL_WIDTH),
		4974 => to_signed(15040, LUT_AMPL_WIDTH),
		4975 => to_signed(15043, LUT_AMPL_WIDTH),
		4976 => to_signed(15046, LUT_AMPL_WIDTH),
		4977 => to_signed(15049, LUT_AMPL_WIDTH),
		4978 => to_signed(15051, LUT_AMPL_WIDTH),
		4979 => to_signed(15054, LUT_AMPL_WIDTH),
		4980 => to_signed(15057, LUT_AMPL_WIDTH),
		4981 => to_signed(15060, LUT_AMPL_WIDTH),
		4982 => to_signed(15063, LUT_AMPL_WIDTH),
		4983 => to_signed(15065, LUT_AMPL_WIDTH),
		4984 => to_signed(15068, LUT_AMPL_WIDTH),
		4985 => to_signed(15071, LUT_AMPL_WIDTH),
		4986 => to_signed(15074, LUT_AMPL_WIDTH),
		4987 => to_signed(15077, LUT_AMPL_WIDTH),
		4988 => to_signed(15079, LUT_AMPL_WIDTH),
		4989 => to_signed(15082, LUT_AMPL_WIDTH),
		4990 => to_signed(15085, LUT_AMPL_WIDTH),
		4991 => to_signed(15088, LUT_AMPL_WIDTH),
		4992 => to_signed(15090, LUT_AMPL_WIDTH),
		4993 => to_signed(15093, LUT_AMPL_WIDTH),
		4994 => to_signed(15096, LUT_AMPL_WIDTH),
		4995 => to_signed(15099, LUT_AMPL_WIDTH),
		4996 => to_signed(15102, LUT_AMPL_WIDTH),
		4997 => to_signed(15104, LUT_AMPL_WIDTH),
		4998 => to_signed(15107, LUT_AMPL_WIDTH),
		4999 => to_signed(15110, LUT_AMPL_WIDTH),
		5000 => to_signed(15113, LUT_AMPL_WIDTH),
		5001 => to_signed(15116, LUT_AMPL_WIDTH),
		5002 => to_signed(15118, LUT_AMPL_WIDTH),
		5003 => to_signed(15121, LUT_AMPL_WIDTH),
		5004 => to_signed(15124, LUT_AMPL_WIDTH),
		5005 => to_signed(15127, LUT_AMPL_WIDTH),
		5006 => to_signed(15129, LUT_AMPL_WIDTH),
		5007 => to_signed(15132, LUT_AMPL_WIDTH),
		5008 => to_signed(15135, LUT_AMPL_WIDTH),
		5009 => to_signed(15138, LUT_AMPL_WIDTH),
		5010 => to_signed(15141, LUT_AMPL_WIDTH),
		5011 => to_signed(15143, LUT_AMPL_WIDTH),
		5012 => to_signed(15146, LUT_AMPL_WIDTH),
		5013 => to_signed(15149, LUT_AMPL_WIDTH),
		5014 => to_signed(15152, LUT_AMPL_WIDTH),
		5015 => to_signed(15155, LUT_AMPL_WIDTH),
		5016 => to_signed(15157, LUT_AMPL_WIDTH),
		5017 => to_signed(15160, LUT_AMPL_WIDTH),
		5018 => to_signed(15163, LUT_AMPL_WIDTH),
		5019 => to_signed(15166, LUT_AMPL_WIDTH),
		5020 => to_signed(15168, LUT_AMPL_WIDTH),
		5021 => to_signed(15171, LUT_AMPL_WIDTH),
		5022 => to_signed(15174, LUT_AMPL_WIDTH),
		5023 => to_signed(15177, LUT_AMPL_WIDTH),
		5024 => to_signed(15180, LUT_AMPL_WIDTH),
		5025 => to_signed(15182, LUT_AMPL_WIDTH),
		5026 => to_signed(15185, LUT_AMPL_WIDTH),
		5027 => to_signed(15188, LUT_AMPL_WIDTH),
		5028 => to_signed(15191, LUT_AMPL_WIDTH),
		5029 => to_signed(15194, LUT_AMPL_WIDTH),
		5030 => to_signed(15196, LUT_AMPL_WIDTH),
		5031 => to_signed(15199, LUT_AMPL_WIDTH),
		5032 => to_signed(15202, LUT_AMPL_WIDTH),
		5033 => to_signed(15205, LUT_AMPL_WIDTH),
		5034 => to_signed(15207, LUT_AMPL_WIDTH),
		5035 => to_signed(15210, LUT_AMPL_WIDTH),
		5036 => to_signed(15213, LUT_AMPL_WIDTH),
		5037 => to_signed(15216, LUT_AMPL_WIDTH),
		5038 => to_signed(15219, LUT_AMPL_WIDTH),
		5039 => to_signed(15221, LUT_AMPL_WIDTH),
		5040 => to_signed(15224, LUT_AMPL_WIDTH),
		5041 => to_signed(15227, LUT_AMPL_WIDTH),
		5042 => to_signed(15230, LUT_AMPL_WIDTH),
		5043 => to_signed(15233, LUT_AMPL_WIDTH),
		5044 => to_signed(15235, LUT_AMPL_WIDTH),
		5045 => to_signed(15238, LUT_AMPL_WIDTH),
		5046 => to_signed(15241, LUT_AMPL_WIDTH),
		5047 => to_signed(15244, LUT_AMPL_WIDTH),
		5048 => to_signed(15246, LUT_AMPL_WIDTH),
		5049 => to_signed(15249, LUT_AMPL_WIDTH),
		5050 => to_signed(15252, LUT_AMPL_WIDTH),
		5051 => to_signed(15255, LUT_AMPL_WIDTH),
		5052 => to_signed(15258, LUT_AMPL_WIDTH),
		5053 => to_signed(15260, LUT_AMPL_WIDTH),
		5054 => to_signed(15263, LUT_AMPL_WIDTH),
		5055 => to_signed(15266, LUT_AMPL_WIDTH),
		5056 => to_signed(15269, LUT_AMPL_WIDTH),
		5057 => to_signed(15271, LUT_AMPL_WIDTH),
		5058 => to_signed(15274, LUT_AMPL_WIDTH),
		5059 => to_signed(15277, LUT_AMPL_WIDTH),
		5060 => to_signed(15280, LUT_AMPL_WIDTH),
		5061 => to_signed(15283, LUT_AMPL_WIDTH),
		5062 => to_signed(15285, LUT_AMPL_WIDTH),
		5063 => to_signed(15288, LUT_AMPL_WIDTH),
		5064 => to_signed(15291, LUT_AMPL_WIDTH),
		5065 => to_signed(15294, LUT_AMPL_WIDTH),
		5066 => to_signed(15296, LUT_AMPL_WIDTH),
		5067 => to_signed(15299, LUT_AMPL_WIDTH),
		5068 => to_signed(15302, LUT_AMPL_WIDTH),
		5069 => to_signed(15305, LUT_AMPL_WIDTH),
		5070 => to_signed(15308, LUT_AMPL_WIDTH),
		5071 => to_signed(15310, LUT_AMPL_WIDTH),
		5072 => to_signed(15313, LUT_AMPL_WIDTH),
		5073 => to_signed(15316, LUT_AMPL_WIDTH),
		5074 => to_signed(15319, LUT_AMPL_WIDTH),
		5075 => to_signed(15321, LUT_AMPL_WIDTH),
		5076 => to_signed(15324, LUT_AMPL_WIDTH),
		5077 => to_signed(15327, LUT_AMPL_WIDTH),
		5078 => to_signed(15330, LUT_AMPL_WIDTH),
		5079 => to_signed(15333, LUT_AMPL_WIDTH),
		5080 => to_signed(15335, LUT_AMPL_WIDTH),
		5081 => to_signed(15338, LUT_AMPL_WIDTH),
		5082 => to_signed(15341, LUT_AMPL_WIDTH),
		5083 => to_signed(15344, LUT_AMPL_WIDTH),
		5084 => to_signed(15346, LUT_AMPL_WIDTH),
		5085 => to_signed(15349, LUT_AMPL_WIDTH),
		5086 => to_signed(15352, LUT_AMPL_WIDTH),
		5087 => to_signed(15355, LUT_AMPL_WIDTH),
		5088 => to_signed(15358, LUT_AMPL_WIDTH),
		5089 => to_signed(15360, LUT_AMPL_WIDTH),
		5090 => to_signed(15363, LUT_AMPL_WIDTH),
		5091 => to_signed(15366, LUT_AMPL_WIDTH),
		5092 => to_signed(15369, LUT_AMPL_WIDTH),
		5093 => to_signed(15371, LUT_AMPL_WIDTH),
		5094 => to_signed(15374, LUT_AMPL_WIDTH),
		5095 => to_signed(15377, LUT_AMPL_WIDTH),
		5096 => to_signed(15380, LUT_AMPL_WIDTH),
		5097 => to_signed(15382, LUT_AMPL_WIDTH),
		5098 => to_signed(15385, LUT_AMPL_WIDTH),
		5099 => to_signed(15388, LUT_AMPL_WIDTH),
		5100 => to_signed(15391, LUT_AMPL_WIDTH),
		5101 => to_signed(15394, LUT_AMPL_WIDTH),
		5102 => to_signed(15396, LUT_AMPL_WIDTH),
		5103 => to_signed(15399, LUT_AMPL_WIDTH),
		5104 => to_signed(15402, LUT_AMPL_WIDTH),
		5105 => to_signed(15405, LUT_AMPL_WIDTH),
		5106 => to_signed(15407, LUT_AMPL_WIDTH),
		5107 => to_signed(15410, LUT_AMPL_WIDTH),
		5108 => to_signed(15413, LUT_AMPL_WIDTH),
		5109 => to_signed(15416, LUT_AMPL_WIDTH),
		5110 => to_signed(15419, LUT_AMPL_WIDTH),
		5111 => to_signed(15421, LUT_AMPL_WIDTH),
		5112 => to_signed(15424, LUT_AMPL_WIDTH),
		5113 => to_signed(15427, LUT_AMPL_WIDTH),
		5114 => to_signed(15430, LUT_AMPL_WIDTH),
		5115 => to_signed(15432, LUT_AMPL_WIDTH),
		5116 => to_signed(15435, LUT_AMPL_WIDTH),
		5117 => to_signed(15438, LUT_AMPL_WIDTH),
		5118 => to_signed(15441, LUT_AMPL_WIDTH),
		5119 => to_signed(15443, LUT_AMPL_WIDTH),
		5120 => to_signed(15446, LUT_AMPL_WIDTH),
		5121 => to_signed(15449, LUT_AMPL_WIDTH),
		5122 => to_signed(15452, LUT_AMPL_WIDTH),
		5123 => to_signed(15455, LUT_AMPL_WIDTH),
		5124 => to_signed(15457, LUT_AMPL_WIDTH),
		5125 => to_signed(15460, LUT_AMPL_WIDTH),
		5126 => to_signed(15463, LUT_AMPL_WIDTH),
		5127 => to_signed(15466, LUT_AMPL_WIDTH),
		5128 => to_signed(15468, LUT_AMPL_WIDTH),
		5129 => to_signed(15471, LUT_AMPL_WIDTH),
		5130 => to_signed(15474, LUT_AMPL_WIDTH),
		5131 => to_signed(15477, LUT_AMPL_WIDTH),
		5132 => to_signed(15479, LUT_AMPL_WIDTH),
		5133 => to_signed(15482, LUT_AMPL_WIDTH),
		5134 => to_signed(15485, LUT_AMPL_WIDTH),
		5135 => to_signed(15488, LUT_AMPL_WIDTH),
		5136 => to_signed(15491, LUT_AMPL_WIDTH),
		5137 => to_signed(15493, LUT_AMPL_WIDTH),
		5138 => to_signed(15496, LUT_AMPL_WIDTH),
		5139 => to_signed(15499, LUT_AMPL_WIDTH),
		5140 => to_signed(15502, LUT_AMPL_WIDTH),
		5141 => to_signed(15504, LUT_AMPL_WIDTH),
		5142 => to_signed(15507, LUT_AMPL_WIDTH),
		5143 => to_signed(15510, LUT_AMPL_WIDTH),
		5144 => to_signed(15513, LUT_AMPL_WIDTH),
		5145 => to_signed(15515, LUT_AMPL_WIDTH),
		5146 => to_signed(15518, LUT_AMPL_WIDTH),
		5147 => to_signed(15521, LUT_AMPL_WIDTH),
		5148 => to_signed(15524, LUT_AMPL_WIDTH),
		5149 => to_signed(15527, LUT_AMPL_WIDTH),
		5150 => to_signed(15529, LUT_AMPL_WIDTH),
		5151 => to_signed(15532, LUT_AMPL_WIDTH),
		5152 => to_signed(15535, LUT_AMPL_WIDTH),
		5153 => to_signed(15538, LUT_AMPL_WIDTH),
		5154 => to_signed(15540, LUT_AMPL_WIDTH),
		5155 => to_signed(15543, LUT_AMPL_WIDTH),
		5156 => to_signed(15546, LUT_AMPL_WIDTH),
		5157 => to_signed(15549, LUT_AMPL_WIDTH),
		5158 => to_signed(15551, LUT_AMPL_WIDTH),
		5159 => to_signed(15554, LUT_AMPL_WIDTH),
		5160 => to_signed(15557, LUT_AMPL_WIDTH),
		5161 => to_signed(15560, LUT_AMPL_WIDTH),
		5162 => to_signed(15562, LUT_AMPL_WIDTH),
		5163 => to_signed(15565, LUT_AMPL_WIDTH),
		5164 => to_signed(15568, LUT_AMPL_WIDTH),
		5165 => to_signed(15571, LUT_AMPL_WIDTH),
		5166 => to_signed(15574, LUT_AMPL_WIDTH),
		5167 => to_signed(15576, LUT_AMPL_WIDTH),
		5168 => to_signed(15579, LUT_AMPL_WIDTH),
		5169 => to_signed(15582, LUT_AMPL_WIDTH),
		5170 => to_signed(15585, LUT_AMPL_WIDTH),
		5171 => to_signed(15587, LUT_AMPL_WIDTH),
		5172 => to_signed(15590, LUT_AMPL_WIDTH),
		5173 => to_signed(15593, LUT_AMPL_WIDTH),
		5174 => to_signed(15596, LUT_AMPL_WIDTH),
		5175 => to_signed(15598, LUT_AMPL_WIDTH),
		5176 => to_signed(15601, LUT_AMPL_WIDTH),
		5177 => to_signed(15604, LUT_AMPL_WIDTH),
		5178 => to_signed(15607, LUT_AMPL_WIDTH),
		5179 => to_signed(15609, LUT_AMPL_WIDTH),
		5180 => to_signed(15612, LUT_AMPL_WIDTH),
		5181 => to_signed(15615, LUT_AMPL_WIDTH),
		5182 => to_signed(15618, LUT_AMPL_WIDTH),
		5183 => to_signed(15621, LUT_AMPL_WIDTH),
		5184 => to_signed(15623, LUT_AMPL_WIDTH),
		5185 => to_signed(15626, LUT_AMPL_WIDTH),
		5186 => to_signed(15629, LUT_AMPL_WIDTH),
		5187 => to_signed(15632, LUT_AMPL_WIDTH),
		5188 => to_signed(15634, LUT_AMPL_WIDTH),
		5189 => to_signed(15637, LUT_AMPL_WIDTH),
		5190 => to_signed(15640, LUT_AMPL_WIDTH),
		5191 => to_signed(15643, LUT_AMPL_WIDTH),
		5192 => to_signed(15645, LUT_AMPL_WIDTH),
		5193 => to_signed(15648, LUT_AMPL_WIDTH),
		5194 => to_signed(15651, LUT_AMPL_WIDTH),
		5195 => to_signed(15654, LUT_AMPL_WIDTH),
		5196 => to_signed(15656, LUT_AMPL_WIDTH),
		5197 => to_signed(15659, LUT_AMPL_WIDTH),
		5198 => to_signed(15662, LUT_AMPL_WIDTH),
		5199 => to_signed(15665, LUT_AMPL_WIDTH),
		5200 => to_signed(15667, LUT_AMPL_WIDTH),
		5201 => to_signed(15670, LUT_AMPL_WIDTH),
		5202 => to_signed(15673, LUT_AMPL_WIDTH),
		5203 => to_signed(15676, LUT_AMPL_WIDTH),
		5204 => to_signed(15678, LUT_AMPL_WIDTH),
		5205 => to_signed(15681, LUT_AMPL_WIDTH),
		5206 => to_signed(15684, LUT_AMPL_WIDTH),
		5207 => to_signed(15687, LUT_AMPL_WIDTH),
		5208 => to_signed(15690, LUT_AMPL_WIDTH),
		5209 => to_signed(15692, LUT_AMPL_WIDTH),
		5210 => to_signed(15695, LUT_AMPL_WIDTH),
		5211 => to_signed(15698, LUT_AMPL_WIDTH),
		5212 => to_signed(15701, LUT_AMPL_WIDTH),
		5213 => to_signed(15703, LUT_AMPL_WIDTH),
		5214 => to_signed(15706, LUT_AMPL_WIDTH),
		5215 => to_signed(15709, LUT_AMPL_WIDTH),
		5216 => to_signed(15712, LUT_AMPL_WIDTH),
		5217 => to_signed(15714, LUT_AMPL_WIDTH),
		5218 => to_signed(15717, LUT_AMPL_WIDTH),
		5219 => to_signed(15720, LUT_AMPL_WIDTH),
		5220 => to_signed(15723, LUT_AMPL_WIDTH),
		5221 => to_signed(15725, LUT_AMPL_WIDTH),
		5222 => to_signed(15728, LUT_AMPL_WIDTH),
		5223 => to_signed(15731, LUT_AMPL_WIDTH),
		5224 => to_signed(15734, LUT_AMPL_WIDTH),
		5225 => to_signed(15736, LUT_AMPL_WIDTH),
		5226 => to_signed(15739, LUT_AMPL_WIDTH),
		5227 => to_signed(15742, LUT_AMPL_WIDTH),
		5228 => to_signed(15745, LUT_AMPL_WIDTH),
		5229 => to_signed(15747, LUT_AMPL_WIDTH),
		5230 => to_signed(15750, LUT_AMPL_WIDTH),
		5231 => to_signed(15753, LUT_AMPL_WIDTH),
		5232 => to_signed(15756, LUT_AMPL_WIDTH),
		5233 => to_signed(15758, LUT_AMPL_WIDTH),
		5234 => to_signed(15761, LUT_AMPL_WIDTH),
		5235 => to_signed(15764, LUT_AMPL_WIDTH),
		5236 => to_signed(15767, LUT_AMPL_WIDTH),
		5237 => to_signed(15769, LUT_AMPL_WIDTH),
		5238 => to_signed(15772, LUT_AMPL_WIDTH),
		5239 => to_signed(15775, LUT_AMPL_WIDTH),
		5240 => to_signed(15778, LUT_AMPL_WIDTH),
		5241 => to_signed(15780, LUT_AMPL_WIDTH),
		5242 => to_signed(15783, LUT_AMPL_WIDTH),
		5243 => to_signed(15786, LUT_AMPL_WIDTH),
		5244 => to_signed(15789, LUT_AMPL_WIDTH),
		5245 => to_signed(15791, LUT_AMPL_WIDTH),
		5246 => to_signed(15794, LUT_AMPL_WIDTH),
		5247 => to_signed(15797, LUT_AMPL_WIDTH),
		5248 => to_signed(15800, LUT_AMPL_WIDTH),
		5249 => to_signed(15802, LUT_AMPL_WIDTH),
		5250 => to_signed(15805, LUT_AMPL_WIDTH),
		5251 => to_signed(15808, LUT_AMPL_WIDTH),
		5252 => to_signed(15811, LUT_AMPL_WIDTH),
		5253 => to_signed(15813, LUT_AMPL_WIDTH),
		5254 => to_signed(15816, LUT_AMPL_WIDTH),
		5255 => to_signed(15819, LUT_AMPL_WIDTH),
		5256 => to_signed(15822, LUT_AMPL_WIDTH),
		5257 => to_signed(15824, LUT_AMPL_WIDTH),
		5258 => to_signed(15827, LUT_AMPL_WIDTH),
		5259 => to_signed(15830, LUT_AMPL_WIDTH),
		5260 => to_signed(15833, LUT_AMPL_WIDTH),
		5261 => to_signed(15835, LUT_AMPL_WIDTH),
		5262 => to_signed(15838, LUT_AMPL_WIDTH),
		5263 => to_signed(15841, LUT_AMPL_WIDTH),
		5264 => to_signed(15844, LUT_AMPL_WIDTH),
		5265 => to_signed(15846, LUT_AMPL_WIDTH),
		5266 => to_signed(15849, LUT_AMPL_WIDTH),
		5267 => to_signed(15852, LUT_AMPL_WIDTH),
		5268 => to_signed(15855, LUT_AMPL_WIDTH),
		5269 => to_signed(15857, LUT_AMPL_WIDTH),
		5270 => to_signed(15860, LUT_AMPL_WIDTH),
		5271 => to_signed(15863, LUT_AMPL_WIDTH),
		5272 => to_signed(15866, LUT_AMPL_WIDTH),
		5273 => to_signed(15868, LUT_AMPL_WIDTH),
		5274 => to_signed(15871, LUT_AMPL_WIDTH),
		5275 => to_signed(15874, LUT_AMPL_WIDTH),
		5276 => to_signed(15877, LUT_AMPL_WIDTH),
		5277 => to_signed(15879, LUT_AMPL_WIDTH),
		5278 => to_signed(15882, LUT_AMPL_WIDTH),
		5279 => to_signed(15885, LUT_AMPL_WIDTH),
		5280 => to_signed(15888, LUT_AMPL_WIDTH),
		5281 => to_signed(15890, LUT_AMPL_WIDTH),
		5282 => to_signed(15893, LUT_AMPL_WIDTH),
		5283 => to_signed(15896, LUT_AMPL_WIDTH),
		5284 => to_signed(15899, LUT_AMPL_WIDTH),
		5285 => to_signed(15901, LUT_AMPL_WIDTH),
		5286 => to_signed(15904, LUT_AMPL_WIDTH),
		5287 => to_signed(15907, LUT_AMPL_WIDTH),
		5288 => to_signed(15910, LUT_AMPL_WIDTH),
		5289 => to_signed(15912, LUT_AMPL_WIDTH),
		5290 => to_signed(15915, LUT_AMPL_WIDTH),
		5291 => to_signed(15918, LUT_AMPL_WIDTH),
		5292 => to_signed(15921, LUT_AMPL_WIDTH),
		5293 => to_signed(15923, LUT_AMPL_WIDTH),
		5294 => to_signed(15926, LUT_AMPL_WIDTH),
		5295 => to_signed(15929, LUT_AMPL_WIDTH),
		5296 => to_signed(15932, LUT_AMPL_WIDTH),
		5297 => to_signed(15934, LUT_AMPL_WIDTH),
		5298 => to_signed(15937, LUT_AMPL_WIDTH),
		5299 => to_signed(15940, LUT_AMPL_WIDTH),
		5300 => to_signed(15943, LUT_AMPL_WIDTH),
		5301 => to_signed(15945, LUT_AMPL_WIDTH),
		5302 => to_signed(15948, LUT_AMPL_WIDTH),
		5303 => to_signed(15951, LUT_AMPL_WIDTH),
		5304 => to_signed(15954, LUT_AMPL_WIDTH),
		5305 => to_signed(15956, LUT_AMPL_WIDTH),
		5306 => to_signed(15959, LUT_AMPL_WIDTH),
		5307 => to_signed(15962, LUT_AMPL_WIDTH),
		5308 => to_signed(15965, LUT_AMPL_WIDTH),
		5309 => to_signed(15967, LUT_AMPL_WIDTH),
		5310 => to_signed(15970, LUT_AMPL_WIDTH),
		5311 => to_signed(15973, LUT_AMPL_WIDTH),
		5312 => to_signed(15976, LUT_AMPL_WIDTH),
		5313 => to_signed(15978, LUT_AMPL_WIDTH),
		5314 => to_signed(15981, LUT_AMPL_WIDTH),
		5315 => to_signed(15984, LUT_AMPL_WIDTH),
		5316 => to_signed(15987, LUT_AMPL_WIDTH),
		5317 => to_signed(15989, LUT_AMPL_WIDTH),
		5318 => to_signed(15992, LUT_AMPL_WIDTH),
		5319 => to_signed(15995, LUT_AMPL_WIDTH),
		5320 => to_signed(15997, LUT_AMPL_WIDTH),
		5321 => to_signed(16000, LUT_AMPL_WIDTH),
		5322 => to_signed(16003, LUT_AMPL_WIDTH),
		5323 => to_signed(16006, LUT_AMPL_WIDTH),
		5324 => to_signed(16008, LUT_AMPL_WIDTH),
		5325 => to_signed(16011, LUT_AMPL_WIDTH),
		5326 => to_signed(16014, LUT_AMPL_WIDTH),
		5327 => to_signed(16017, LUT_AMPL_WIDTH),
		5328 => to_signed(16019, LUT_AMPL_WIDTH),
		5329 => to_signed(16022, LUT_AMPL_WIDTH),
		5330 => to_signed(16025, LUT_AMPL_WIDTH),
		5331 => to_signed(16028, LUT_AMPL_WIDTH),
		5332 => to_signed(16030, LUT_AMPL_WIDTH),
		5333 => to_signed(16033, LUT_AMPL_WIDTH),
		5334 => to_signed(16036, LUT_AMPL_WIDTH),
		5335 => to_signed(16039, LUT_AMPL_WIDTH),
		5336 => to_signed(16041, LUT_AMPL_WIDTH),
		5337 => to_signed(16044, LUT_AMPL_WIDTH),
		5338 => to_signed(16047, LUT_AMPL_WIDTH),
		5339 => to_signed(16050, LUT_AMPL_WIDTH),
		5340 => to_signed(16052, LUT_AMPL_WIDTH),
		5341 => to_signed(16055, LUT_AMPL_WIDTH),
		5342 => to_signed(16058, LUT_AMPL_WIDTH),
		5343 => to_signed(16061, LUT_AMPL_WIDTH),
		5344 => to_signed(16063, LUT_AMPL_WIDTH),
		5345 => to_signed(16066, LUT_AMPL_WIDTH),
		5346 => to_signed(16069, LUT_AMPL_WIDTH),
		5347 => to_signed(16071, LUT_AMPL_WIDTH),
		5348 => to_signed(16074, LUT_AMPL_WIDTH),
		5349 => to_signed(16077, LUT_AMPL_WIDTH),
		5350 => to_signed(16080, LUT_AMPL_WIDTH),
		5351 => to_signed(16082, LUT_AMPL_WIDTH),
		5352 => to_signed(16085, LUT_AMPL_WIDTH),
		5353 => to_signed(16088, LUT_AMPL_WIDTH),
		5354 => to_signed(16091, LUT_AMPL_WIDTH),
		5355 => to_signed(16093, LUT_AMPL_WIDTH),
		5356 => to_signed(16096, LUT_AMPL_WIDTH),
		5357 => to_signed(16099, LUT_AMPL_WIDTH),
		5358 => to_signed(16102, LUT_AMPL_WIDTH),
		5359 => to_signed(16104, LUT_AMPL_WIDTH),
		5360 => to_signed(16107, LUT_AMPL_WIDTH),
		5361 => to_signed(16110, LUT_AMPL_WIDTH),
		5362 => to_signed(16113, LUT_AMPL_WIDTH),
		5363 => to_signed(16115, LUT_AMPL_WIDTH),
		5364 => to_signed(16118, LUT_AMPL_WIDTH),
		5365 => to_signed(16121, LUT_AMPL_WIDTH),
		5366 => to_signed(16123, LUT_AMPL_WIDTH),
		5367 => to_signed(16126, LUT_AMPL_WIDTH),
		5368 => to_signed(16129, LUT_AMPL_WIDTH),
		5369 => to_signed(16132, LUT_AMPL_WIDTH),
		5370 => to_signed(16134, LUT_AMPL_WIDTH),
		5371 => to_signed(16137, LUT_AMPL_WIDTH),
		5372 => to_signed(16140, LUT_AMPL_WIDTH),
		5373 => to_signed(16143, LUT_AMPL_WIDTH),
		5374 => to_signed(16145, LUT_AMPL_WIDTH),
		5375 => to_signed(16148, LUT_AMPL_WIDTH),
		5376 => to_signed(16151, LUT_AMPL_WIDTH),
		5377 => to_signed(16154, LUT_AMPL_WIDTH),
		5378 => to_signed(16156, LUT_AMPL_WIDTH),
		5379 => to_signed(16159, LUT_AMPL_WIDTH),
		5380 => to_signed(16162, LUT_AMPL_WIDTH),
		5381 => to_signed(16164, LUT_AMPL_WIDTH),
		5382 => to_signed(16167, LUT_AMPL_WIDTH),
		5383 => to_signed(16170, LUT_AMPL_WIDTH),
		5384 => to_signed(16173, LUT_AMPL_WIDTH),
		5385 => to_signed(16175, LUT_AMPL_WIDTH),
		5386 => to_signed(16178, LUT_AMPL_WIDTH),
		5387 => to_signed(16181, LUT_AMPL_WIDTH),
		5388 => to_signed(16184, LUT_AMPL_WIDTH),
		5389 => to_signed(16186, LUT_AMPL_WIDTH),
		5390 => to_signed(16189, LUT_AMPL_WIDTH),
		5391 => to_signed(16192, LUT_AMPL_WIDTH),
		5392 => to_signed(16195, LUT_AMPL_WIDTH),
		5393 => to_signed(16197, LUT_AMPL_WIDTH),
		5394 => to_signed(16200, LUT_AMPL_WIDTH),
		5395 => to_signed(16203, LUT_AMPL_WIDTH),
		5396 => to_signed(16205, LUT_AMPL_WIDTH),
		5397 => to_signed(16208, LUT_AMPL_WIDTH),
		5398 => to_signed(16211, LUT_AMPL_WIDTH),
		5399 => to_signed(16214, LUT_AMPL_WIDTH),
		5400 => to_signed(16216, LUT_AMPL_WIDTH),
		5401 => to_signed(16219, LUT_AMPL_WIDTH),
		5402 => to_signed(16222, LUT_AMPL_WIDTH),
		5403 => to_signed(16225, LUT_AMPL_WIDTH),
		5404 => to_signed(16227, LUT_AMPL_WIDTH),
		5405 => to_signed(16230, LUT_AMPL_WIDTH),
		5406 => to_signed(16233, LUT_AMPL_WIDTH),
		5407 => to_signed(16235, LUT_AMPL_WIDTH),
		5408 => to_signed(16238, LUT_AMPL_WIDTH),
		5409 => to_signed(16241, LUT_AMPL_WIDTH),
		5410 => to_signed(16244, LUT_AMPL_WIDTH),
		5411 => to_signed(16246, LUT_AMPL_WIDTH),
		5412 => to_signed(16249, LUT_AMPL_WIDTH),
		5413 => to_signed(16252, LUT_AMPL_WIDTH),
		5414 => to_signed(16255, LUT_AMPL_WIDTH),
		5415 => to_signed(16257, LUT_AMPL_WIDTH),
		5416 => to_signed(16260, LUT_AMPL_WIDTH),
		5417 => to_signed(16263, LUT_AMPL_WIDTH),
		5418 => to_signed(16265, LUT_AMPL_WIDTH),
		5419 => to_signed(16268, LUT_AMPL_WIDTH),
		5420 => to_signed(16271, LUT_AMPL_WIDTH),
		5421 => to_signed(16274, LUT_AMPL_WIDTH),
		5422 => to_signed(16276, LUT_AMPL_WIDTH),
		5423 => to_signed(16279, LUT_AMPL_WIDTH),
		5424 => to_signed(16282, LUT_AMPL_WIDTH),
		5425 => to_signed(16285, LUT_AMPL_WIDTH),
		5426 => to_signed(16287, LUT_AMPL_WIDTH),
		5427 => to_signed(16290, LUT_AMPL_WIDTH),
		5428 => to_signed(16293, LUT_AMPL_WIDTH),
		5429 => to_signed(16295, LUT_AMPL_WIDTH),
		5430 => to_signed(16298, LUT_AMPL_WIDTH),
		5431 => to_signed(16301, LUT_AMPL_WIDTH),
		5432 => to_signed(16304, LUT_AMPL_WIDTH),
		5433 => to_signed(16306, LUT_AMPL_WIDTH),
		5434 => to_signed(16309, LUT_AMPL_WIDTH),
		5435 => to_signed(16312, LUT_AMPL_WIDTH),
		5436 => to_signed(16315, LUT_AMPL_WIDTH),
		5437 => to_signed(16317, LUT_AMPL_WIDTH),
		5438 => to_signed(16320, LUT_AMPL_WIDTH),
		5439 => to_signed(16323, LUT_AMPL_WIDTH),
		5440 => to_signed(16325, LUT_AMPL_WIDTH),
		5441 => to_signed(16328, LUT_AMPL_WIDTH),
		5442 => to_signed(16331, LUT_AMPL_WIDTH),
		5443 => to_signed(16334, LUT_AMPL_WIDTH),
		5444 => to_signed(16336, LUT_AMPL_WIDTH),
		5445 => to_signed(16339, LUT_AMPL_WIDTH),
		5446 => to_signed(16342, LUT_AMPL_WIDTH),
		5447 => to_signed(16344, LUT_AMPL_WIDTH),
		5448 => to_signed(16347, LUT_AMPL_WIDTH),
		5449 => to_signed(16350, LUT_AMPL_WIDTH),
		5450 => to_signed(16353, LUT_AMPL_WIDTH),
		5451 => to_signed(16355, LUT_AMPL_WIDTH),
		5452 => to_signed(16358, LUT_AMPL_WIDTH),
		5453 => to_signed(16361, LUT_AMPL_WIDTH),
		5454 => to_signed(16364, LUT_AMPL_WIDTH),
		5455 => to_signed(16366, LUT_AMPL_WIDTH),
		5456 => to_signed(16369, LUT_AMPL_WIDTH),
		5457 => to_signed(16372, LUT_AMPL_WIDTH),
		5458 => to_signed(16374, LUT_AMPL_WIDTH),
		5459 => to_signed(16377, LUT_AMPL_WIDTH),
		5460 => to_signed(16380, LUT_AMPL_WIDTH),
		5461 => to_signed(16383, LUT_AMPL_WIDTH),
		5462 => to_signed(16385, LUT_AMPL_WIDTH),
		5463 => to_signed(16388, LUT_AMPL_WIDTH),
		5464 => to_signed(16391, LUT_AMPL_WIDTH),
		5465 => to_signed(16393, LUT_AMPL_WIDTH),
		5466 => to_signed(16396, LUT_AMPL_WIDTH),
		5467 => to_signed(16399, LUT_AMPL_WIDTH),
		5468 => to_signed(16402, LUT_AMPL_WIDTH),
		5469 => to_signed(16404, LUT_AMPL_WIDTH),
		5470 => to_signed(16407, LUT_AMPL_WIDTH),
		5471 => to_signed(16410, LUT_AMPL_WIDTH),
		5472 => to_signed(16413, LUT_AMPL_WIDTH),
		5473 => to_signed(16415, LUT_AMPL_WIDTH),
		5474 => to_signed(16418, LUT_AMPL_WIDTH),
		5475 => to_signed(16421, LUT_AMPL_WIDTH),
		5476 => to_signed(16423, LUT_AMPL_WIDTH),
		5477 => to_signed(16426, LUT_AMPL_WIDTH),
		5478 => to_signed(16429, LUT_AMPL_WIDTH),
		5479 => to_signed(16432, LUT_AMPL_WIDTH),
		5480 => to_signed(16434, LUT_AMPL_WIDTH),
		5481 => to_signed(16437, LUT_AMPL_WIDTH),
		5482 => to_signed(16440, LUT_AMPL_WIDTH),
		5483 => to_signed(16442, LUT_AMPL_WIDTH),
		5484 => to_signed(16445, LUT_AMPL_WIDTH),
		5485 => to_signed(16448, LUT_AMPL_WIDTH),
		5486 => to_signed(16451, LUT_AMPL_WIDTH),
		5487 => to_signed(16453, LUT_AMPL_WIDTH),
		5488 => to_signed(16456, LUT_AMPL_WIDTH),
		5489 => to_signed(16459, LUT_AMPL_WIDTH),
		5490 => to_signed(16461, LUT_AMPL_WIDTH),
		5491 => to_signed(16464, LUT_AMPL_WIDTH),
		5492 => to_signed(16467, LUT_AMPL_WIDTH),
		5493 => to_signed(16470, LUT_AMPL_WIDTH),
		5494 => to_signed(16472, LUT_AMPL_WIDTH),
		5495 => to_signed(16475, LUT_AMPL_WIDTH),
		5496 => to_signed(16478, LUT_AMPL_WIDTH),
		5497 => to_signed(16480, LUT_AMPL_WIDTH),
		5498 => to_signed(16483, LUT_AMPL_WIDTH),
		5499 => to_signed(16486, LUT_AMPL_WIDTH),
		5500 => to_signed(16489, LUT_AMPL_WIDTH),
		5501 => to_signed(16491, LUT_AMPL_WIDTH),
		5502 => to_signed(16494, LUT_AMPL_WIDTH),
		5503 => to_signed(16497, LUT_AMPL_WIDTH),
		5504 => to_signed(16499, LUT_AMPL_WIDTH),
		5505 => to_signed(16502, LUT_AMPL_WIDTH),
		5506 => to_signed(16505, LUT_AMPL_WIDTH),
		5507 => to_signed(16508, LUT_AMPL_WIDTH),
		5508 => to_signed(16510, LUT_AMPL_WIDTH),
		5509 => to_signed(16513, LUT_AMPL_WIDTH),
		5510 => to_signed(16516, LUT_AMPL_WIDTH),
		5511 => to_signed(16518, LUT_AMPL_WIDTH),
		5512 => to_signed(16521, LUT_AMPL_WIDTH),
		5513 => to_signed(16524, LUT_AMPL_WIDTH),
		5514 => to_signed(16527, LUT_AMPL_WIDTH),
		5515 => to_signed(16529, LUT_AMPL_WIDTH),
		5516 => to_signed(16532, LUT_AMPL_WIDTH),
		5517 => to_signed(16535, LUT_AMPL_WIDTH),
		5518 => to_signed(16537, LUT_AMPL_WIDTH),
		5519 => to_signed(16540, LUT_AMPL_WIDTH),
		5520 => to_signed(16543, LUT_AMPL_WIDTH),
		5521 => to_signed(16546, LUT_AMPL_WIDTH),
		5522 => to_signed(16548, LUT_AMPL_WIDTH),
		5523 => to_signed(16551, LUT_AMPL_WIDTH),
		5524 => to_signed(16554, LUT_AMPL_WIDTH),
		5525 => to_signed(16556, LUT_AMPL_WIDTH),
		5526 => to_signed(16559, LUT_AMPL_WIDTH),
		5527 => to_signed(16562, LUT_AMPL_WIDTH),
		5528 => to_signed(16565, LUT_AMPL_WIDTH),
		5529 => to_signed(16567, LUT_AMPL_WIDTH),
		5530 => to_signed(16570, LUT_AMPL_WIDTH),
		5531 => to_signed(16573, LUT_AMPL_WIDTH),
		5532 => to_signed(16575, LUT_AMPL_WIDTH),
		5533 => to_signed(16578, LUT_AMPL_WIDTH),
		5534 => to_signed(16581, LUT_AMPL_WIDTH),
		5535 => to_signed(16584, LUT_AMPL_WIDTH),
		5536 => to_signed(16586, LUT_AMPL_WIDTH),
		5537 => to_signed(16589, LUT_AMPL_WIDTH),
		5538 => to_signed(16592, LUT_AMPL_WIDTH),
		5539 => to_signed(16594, LUT_AMPL_WIDTH),
		5540 => to_signed(16597, LUT_AMPL_WIDTH),
		5541 => to_signed(16600, LUT_AMPL_WIDTH),
		5542 => to_signed(16602, LUT_AMPL_WIDTH),
		5543 => to_signed(16605, LUT_AMPL_WIDTH),
		5544 => to_signed(16608, LUT_AMPL_WIDTH),
		5545 => to_signed(16611, LUT_AMPL_WIDTH),
		5546 => to_signed(16613, LUT_AMPL_WIDTH),
		5547 => to_signed(16616, LUT_AMPL_WIDTH),
		5548 => to_signed(16619, LUT_AMPL_WIDTH),
		5549 => to_signed(16621, LUT_AMPL_WIDTH),
		5550 => to_signed(16624, LUT_AMPL_WIDTH),
		5551 => to_signed(16627, LUT_AMPL_WIDTH),
		5552 => to_signed(16630, LUT_AMPL_WIDTH),
		5553 => to_signed(16632, LUT_AMPL_WIDTH),
		5554 => to_signed(16635, LUT_AMPL_WIDTH),
		5555 => to_signed(16638, LUT_AMPL_WIDTH),
		5556 => to_signed(16640, LUT_AMPL_WIDTH),
		5557 => to_signed(16643, LUT_AMPL_WIDTH),
		5558 => to_signed(16646, LUT_AMPL_WIDTH),
		5559 => to_signed(16648, LUT_AMPL_WIDTH),
		5560 => to_signed(16651, LUT_AMPL_WIDTH),
		5561 => to_signed(16654, LUT_AMPL_WIDTH),
		5562 => to_signed(16657, LUT_AMPL_WIDTH),
		5563 => to_signed(16659, LUT_AMPL_WIDTH),
		5564 => to_signed(16662, LUT_AMPL_WIDTH),
		5565 => to_signed(16665, LUT_AMPL_WIDTH),
		5566 => to_signed(16667, LUT_AMPL_WIDTH),
		5567 => to_signed(16670, LUT_AMPL_WIDTH),
		5568 => to_signed(16673, LUT_AMPL_WIDTH),
		5569 => to_signed(16676, LUT_AMPL_WIDTH),
		5570 => to_signed(16678, LUT_AMPL_WIDTH),
		5571 => to_signed(16681, LUT_AMPL_WIDTH),
		5572 => to_signed(16684, LUT_AMPL_WIDTH),
		5573 => to_signed(16686, LUT_AMPL_WIDTH),
		5574 => to_signed(16689, LUT_AMPL_WIDTH),
		5575 => to_signed(16692, LUT_AMPL_WIDTH),
		5576 => to_signed(16694, LUT_AMPL_WIDTH),
		5577 => to_signed(16697, LUT_AMPL_WIDTH),
		5578 => to_signed(16700, LUT_AMPL_WIDTH),
		5579 => to_signed(16703, LUT_AMPL_WIDTH),
		5580 => to_signed(16705, LUT_AMPL_WIDTH),
		5581 => to_signed(16708, LUT_AMPL_WIDTH),
		5582 => to_signed(16711, LUT_AMPL_WIDTH),
		5583 => to_signed(16713, LUT_AMPL_WIDTH),
		5584 => to_signed(16716, LUT_AMPL_WIDTH),
		5585 => to_signed(16719, LUT_AMPL_WIDTH),
		5586 => to_signed(16721, LUT_AMPL_WIDTH),
		5587 => to_signed(16724, LUT_AMPL_WIDTH),
		5588 => to_signed(16727, LUT_AMPL_WIDTH),
		5589 => to_signed(16730, LUT_AMPL_WIDTH),
		5590 => to_signed(16732, LUT_AMPL_WIDTH),
		5591 => to_signed(16735, LUT_AMPL_WIDTH),
		5592 => to_signed(16738, LUT_AMPL_WIDTH),
		5593 => to_signed(16740, LUT_AMPL_WIDTH),
		5594 => to_signed(16743, LUT_AMPL_WIDTH),
		5595 => to_signed(16746, LUT_AMPL_WIDTH),
		5596 => to_signed(16749, LUT_AMPL_WIDTH),
		5597 => to_signed(16751, LUT_AMPL_WIDTH),
		5598 => to_signed(16754, LUT_AMPL_WIDTH),
		5599 => to_signed(16757, LUT_AMPL_WIDTH),
		5600 => to_signed(16759, LUT_AMPL_WIDTH),
		5601 => to_signed(16762, LUT_AMPL_WIDTH),
		5602 => to_signed(16765, LUT_AMPL_WIDTH),
		5603 => to_signed(16767, LUT_AMPL_WIDTH),
		5604 => to_signed(16770, LUT_AMPL_WIDTH),
		5605 => to_signed(16773, LUT_AMPL_WIDTH),
		5606 => to_signed(16775, LUT_AMPL_WIDTH),
		5607 => to_signed(16778, LUT_AMPL_WIDTH),
		5608 => to_signed(16781, LUT_AMPL_WIDTH),
		5609 => to_signed(16784, LUT_AMPL_WIDTH),
		5610 => to_signed(16786, LUT_AMPL_WIDTH),
		5611 => to_signed(16789, LUT_AMPL_WIDTH),
		5612 => to_signed(16792, LUT_AMPL_WIDTH),
		5613 => to_signed(16794, LUT_AMPL_WIDTH),
		5614 => to_signed(16797, LUT_AMPL_WIDTH),
		5615 => to_signed(16800, LUT_AMPL_WIDTH),
		5616 => to_signed(16802, LUT_AMPL_WIDTH),
		5617 => to_signed(16805, LUT_AMPL_WIDTH),
		5618 => to_signed(16808, LUT_AMPL_WIDTH),
		5619 => to_signed(16811, LUT_AMPL_WIDTH),
		5620 => to_signed(16813, LUT_AMPL_WIDTH),
		5621 => to_signed(16816, LUT_AMPL_WIDTH),
		5622 => to_signed(16819, LUT_AMPL_WIDTH),
		5623 => to_signed(16821, LUT_AMPL_WIDTH),
		5624 => to_signed(16824, LUT_AMPL_WIDTH),
		5625 => to_signed(16827, LUT_AMPL_WIDTH),
		5626 => to_signed(16829, LUT_AMPL_WIDTH),
		5627 => to_signed(16832, LUT_AMPL_WIDTH),
		5628 => to_signed(16835, LUT_AMPL_WIDTH),
		5629 => to_signed(16838, LUT_AMPL_WIDTH),
		5630 => to_signed(16840, LUT_AMPL_WIDTH),
		5631 => to_signed(16843, LUT_AMPL_WIDTH),
		5632 => to_signed(16846, LUT_AMPL_WIDTH),
		5633 => to_signed(16848, LUT_AMPL_WIDTH),
		5634 => to_signed(16851, LUT_AMPL_WIDTH),
		5635 => to_signed(16854, LUT_AMPL_WIDTH),
		5636 => to_signed(16856, LUT_AMPL_WIDTH),
		5637 => to_signed(16859, LUT_AMPL_WIDTH),
		5638 => to_signed(16862, LUT_AMPL_WIDTH),
		5639 => to_signed(16864, LUT_AMPL_WIDTH),
		5640 => to_signed(16867, LUT_AMPL_WIDTH),
		5641 => to_signed(16870, LUT_AMPL_WIDTH),
		5642 => to_signed(16873, LUT_AMPL_WIDTH),
		5643 => to_signed(16875, LUT_AMPL_WIDTH),
		5644 => to_signed(16878, LUT_AMPL_WIDTH),
		5645 => to_signed(16881, LUT_AMPL_WIDTH),
		5646 => to_signed(16883, LUT_AMPL_WIDTH),
		5647 => to_signed(16886, LUT_AMPL_WIDTH),
		5648 => to_signed(16889, LUT_AMPL_WIDTH),
		5649 => to_signed(16891, LUT_AMPL_WIDTH),
		5650 => to_signed(16894, LUT_AMPL_WIDTH),
		5651 => to_signed(16897, LUT_AMPL_WIDTH),
		5652 => to_signed(16899, LUT_AMPL_WIDTH),
		5653 => to_signed(16902, LUT_AMPL_WIDTH),
		5654 => to_signed(16905, LUT_AMPL_WIDTH),
		5655 => to_signed(16908, LUT_AMPL_WIDTH),
		5656 => to_signed(16910, LUT_AMPL_WIDTH),
		5657 => to_signed(16913, LUT_AMPL_WIDTH),
		5658 => to_signed(16916, LUT_AMPL_WIDTH),
		5659 => to_signed(16918, LUT_AMPL_WIDTH),
		5660 => to_signed(16921, LUT_AMPL_WIDTH),
		5661 => to_signed(16924, LUT_AMPL_WIDTH),
		5662 => to_signed(16926, LUT_AMPL_WIDTH),
		5663 => to_signed(16929, LUT_AMPL_WIDTH),
		5664 => to_signed(16932, LUT_AMPL_WIDTH),
		5665 => to_signed(16934, LUT_AMPL_WIDTH),
		5666 => to_signed(16937, LUT_AMPL_WIDTH),
		5667 => to_signed(16940, LUT_AMPL_WIDTH),
		5668 => to_signed(16943, LUT_AMPL_WIDTH),
		5669 => to_signed(16945, LUT_AMPL_WIDTH),
		5670 => to_signed(16948, LUT_AMPL_WIDTH),
		5671 => to_signed(16951, LUT_AMPL_WIDTH),
		5672 => to_signed(16953, LUT_AMPL_WIDTH),
		5673 => to_signed(16956, LUT_AMPL_WIDTH),
		5674 => to_signed(16959, LUT_AMPL_WIDTH),
		5675 => to_signed(16961, LUT_AMPL_WIDTH),
		5676 => to_signed(16964, LUT_AMPL_WIDTH),
		5677 => to_signed(16967, LUT_AMPL_WIDTH),
		5678 => to_signed(16969, LUT_AMPL_WIDTH),
		5679 => to_signed(16972, LUT_AMPL_WIDTH),
		5680 => to_signed(16975, LUT_AMPL_WIDTH),
		5681 => to_signed(16977, LUT_AMPL_WIDTH),
		5682 => to_signed(16980, LUT_AMPL_WIDTH),
		5683 => to_signed(16983, LUT_AMPL_WIDTH),
		5684 => to_signed(16986, LUT_AMPL_WIDTH),
		5685 => to_signed(16988, LUT_AMPL_WIDTH),
		5686 => to_signed(16991, LUT_AMPL_WIDTH),
		5687 => to_signed(16994, LUT_AMPL_WIDTH),
		5688 => to_signed(16996, LUT_AMPL_WIDTH),
		5689 => to_signed(16999, LUT_AMPL_WIDTH),
		5690 => to_signed(17002, LUT_AMPL_WIDTH),
		5691 => to_signed(17004, LUT_AMPL_WIDTH),
		5692 => to_signed(17007, LUT_AMPL_WIDTH),
		5693 => to_signed(17010, LUT_AMPL_WIDTH),
		5694 => to_signed(17012, LUT_AMPL_WIDTH),
		5695 => to_signed(17015, LUT_AMPL_WIDTH),
		5696 => to_signed(17018, LUT_AMPL_WIDTH),
		5697 => to_signed(17020, LUT_AMPL_WIDTH),
		5698 => to_signed(17023, LUT_AMPL_WIDTH),
		5699 => to_signed(17026, LUT_AMPL_WIDTH),
		5700 => to_signed(17028, LUT_AMPL_WIDTH),
		5701 => to_signed(17031, LUT_AMPL_WIDTH),
		5702 => to_signed(17034, LUT_AMPL_WIDTH),
		5703 => to_signed(17037, LUT_AMPL_WIDTH),
		5704 => to_signed(17039, LUT_AMPL_WIDTH),
		5705 => to_signed(17042, LUT_AMPL_WIDTH),
		5706 => to_signed(17045, LUT_AMPL_WIDTH),
		5707 => to_signed(17047, LUT_AMPL_WIDTH),
		5708 => to_signed(17050, LUT_AMPL_WIDTH),
		5709 => to_signed(17053, LUT_AMPL_WIDTH),
		5710 => to_signed(17055, LUT_AMPL_WIDTH),
		5711 => to_signed(17058, LUT_AMPL_WIDTH),
		5712 => to_signed(17061, LUT_AMPL_WIDTH),
		5713 => to_signed(17063, LUT_AMPL_WIDTH),
		5714 => to_signed(17066, LUT_AMPL_WIDTH),
		5715 => to_signed(17069, LUT_AMPL_WIDTH),
		5716 => to_signed(17071, LUT_AMPL_WIDTH),
		5717 => to_signed(17074, LUT_AMPL_WIDTH),
		5718 => to_signed(17077, LUT_AMPL_WIDTH),
		5719 => to_signed(17079, LUT_AMPL_WIDTH),
		5720 => to_signed(17082, LUT_AMPL_WIDTH),
		5721 => to_signed(17085, LUT_AMPL_WIDTH),
		5722 => to_signed(17087, LUT_AMPL_WIDTH),
		5723 => to_signed(17090, LUT_AMPL_WIDTH),
		5724 => to_signed(17093, LUT_AMPL_WIDTH),
		5725 => to_signed(17096, LUT_AMPL_WIDTH),
		5726 => to_signed(17098, LUT_AMPL_WIDTH),
		5727 => to_signed(17101, LUT_AMPL_WIDTH),
		5728 => to_signed(17104, LUT_AMPL_WIDTH),
		5729 => to_signed(17106, LUT_AMPL_WIDTH),
		5730 => to_signed(17109, LUT_AMPL_WIDTH),
		5731 => to_signed(17112, LUT_AMPL_WIDTH),
		5732 => to_signed(17114, LUT_AMPL_WIDTH),
		5733 => to_signed(17117, LUT_AMPL_WIDTH),
		5734 => to_signed(17120, LUT_AMPL_WIDTH),
		5735 => to_signed(17122, LUT_AMPL_WIDTH),
		5736 => to_signed(17125, LUT_AMPL_WIDTH),
		5737 => to_signed(17128, LUT_AMPL_WIDTH),
		5738 => to_signed(17130, LUT_AMPL_WIDTH),
		5739 => to_signed(17133, LUT_AMPL_WIDTH),
		5740 => to_signed(17136, LUT_AMPL_WIDTH),
		5741 => to_signed(17138, LUT_AMPL_WIDTH),
		5742 => to_signed(17141, LUT_AMPL_WIDTH),
		5743 => to_signed(17144, LUT_AMPL_WIDTH),
		5744 => to_signed(17146, LUT_AMPL_WIDTH),
		5745 => to_signed(17149, LUT_AMPL_WIDTH),
		5746 => to_signed(17152, LUT_AMPL_WIDTH),
		5747 => to_signed(17154, LUT_AMPL_WIDTH),
		5748 => to_signed(17157, LUT_AMPL_WIDTH),
		5749 => to_signed(17160, LUT_AMPL_WIDTH),
		5750 => to_signed(17162, LUT_AMPL_WIDTH),
		5751 => to_signed(17165, LUT_AMPL_WIDTH),
		5752 => to_signed(17168, LUT_AMPL_WIDTH),
		5753 => to_signed(17171, LUT_AMPL_WIDTH),
		5754 => to_signed(17173, LUT_AMPL_WIDTH),
		5755 => to_signed(17176, LUT_AMPL_WIDTH),
		5756 => to_signed(17179, LUT_AMPL_WIDTH),
		5757 => to_signed(17181, LUT_AMPL_WIDTH),
		5758 => to_signed(17184, LUT_AMPL_WIDTH),
		5759 => to_signed(17187, LUT_AMPL_WIDTH),
		5760 => to_signed(17189, LUT_AMPL_WIDTH),
		5761 => to_signed(17192, LUT_AMPL_WIDTH),
		5762 => to_signed(17195, LUT_AMPL_WIDTH),
		5763 => to_signed(17197, LUT_AMPL_WIDTH),
		5764 => to_signed(17200, LUT_AMPL_WIDTH),
		5765 => to_signed(17203, LUT_AMPL_WIDTH),
		5766 => to_signed(17205, LUT_AMPL_WIDTH),
		5767 => to_signed(17208, LUT_AMPL_WIDTH),
		5768 => to_signed(17211, LUT_AMPL_WIDTH),
		5769 => to_signed(17213, LUT_AMPL_WIDTH),
		5770 => to_signed(17216, LUT_AMPL_WIDTH),
		5771 => to_signed(17219, LUT_AMPL_WIDTH),
		5772 => to_signed(17221, LUT_AMPL_WIDTH),
		5773 => to_signed(17224, LUT_AMPL_WIDTH),
		5774 => to_signed(17227, LUT_AMPL_WIDTH),
		5775 => to_signed(17229, LUT_AMPL_WIDTH),
		5776 => to_signed(17232, LUT_AMPL_WIDTH),
		5777 => to_signed(17235, LUT_AMPL_WIDTH),
		5778 => to_signed(17237, LUT_AMPL_WIDTH),
		5779 => to_signed(17240, LUT_AMPL_WIDTH),
		5780 => to_signed(17243, LUT_AMPL_WIDTH),
		5781 => to_signed(17245, LUT_AMPL_WIDTH),
		5782 => to_signed(17248, LUT_AMPL_WIDTH),
		5783 => to_signed(17251, LUT_AMPL_WIDTH),
		5784 => to_signed(17253, LUT_AMPL_WIDTH),
		5785 => to_signed(17256, LUT_AMPL_WIDTH),
		5786 => to_signed(17259, LUT_AMPL_WIDTH),
		5787 => to_signed(17261, LUT_AMPL_WIDTH),
		5788 => to_signed(17264, LUT_AMPL_WIDTH),
		5789 => to_signed(17267, LUT_AMPL_WIDTH),
		5790 => to_signed(17269, LUT_AMPL_WIDTH),
		5791 => to_signed(17272, LUT_AMPL_WIDTH),
		5792 => to_signed(17275, LUT_AMPL_WIDTH),
		5793 => to_signed(17277, LUT_AMPL_WIDTH),
		5794 => to_signed(17280, LUT_AMPL_WIDTH),
		5795 => to_signed(17283, LUT_AMPL_WIDTH),
		5796 => to_signed(17285, LUT_AMPL_WIDTH),
		5797 => to_signed(17288, LUT_AMPL_WIDTH),
		5798 => to_signed(17291, LUT_AMPL_WIDTH),
		5799 => to_signed(17293, LUT_AMPL_WIDTH),
		5800 => to_signed(17296, LUT_AMPL_WIDTH),
		5801 => to_signed(17299, LUT_AMPL_WIDTH),
		5802 => to_signed(17301, LUT_AMPL_WIDTH),
		5803 => to_signed(17304, LUT_AMPL_WIDTH),
		5804 => to_signed(17307, LUT_AMPL_WIDTH),
		5805 => to_signed(17309, LUT_AMPL_WIDTH),
		5806 => to_signed(17312, LUT_AMPL_WIDTH),
		5807 => to_signed(17315, LUT_AMPL_WIDTH),
		5808 => to_signed(17317, LUT_AMPL_WIDTH),
		5809 => to_signed(17320, LUT_AMPL_WIDTH),
		5810 => to_signed(17323, LUT_AMPL_WIDTH),
		5811 => to_signed(17325, LUT_AMPL_WIDTH),
		5812 => to_signed(17328, LUT_AMPL_WIDTH),
		5813 => to_signed(17331, LUT_AMPL_WIDTH),
		5814 => to_signed(17333, LUT_AMPL_WIDTH),
		5815 => to_signed(17336, LUT_AMPL_WIDTH),
		5816 => to_signed(17339, LUT_AMPL_WIDTH),
		5817 => to_signed(17341, LUT_AMPL_WIDTH),
		5818 => to_signed(17344, LUT_AMPL_WIDTH),
		5819 => to_signed(17347, LUT_AMPL_WIDTH),
		5820 => to_signed(17349, LUT_AMPL_WIDTH),
		5821 => to_signed(17352, LUT_AMPL_WIDTH),
		5822 => to_signed(17355, LUT_AMPL_WIDTH),
		5823 => to_signed(17357, LUT_AMPL_WIDTH),
		5824 => to_signed(17360, LUT_AMPL_WIDTH),
		5825 => to_signed(17363, LUT_AMPL_WIDTH),
		5826 => to_signed(17365, LUT_AMPL_WIDTH),
		5827 => to_signed(17368, LUT_AMPL_WIDTH),
		5828 => to_signed(17371, LUT_AMPL_WIDTH),
		5829 => to_signed(17373, LUT_AMPL_WIDTH),
		5830 => to_signed(17376, LUT_AMPL_WIDTH),
		5831 => to_signed(17379, LUT_AMPL_WIDTH),
		5832 => to_signed(17381, LUT_AMPL_WIDTH),
		5833 => to_signed(17384, LUT_AMPL_WIDTH),
		5834 => to_signed(17387, LUT_AMPL_WIDTH),
		5835 => to_signed(17389, LUT_AMPL_WIDTH),
		5836 => to_signed(17392, LUT_AMPL_WIDTH),
		5837 => to_signed(17395, LUT_AMPL_WIDTH),
		5838 => to_signed(17397, LUT_AMPL_WIDTH),
		5839 => to_signed(17400, LUT_AMPL_WIDTH),
		5840 => to_signed(17403, LUT_AMPL_WIDTH),
		5841 => to_signed(17405, LUT_AMPL_WIDTH),
		5842 => to_signed(17408, LUT_AMPL_WIDTH),
		5843 => to_signed(17411, LUT_AMPL_WIDTH),
		5844 => to_signed(17413, LUT_AMPL_WIDTH),
		5845 => to_signed(17416, LUT_AMPL_WIDTH),
		5846 => to_signed(17419, LUT_AMPL_WIDTH),
		5847 => to_signed(17421, LUT_AMPL_WIDTH),
		5848 => to_signed(17424, LUT_AMPL_WIDTH),
		5849 => to_signed(17427, LUT_AMPL_WIDTH),
		5850 => to_signed(17429, LUT_AMPL_WIDTH),
		5851 => to_signed(17432, LUT_AMPL_WIDTH),
		5852 => to_signed(17435, LUT_AMPL_WIDTH),
		5853 => to_signed(17437, LUT_AMPL_WIDTH),
		5854 => to_signed(17440, LUT_AMPL_WIDTH),
		5855 => to_signed(17443, LUT_AMPL_WIDTH),
		5856 => to_signed(17445, LUT_AMPL_WIDTH),
		5857 => to_signed(17448, LUT_AMPL_WIDTH),
		5858 => to_signed(17451, LUT_AMPL_WIDTH),
		5859 => to_signed(17453, LUT_AMPL_WIDTH),
		5860 => to_signed(17456, LUT_AMPL_WIDTH),
		5861 => to_signed(17459, LUT_AMPL_WIDTH),
		5862 => to_signed(17461, LUT_AMPL_WIDTH),
		5863 => to_signed(17464, LUT_AMPL_WIDTH),
		5864 => to_signed(17467, LUT_AMPL_WIDTH),
		5865 => to_signed(17469, LUT_AMPL_WIDTH),
		5866 => to_signed(17472, LUT_AMPL_WIDTH),
		5867 => to_signed(17474, LUT_AMPL_WIDTH),
		5868 => to_signed(17477, LUT_AMPL_WIDTH),
		5869 => to_signed(17480, LUT_AMPL_WIDTH),
		5870 => to_signed(17482, LUT_AMPL_WIDTH),
		5871 => to_signed(17485, LUT_AMPL_WIDTH),
		5872 => to_signed(17488, LUT_AMPL_WIDTH),
		5873 => to_signed(17490, LUT_AMPL_WIDTH),
		5874 => to_signed(17493, LUT_AMPL_WIDTH),
		5875 => to_signed(17496, LUT_AMPL_WIDTH),
		5876 => to_signed(17498, LUT_AMPL_WIDTH),
		5877 => to_signed(17501, LUT_AMPL_WIDTH),
		5878 => to_signed(17504, LUT_AMPL_WIDTH),
		5879 => to_signed(17506, LUT_AMPL_WIDTH),
		5880 => to_signed(17509, LUT_AMPL_WIDTH),
		5881 => to_signed(17512, LUT_AMPL_WIDTH),
		5882 => to_signed(17514, LUT_AMPL_WIDTH),
		5883 => to_signed(17517, LUT_AMPL_WIDTH),
		5884 => to_signed(17520, LUT_AMPL_WIDTH),
		5885 => to_signed(17522, LUT_AMPL_WIDTH),
		5886 => to_signed(17525, LUT_AMPL_WIDTH),
		5887 => to_signed(17528, LUT_AMPL_WIDTH),
		5888 => to_signed(17530, LUT_AMPL_WIDTH),
		5889 => to_signed(17533, LUT_AMPL_WIDTH),
		5890 => to_signed(17536, LUT_AMPL_WIDTH),
		5891 => to_signed(17538, LUT_AMPL_WIDTH),
		5892 => to_signed(17541, LUT_AMPL_WIDTH),
		5893 => to_signed(17544, LUT_AMPL_WIDTH),
		5894 => to_signed(17546, LUT_AMPL_WIDTH),
		5895 => to_signed(17549, LUT_AMPL_WIDTH),
		5896 => to_signed(17551, LUT_AMPL_WIDTH),
		5897 => to_signed(17554, LUT_AMPL_WIDTH),
		5898 => to_signed(17557, LUT_AMPL_WIDTH),
		5899 => to_signed(17559, LUT_AMPL_WIDTH),
		5900 => to_signed(17562, LUT_AMPL_WIDTH),
		5901 => to_signed(17565, LUT_AMPL_WIDTH),
		5902 => to_signed(17567, LUT_AMPL_WIDTH),
		5903 => to_signed(17570, LUT_AMPL_WIDTH),
		5904 => to_signed(17573, LUT_AMPL_WIDTH),
		5905 => to_signed(17575, LUT_AMPL_WIDTH),
		5906 => to_signed(17578, LUT_AMPL_WIDTH),
		5907 => to_signed(17581, LUT_AMPL_WIDTH),
		5908 => to_signed(17583, LUT_AMPL_WIDTH),
		5909 => to_signed(17586, LUT_AMPL_WIDTH),
		5910 => to_signed(17589, LUT_AMPL_WIDTH),
		5911 => to_signed(17591, LUT_AMPL_WIDTH),
		5912 => to_signed(17594, LUT_AMPL_WIDTH),
		5913 => to_signed(17597, LUT_AMPL_WIDTH),
		5914 => to_signed(17599, LUT_AMPL_WIDTH),
		5915 => to_signed(17602, LUT_AMPL_WIDTH),
		5916 => to_signed(17605, LUT_AMPL_WIDTH),
		5917 => to_signed(17607, LUT_AMPL_WIDTH),
		5918 => to_signed(17610, LUT_AMPL_WIDTH),
		5919 => to_signed(17612, LUT_AMPL_WIDTH),
		5920 => to_signed(17615, LUT_AMPL_WIDTH),
		5921 => to_signed(17618, LUT_AMPL_WIDTH),
		5922 => to_signed(17620, LUT_AMPL_WIDTH),
		5923 => to_signed(17623, LUT_AMPL_WIDTH),
		5924 => to_signed(17626, LUT_AMPL_WIDTH),
		5925 => to_signed(17628, LUT_AMPL_WIDTH),
		5926 => to_signed(17631, LUT_AMPL_WIDTH),
		5927 => to_signed(17634, LUT_AMPL_WIDTH),
		5928 => to_signed(17636, LUT_AMPL_WIDTH),
		5929 => to_signed(17639, LUT_AMPL_WIDTH),
		5930 => to_signed(17642, LUT_AMPL_WIDTH),
		5931 => to_signed(17644, LUT_AMPL_WIDTH),
		5932 => to_signed(17647, LUT_AMPL_WIDTH),
		5933 => to_signed(17650, LUT_AMPL_WIDTH),
		5934 => to_signed(17652, LUT_AMPL_WIDTH),
		5935 => to_signed(17655, LUT_AMPL_WIDTH),
		5936 => to_signed(17657, LUT_AMPL_WIDTH),
		5937 => to_signed(17660, LUT_AMPL_WIDTH),
		5938 => to_signed(17663, LUT_AMPL_WIDTH),
		5939 => to_signed(17665, LUT_AMPL_WIDTH),
		5940 => to_signed(17668, LUT_AMPL_WIDTH),
		5941 => to_signed(17671, LUT_AMPL_WIDTH),
		5942 => to_signed(17673, LUT_AMPL_WIDTH),
		5943 => to_signed(17676, LUT_AMPL_WIDTH),
		5944 => to_signed(17679, LUT_AMPL_WIDTH),
		5945 => to_signed(17681, LUT_AMPL_WIDTH),
		5946 => to_signed(17684, LUT_AMPL_WIDTH),
		5947 => to_signed(17687, LUT_AMPL_WIDTH),
		5948 => to_signed(17689, LUT_AMPL_WIDTH),
		5949 => to_signed(17692, LUT_AMPL_WIDTH),
		5950 => to_signed(17695, LUT_AMPL_WIDTH),
		5951 => to_signed(17697, LUT_AMPL_WIDTH),
		5952 => to_signed(17700, LUT_AMPL_WIDTH),
		5953 => to_signed(17702, LUT_AMPL_WIDTH),
		5954 => to_signed(17705, LUT_AMPL_WIDTH),
		5955 => to_signed(17708, LUT_AMPL_WIDTH),
		5956 => to_signed(17710, LUT_AMPL_WIDTH),
		5957 => to_signed(17713, LUT_AMPL_WIDTH),
		5958 => to_signed(17716, LUT_AMPL_WIDTH),
		5959 => to_signed(17718, LUT_AMPL_WIDTH),
		5960 => to_signed(17721, LUT_AMPL_WIDTH),
		5961 => to_signed(17724, LUT_AMPL_WIDTH),
		5962 => to_signed(17726, LUT_AMPL_WIDTH),
		5963 => to_signed(17729, LUT_AMPL_WIDTH),
		5964 => to_signed(17732, LUT_AMPL_WIDTH),
		5965 => to_signed(17734, LUT_AMPL_WIDTH),
		5966 => to_signed(17737, LUT_AMPL_WIDTH),
		5967 => to_signed(17739, LUT_AMPL_WIDTH),
		5968 => to_signed(17742, LUT_AMPL_WIDTH),
		5969 => to_signed(17745, LUT_AMPL_WIDTH),
		5970 => to_signed(17747, LUT_AMPL_WIDTH),
		5971 => to_signed(17750, LUT_AMPL_WIDTH),
		5972 => to_signed(17753, LUT_AMPL_WIDTH),
		5973 => to_signed(17755, LUT_AMPL_WIDTH),
		5974 => to_signed(17758, LUT_AMPL_WIDTH),
		5975 => to_signed(17761, LUT_AMPL_WIDTH),
		5976 => to_signed(17763, LUT_AMPL_WIDTH),
		5977 => to_signed(17766, LUT_AMPL_WIDTH),
		5978 => to_signed(17768, LUT_AMPL_WIDTH),
		5979 => to_signed(17771, LUT_AMPL_WIDTH),
		5980 => to_signed(17774, LUT_AMPL_WIDTH),
		5981 => to_signed(17776, LUT_AMPL_WIDTH),
		5982 => to_signed(17779, LUT_AMPL_WIDTH),
		5983 => to_signed(17782, LUT_AMPL_WIDTH),
		5984 => to_signed(17784, LUT_AMPL_WIDTH),
		5985 => to_signed(17787, LUT_AMPL_WIDTH),
		5986 => to_signed(17790, LUT_AMPL_WIDTH),
		5987 => to_signed(17792, LUT_AMPL_WIDTH),
		5988 => to_signed(17795, LUT_AMPL_WIDTH),
		5989 => to_signed(17798, LUT_AMPL_WIDTH),
		5990 => to_signed(17800, LUT_AMPL_WIDTH),
		5991 => to_signed(17803, LUT_AMPL_WIDTH),
		5992 => to_signed(17805, LUT_AMPL_WIDTH),
		5993 => to_signed(17808, LUT_AMPL_WIDTH),
		5994 => to_signed(17811, LUT_AMPL_WIDTH),
		5995 => to_signed(17813, LUT_AMPL_WIDTH),
		5996 => to_signed(17816, LUT_AMPL_WIDTH),
		5997 => to_signed(17819, LUT_AMPL_WIDTH),
		5998 => to_signed(17821, LUT_AMPL_WIDTH),
		5999 => to_signed(17824, LUT_AMPL_WIDTH),
		6000 => to_signed(17827, LUT_AMPL_WIDTH),
		6001 => to_signed(17829, LUT_AMPL_WIDTH),
		6002 => to_signed(17832, LUT_AMPL_WIDTH),
		6003 => to_signed(17834, LUT_AMPL_WIDTH),
		6004 => to_signed(17837, LUT_AMPL_WIDTH),
		6005 => to_signed(17840, LUT_AMPL_WIDTH),
		6006 => to_signed(17842, LUT_AMPL_WIDTH),
		6007 => to_signed(17845, LUT_AMPL_WIDTH),
		6008 => to_signed(17848, LUT_AMPL_WIDTH),
		6009 => to_signed(17850, LUT_AMPL_WIDTH),
		6010 => to_signed(17853, LUT_AMPL_WIDTH),
		6011 => to_signed(17855, LUT_AMPL_WIDTH),
		6012 => to_signed(17858, LUT_AMPL_WIDTH),
		6013 => to_signed(17861, LUT_AMPL_WIDTH),
		6014 => to_signed(17863, LUT_AMPL_WIDTH),
		6015 => to_signed(17866, LUT_AMPL_WIDTH),
		6016 => to_signed(17869, LUT_AMPL_WIDTH),
		6017 => to_signed(17871, LUT_AMPL_WIDTH),
		6018 => to_signed(17874, LUT_AMPL_WIDTH),
		6019 => to_signed(17877, LUT_AMPL_WIDTH),
		6020 => to_signed(17879, LUT_AMPL_WIDTH),
		6021 => to_signed(17882, LUT_AMPL_WIDTH),
		6022 => to_signed(17884, LUT_AMPL_WIDTH),
		6023 => to_signed(17887, LUT_AMPL_WIDTH),
		6024 => to_signed(17890, LUT_AMPL_WIDTH),
		6025 => to_signed(17892, LUT_AMPL_WIDTH),
		6026 => to_signed(17895, LUT_AMPL_WIDTH),
		6027 => to_signed(17898, LUT_AMPL_WIDTH),
		6028 => to_signed(17900, LUT_AMPL_WIDTH),
		6029 => to_signed(17903, LUT_AMPL_WIDTH),
		6030 => to_signed(17906, LUT_AMPL_WIDTH),
		6031 => to_signed(17908, LUT_AMPL_WIDTH),
		6032 => to_signed(17911, LUT_AMPL_WIDTH),
		6033 => to_signed(17913, LUT_AMPL_WIDTH),
		6034 => to_signed(17916, LUT_AMPL_WIDTH),
		6035 => to_signed(17919, LUT_AMPL_WIDTH),
		6036 => to_signed(17921, LUT_AMPL_WIDTH),
		6037 => to_signed(17924, LUT_AMPL_WIDTH),
		6038 => to_signed(17927, LUT_AMPL_WIDTH),
		6039 => to_signed(17929, LUT_AMPL_WIDTH),
		6040 => to_signed(17932, LUT_AMPL_WIDTH),
		6041 => to_signed(17934, LUT_AMPL_WIDTH),
		6042 => to_signed(17937, LUT_AMPL_WIDTH),
		6043 => to_signed(17940, LUT_AMPL_WIDTH),
		6044 => to_signed(17942, LUT_AMPL_WIDTH),
		6045 => to_signed(17945, LUT_AMPL_WIDTH),
		6046 => to_signed(17948, LUT_AMPL_WIDTH),
		6047 => to_signed(17950, LUT_AMPL_WIDTH),
		6048 => to_signed(17953, LUT_AMPL_WIDTH),
		6049 => to_signed(17955, LUT_AMPL_WIDTH),
		6050 => to_signed(17958, LUT_AMPL_WIDTH),
		6051 => to_signed(17961, LUT_AMPL_WIDTH),
		6052 => to_signed(17963, LUT_AMPL_WIDTH),
		6053 => to_signed(17966, LUT_AMPL_WIDTH),
		6054 => to_signed(17969, LUT_AMPL_WIDTH),
		6055 => to_signed(17971, LUT_AMPL_WIDTH),
		6056 => to_signed(17974, LUT_AMPL_WIDTH),
		6057 => to_signed(17976, LUT_AMPL_WIDTH),
		6058 => to_signed(17979, LUT_AMPL_WIDTH),
		6059 => to_signed(17982, LUT_AMPL_WIDTH),
		6060 => to_signed(17984, LUT_AMPL_WIDTH),
		6061 => to_signed(17987, LUT_AMPL_WIDTH),
		6062 => to_signed(17990, LUT_AMPL_WIDTH),
		6063 => to_signed(17992, LUT_AMPL_WIDTH),
		6064 => to_signed(17995, LUT_AMPL_WIDTH),
		6065 => to_signed(17997, LUT_AMPL_WIDTH),
		6066 => to_signed(18000, LUT_AMPL_WIDTH),
		6067 => to_signed(18003, LUT_AMPL_WIDTH),
		6068 => to_signed(18005, LUT_AMPL_WIDTH),
		6069 => to_signed(18008, LUT_AMPL_WIDTH),
		6070 => to_signed(18011, LUT_AMPL_WIDTH),
		6071 => to_signed(18013, LUT_AMPL_WIDTH),
		6072 => to_signed(18016, LUT_AMPL_WIDTH),
		6073 => to_signed(18018, LUT_AMPL_WIDTH),
		6074 => to_signed(18021, LUT_AMPL_WIDTH),
		6075 => to_signed(18024, LUT_AMPL_WIDTH),
		6076 => to_signed(18026, LUT_AMPL_WIDTH),
		6077 => to_signed(18029, LUT_AMPL_WIDTH),
		6078 => to_signed(18032, LUT_AMPL_WIDTH),
		6079 => to_signed(18034, LUT_AMPL_WIDTH),
		6080 => to_signed(18037, LUT_AMPL_WIDTH),
		6081 => to_signed(18039, LUT_AMPL_WIDTH),
		6082 => to_signed(18042, LUT_AMPL_WIDTH),
		6083 => to_signed(18045, LUT_AMPL_WIDTH),
		6084 => to_signed(18047, LUT_AMPL_WIDTH),
		6085 => to_signed(18050, LUT_AMPL_WIDTH),
		6086 => to_signed(18053, LUT_AMPL_WIDTH),
		6087 => to_signed(18055, LUT_AMPL_WIDTH),
		6088 => to_signed(18058, LUT_AMPL_WIDTH),
		6089 => to_signed(18060, LUT_AMPL_WIDTH),
		6090 => to_signed(18063, LUT_AMPL_WIDTH),
		6091 => to_signed(18066, LUT_AMPL_WIDTH),
		6092 => to_signed(18068, LUT_AMPL_WIDTH),
		6093 => to_signed(18071, LUT_AMPL_WIDTH),
		6094 => to_signed(18074, LUT_AMPL_WIDTH),
		6095 => to_signed(18076, LUT_AMPL_WIDTH),
		6096 => to_signed(18079, LUT_AMPL_WIDTH),
		6097 => to_signed(18081, LUT_AMPL_WIDTH),
		6098 => to_signed(18084, LUT_AMPL_WIDTH),
		6099 => to_signed(18087, LUT_AMPL_WIDTH),
		6100 => to_signed(18089, LUT_AMPL_WIDTH),
		6101 => to_signed(18092, LUT_AMPL_WIDTH),
		6102 => to_signed(18095, LUT_AMPL_WIDTH),
		6103 => to_signed(18097, LUT_AMPL_WIDTH),
		6104 => to_signed(18100, LUT_AMPL_WIDTH),
		6105 => to_signed(18102, LUT_AMPL_WIDTH),
		6106 => to_signed(18105, LUT_AMPL_WIDTH),
		6107 => to_signed(18108, LUT_AMPL_WIDTH),
		6108 => to_signed(18110, LUT_AMPL_WIDTH),
		6109 => to_signed(18113, LUT_AMPL_WIDTH),
		6110 => to_signed(18115, LUT_AMPL_WIDTH),
		6111 => to_signed(18118, LUT_AMPL_WIDTH),
		6112 => to_signed(18121, LUT_AMPL_WIDTH),
		6113 => to_signed(18123, LUT_AMPL_WIDTH),
		6114 => to_signed(18126, LUT_AMPL_WIDTH),
		6115 => to_signed(18129, LUT_AMPL_WIDTH),
		6116 => to_signed(18131, LUT_AMPL_WIDTH),
		6117 => to_signed(18134, LUT_AMPL_WIDTH),
		6118 => to_signed(18136, LUT_AMPL_WIDTH),
		6119 => to_signed(18139, LUT_AMPL_WIDTH),
		6120 => to_signed(18142, LUT_AMPL_WIDTH),
		6121 => to_signed(18144, LUT_AMPL_WIDTH),
		6122 => to_signed(18147, LUT_AMPL_WIDTH),
		6123 => to_signed(18149, LUT_AMPL_WIDTH),
		6124 => to_signed(18152, LUT_AMPL_WIDTH),
		6125 => to_signed(18155, LUT_AMPL_WIDTH),
		6126 => to_signed(18157, LUT_AMPL_WIDTH),
		6127 => to_signed(18160, LUT_AMPL_WIDTH),
		6128 => to_signed(18163, LUT_AMPL_WIDTH),
		6129 => to_signed(18165, LUT_AMPL_WIDTH),
		6130 => to_signed(18168, LUT_AMPL_WIDTH),
		6131 => to_signed(18170, LUT_AMPL_WIDTH),
		6132 => to_signed(18173, LUT_AMPL_WIDTH),
		6133 => to_signed(18176, LUT_AMPL_WIDTH),
		6134 => to_signed(18178, LUT_AMPL_WIDTH),
		6135 => to_signed(18181, LUT_AMPL_WIDTH),
		6136 => to_signed(18183, LUT_AMPL_WIDTH),
		6137 => to_signed(18186, LUT_AMPL_WIDTH),
		6138 => to_signed(18189, LUT_AMPL_WIDTH),
		6139 => to_signed(18191, LUT_AMPL_WIDTH),
		6140 => to_signed(18194, LUT_AMPL_WIDTH),
		6141 => to_signed(18197, LUT_AMPL_WIDTH),
		6142 => to_signed(18199, LUT_AMPL_WIDTH),
		6143 => to_signed(18202, LUT_AMPL_WIDTH),
		6144 => to_signed(18204, LUT_AMPL_WIDTH),
		6145 => to_signed(18207, LUT_AMPL_WIDTH),
		6146 => to_signed(18210, LUT_AMPL_WIDTH),
		6147 => to_signed(18212, LUT_AMPL_WIDTH),
		6148 => to_signed(18215, LUT_AMPL_WIDTH),
		6149 => to_signed(18217, LUT_AMPL_WIDTH),
		6150 => to_signed(18220, LUT_AMPL_WIDTH),
		6151 => to_signed(18223, LUT_AMPL_WIDTH),
		6152 => to_signed(18225, LUT_AMPL_WIDTH),
		6153 => to_signed(18228, LUT_AMPL_WIDTH),
		6154 => to_signed(18230, LUT_AMPL_WIDTH),
		6155 => to_signed(18233, LUT_AMPL_WIDTH),
		6156 => to_signed(18236, LUT_AMPL_WIDTH),
		6157 => to_signed(18238, LUT_AMPL_WIDTH),
		6158 => to_signed(18241, LUT_AMPL_WIDTH),
		6159 => to_signed(18244, LUT_AMPL_WIDTH),
		6160 => to_signed(18246, LUT_AMPL_WIDTH),
		6161 => to_signed(18249, LUT_AMPL_WIDTH),
		6162 => to_signed(18251, LUT_AMPL_WIDTH),
		6163 => to_signed(18254, LUT_AMPL_WIDTH),
		6164 => to_signed(18257, LUT_AMPL_WIDTH),
		6165 => to_signed(18259, LUT_AMPL_WIDTH),
		6166 => to_signed(18262, LUT_AMPL_WIDTH),
		6167 => to_signed(18264, LUT_AMPL_WIDTH),
		6168 => to_signed(18267, LUT_AMPL_WIDTH),
		6169 => to_signed(18270, LUT_AMPL_WIDTH),
		6170 => to_signed(18272, LUT_AMPL_WIDTH),
		6171 => to_signed(18275, LUT_AMPL_WIDTH),
		6172 => to_signed(18277, LUT_AMPL_WIDTH),
		6173 => to_signed(18280, LUT_AMPL_WIDTH),
		6174 => to_signed(18283, LUT_AMPL_WIDTH),
		6175 => to_signed(18285, LUT_AMPL_WIDTH),
		6176 => to_signed(18288, LUT_AMPL_WIDTH),
		6177 => to_signed(18290, LUT_AMPL_WIDTH),
		6178 => to_signed(18293, LUT_AMPL_WIDTH),
		6179 => to_signed(18296, LUT_AMPL_WIDTH),
		6180 => to_signed(18298, LUT_AMPL_WIDTH),
		6181 => to_signed(18301, LUT_AMPL_WIDTH),
		6182 => to_signed(18304, LUT_AMPL_WIDTH),
		6183 => to_signed(18306, LUT_AMPL_WIDTH),
		6184 => to_signed(18309, LUT_AMPL_WIDTH),
		6185 => to_signed(18311, LUT_AMPL_WIDTH),
		6186 => to_signed(18314, LUT_AMPL_WIDTH),
		6187 => to_signed(18317, LUT_AMPL_WIDTH),
		6188 => to_signed(18319, LUT_AMPL_WIDTH),
		6189 => to_signed(18322, LUT_AMPL_WIDTH),
		6190 => to_signed(18324, LUT_AMPL_WIDTH),
		6191 => to_signed(18327, LUT_AMPL_WIDTH),
		6192 => to_signed(18330, LUT_AMPL_WIDTH),
		6193 => to_signed(18332, LUT_AMPL_WIDTH),
		6194 => to_signed(18335, LUT_AMPL_WIDTH),
		6195 => to_signed(18337, LUT_AMPL_WIDTH),
		6196 => to_signed(18340, LUT_AMPL_WIDTH),
		6197 => to_signed(18343, LUT_AMPL_WIDTH),
		6198 => to_signed(18345, LUT_AMPL_WIDTH),
		6199 => to_signed(18348, LUT_AMPL_WIDTH),
		6200 => to_signed(18350, LUT_AMPL_WIDTH),
		6201 => to_signed(18353, LUT_AMPL_WIDTH),
		6202 => to_signed(18356, LUT_AMPL_WIDTH),
		6203 => to_signed(18358, LUT_AMPL_WIDTH),
		6204 => to_signed(18361, LUT_AMPL_WIDTH),
		6205 => to_signed(18363, LUT_AMPL_WIDTH),
		6206 => to_signed(18366, LUT_AMPL_WIDTH),
		6207 => to_signed(18369, LUT_AMPL_WIDTH),
		6208 => to_signed(18371, LUT_AMPL_WIDTH),
		6209 => to_signed(18374, LUT_AMPL_WIDTH),
		6210 => to_signed(18376, LUT_AMPL_WIDTH),
		6211 => to_signed(18379, LUT_AMPL_WIDTH),
		6212 => to_signed(18382, LUT_AMPL_WIDTH),
		6213 => to_signed(18384, LUT_AMPL_WIDTH),
		6214 => to_signed(18387, LUT_AMPL_WIDTH),
		6215 => to_signed(18389, LUT_AMPL_WIDTH),
		6216 => to_signed(18392, LUT_AMPL_WIDTH),
		6217 => to_signed(18395, LUT_AMPL_WIDTH),
		6218 => to_signed(18397, LUT_AMPL_WIDTH),
		6219 => to_signed(18400, LUT_AMPL_WIDTH),
		6220 => to_signed(18402, LUT_AMPL_WIDTH),
		6221 => to_signed(18405, LUT_AMPL_WIDTH),
		6222 => to_signed(18408, LUT_AMPL_WIDTH),
		6223 => to_signed(18410, LUT_AMPL_WIDTH),
		6224 => to_signed(18413, LUT_AMPL_WIDTH),
		6225 => to_signed(18415, LUT_AMPL_WIDTH),
		6226 => to_signed(18418, LUT_AMPL_WIDTH),
		6227 => to_signed(18421, LUT_AMPL_WIDTH),
		6228 => to_signed(18423, LUT_AMPL_WIDTH),
		6229 => to_signed(18426, LUT_AMPL_WIDTH),
		6230 => to_signed(18428, LUT_AMPL_WIDTH),
		6231 => to_signed(18431, LUT_AMPL_WIDTH),
		6232 => to_signed(18434, LUT_AMPL_WIDTH),
		6233 => to_signed(18436, LUT_AMPL_WIDTH),
		6234 => to_signed(18439, LUT_AMPL_WIDTH),
		6235 => to_signed(18441, LUT_AMPL_WIDTH),
		6236 => to_signed(18444, LUT_AMPL_WIDTH),
		6237 => to_signed(18447, LUT_AMPL_WIDTH),
		6238 => to_signed(18449, LUT_AMPL_WIDTH),
		6239 => to_signed(18452, LUT_AMPL_WIDTH),
		6240 => to_signed(18454, LUT_AMPL_WIDTH),
		6241 => to_signed(18457, LUT_AMPL_WIDTH),
		6242 => to_signed(18460, LUT_AMPL_WIDTH),
		6243 => to_signed(18462, LUT_AMPL_WIDTH),
		6244 => to_signed(18465, LUT_AMPL_WIDTH),
		6245 => to_signed(18467, LUT_AMPL_WIDTH),
		6246 => to_signed(18470, LUT_AMPL_WIDTH),
		6247 => to_signed(18473, LUT_AMPL_WIDTH),
		6248 => to_signed(18475, LUT_AMPL_WIDTH),
		6249 => to_signed(18478, LUT_AMPL_WIDTH),
		6250 => to_signed(18480, LUT_AMPL_WIDTH),
		6251 => to_signed(18483, LUT_AMPL_WIDTH),
		6252 => to_signed(18485, LUT_AMPL_WIDTH),
		6253 => to_signed(18488, LUT_AMPL_WIDTH),
		6254 => to_signed(18491, LUT_AMPL_WIDTH),
		6255 => to_signed(18493, LUT_AMPL_WIDTH),
		6256 => to_signed(18496, LUT_AMPL_WIDTH),
		6257 => to_signed(18498, LUT_AMPL_WIDTH),
		6258 => to_signed(18501, LUT_AMPL_WIDTH),
		6259 => to_signed(18504, LUT_AMPL_WIDTH),
		6260 => to_signed(18506, LUT_AMPL_WIDTH),
		6261 => to_signed(18509, LUT_AMPL_WIDTH),
		6262 => to_signed(18511, LUT_AMPL_WIDTH),
		6263 => to_signed(18514, LUT_AMPL_WIDTH),
		6264 => to_signed(18517, LUT_AMPL_WIDTH),
		6265 => to_signed(18519, LUT_AMPL_WIDTH),
		6266 => to_signed(18522, LUT_AMPL_WIDTH),
		6267 => to_signed(18524, LUT_AMPL_WIDTH),
		6268 => to_signed(18527, LUT_AMPL_WIDTH),
		6269 => to_signed(18530, LUT_AMPL_WIDTH),
		6270 => to_signed(18532, LUT_AMPL_WIDTH),
		6271 => to_signed(18535, LUT_AMPL_WIDTH),
		6272 => to_signed(18537, LUT_AMPL_WIDTH),
		6273 => to_signed(18540, LUT_AMPL_WIDTH),
		6274 => to_signed(18543, LUT_AMPL_WIDTH),
		6275 => to_signed(18545, LUT_AMPL_WIDTH),
		6276 => to_signed(18548, LUT_AMPL_WIDTH),
		6277 => to_signed(18550, LUT_AMPL_WIDTH),
		6278 => to_signed(18553, LUT_AMPL_WIDTH),
		6279 => to_signed(18555, LUT_AMPL_WIDTH),
		6280 => to_signed(18558, LUT_AMPL_WIDTH),
		6281 => to_signed(18561, LUT_AMPL_WIDTH),
		6282 => to_signed(18563, LUT_AMPL_WIDTH),
		6283 => to_signed(18566, LUT_AMPL_WIDTH),
		6284 => to_signed(18568, LUT_AMPL_WIDTH),
		6285 => to_signed(18571, LUT_AMPL_WIDTH),
		6286 => to_signed(18574, LUT_AMPL_WIDTH),
		6287 => to_signed(18576, LUT_AMPL_WIDTH),
		6288 => to_signed(18579, LUT_AMPL_WIDTH),
		6289 => to_signed(18581, LUT_AMPL_WIDTH),
		6290 => to_signed(18584, LUT_AMPL_WIDTH),
		6291 => to_signed(18587, LUT_AMPL_WIDTH),
		6292 => to_signed(18589, LUT_AMPL_WIDTH),
		6293 => to_signed(18592, LUT_AMPL_WIDTH),
		6294 => to_signed(18594, LUT_AMPL_WIDTH),
		6295 => to_signed(18597, LUT_AMPL_WIDTH),
		6296 => to_signed(18599, LUT_AMPL_WIDTH),
		6297 => to_signed(18602, LUT_AMPL_WIDTH),
		6298 => to_signed(18605, LUT_AMPL_WIDTH),
		6299 => to_signed(18607, LUT_AMPL_WIDTH),
		6300 => to_signed(18610, LUT_AMPL_WIDTH),
		6301 => to_signed(18612, LUT_AMPL_WIDTH),
		6302 => to_signed(18615, LUT_AMPL_WIDTH),
		6303 => to_signed(18618, LUT_AMPL_WIDTH),
		6304 => to_signed(18620, LUT_AMPL_WIDTH),
		6305 => to_signed(18623, LUT_AMPL_WIDTH),
		6306 => to_signed(18625, LUT_AMPL_WIDTH),
		6307 => to_signed(18628, LUT_AMPL_WIDTH),
		6308 => to_signed(18630, LUT_AMPL_WIDTH),
		6309 => to_signed(18633, LUT_AMPL_WIDTH),
		6310 => to_signed(18636, LUT_AMPL_WIDTH),
		6311 => to_signed(18638, LUT_AMPL_WIDTH),
		6312 => to_signed(18641, LUT_AMPL_WIDTH),
		6313 => to_signed(18643, LUT_AMPL_WIDTH),
		6314 => to_signed(18646, LUT_AMPL_WIDTH),
		6315 => to_signed(18649, LUT_AMPL_WIDTH),
		6316 => to_signed(18651, LUT_AMPL_WIDTH),
		6317 => to_signed(18654, LUT_AMPL_WIDTH),
		6318 => to_signed(18656, LUT_AMPL_WIDTH),
		6319 => to_signed(18659, LUT_AMPL_WIDTH),
		6320 => to_signed(18661, LUT_AMPL_WIDTH),
		6321 => to_signed(18664, LUT_AMPL_WIDTH),
		6322 => to_signed(18667, LUT_AMPL_WIDTH),
		6323 => to_signed(18669, LUT_AMPL_WIDTH),
		6324 => to_signed(18672, LUT_AMPL_WIDTH),
		6325 => to_signed(18674, LUT_AMPL_WIDTH),
		6326 => to_signed(18677, LUT_AMPL_WIDTH),
		6327 => to_signed(18680, LUT_AMPL_WIDTH),
		6328 => to_signed(18682, LUT_AMPL_WIDTH),
		6329 => to_signed(18685, LUT_AMPL_WIDTH),
		6330 => to_signed(18687, LUT_AMPL_WIDTH),
		6331 => to_signed(18690, LUT_AMPL_WIDTH),
		6332 => to_signed(18692, LUT_AMPL_WIDTH),
		6333 => to_signed(18695, LUT_AMPL_WIDTH),
		6334 => to_signed(18698, LUT_AMPL_WIDTH),
		6335 => to_signed(18700, LUT_AMPL_WIDTH),
		6336 => to_signed(18703, LUT_AMPL_WIDTH),
		6337 => to_signed(18705, LUT_AMPL_WIDTH),
		6338 => to_signed(18708, LUT_AMPL_WIDTH),
		6339 => to_signed(18711, LUT_AMPL_WIDTH),
		6340 => to_signed(18713, LUT_AMPL_WIDTH),
		6341 => to_signed(18716, LUT_AMPL_WIDTH),
		6342 => to_signed(18718, LUT_AMPL_WIDTH),
		6343 => to_signed(18721, LUT_AMPL_WIDTH),
		6344 => to_signed(18723, LUT_AMPL_WIDTH),
		6345 => to_signed(18726, LUT_AMPL_WIDTH),
		6346 => to_signed(18729, LUT_AMPL_WIDTH),
		6347 => to_signed(18731, LUT_AMPL_WIDTH),
		6348 => to_signed(18734, LUT_AMPL_WIDTH),
		6349 => to_signed(18736, LUT_AMPL_WIDTH),
		6350 => to_signed(18739, LUT_AMPL_WIDTH),
		6351 => to_signed(18741, LUT_AMPL_WIDTH),
		6352 => to_signed(18744, LUT_AMPL_WIDTH),
		6353 => to_signed(18747, LUT_AMPL_WIDTH),
		6354 => to_signed(18749, LUT_AMPL_WIDTH),
		6355 => to_signed(18752, LUT_AMPL_WIDTH),
		6356 => to_signed(18754, LUT_AMPL_WIDTH),
		6357 => to_signed(18757, LUT_AMPL_WIDTH),
		6358 => to_signed(18759, LUT_AMPL_WIDTH),
		6359 => to_signed(18762, LUT_AMPL_WIDTH),
		6360 => to_signed(18765, LUT_AMPL_WIDTH),
		6361 => to_signed(18767, LUT_AMPL_WIDTH),
		6362 => to_signed(18770, LUT_AMPL_WIDTH),
		6363 => to_signed(18772, LUT_AMPL_WIDTH),
		6364 => to_signed(18775, LUT_AMPL_WIDTH),
		6365 => to_signed(18778, LUT_AMPL_WIDTH),
		6366 => to_signed(18780, LUT_AMPL_WIDTH),
		6367 => to_signed(18783, LUT_AMPL_WIDTH),
		6368 => to_signed(18785, LUT_AMPL_WIDTH),
		6369 => to_signed(18788, LUT_AMPL_WIDTH),
		6370 => to_signed(18790, LUT_AMPL_WIDTH),
		6371 => to_signed(18793, LUT_AMPL_WIDTH),
		6372 => to_signed(18796, LUT_AMPL_WIDTH),
		6373 => to_signed(18798, LUT_AMPL_WIDTH),
		6374 => to_signed(18801, LUT_AMPL_WIDTH),
		6375 => to_signed(18803, LUT_AMPL_WIDTH),
		6376 => to_signed(18806, LUT_AMPL_WIDTH),
		6377 => to_signed(18808, LUT_AMPL_WIDTH),
		6378 => to_signed(18811, LUT_AMPL_WIDTH),
		6379 => to_signed(18814, LUT_AMPL_WIDTH),
		6380 => to_signed(18816, LUT_AMPL_WIDTH),
		6381 => to_signed(18819, LUT_AMPL_WIDTH),
		6382 => to_signed(18821, LUT_AMPL_WIDTH),
		6383 => to_signed(18824, LUT_AMPL_WIDTH),
		6384 => to_signed(18826, LUT_AMPL_WIDTH),
		6385 => to_signed(18829, LUT_AMPL_WIDTH),
		6386 => to_signed(18832, LUT_AMPL_WIDTH),
		6387 => to_signed(18834, LUT_AMPL_WIDTH),
		6388 => to_signed(18837, LUT_AMPL_WIDTH),
		6389 => to_signed(18839, LUT_AMPL_WIDTH),
		6390 => to_signed(18842, LUT_AMPL_WIDTH),
		6391 => to_signed(18844, LUT_AMPL_WIDTH),
		6392 => to_signed(18847, LUT_AMPL_WIDTH),
		6393 => to_signed(18850, LUT_AMPL_WIDTH),
		6394 => to_signed(18852, LUT_AMPL_WIDTH),
		6395 => to_signed(18855, LUT_AMPL_WIDTH),
		6396 => to_signed(18857, LUT_AMPL_WIDTH),
		6397 => to_signed(18860, LUT_AMPL_WIDTH),
		6398 => to_signed(18862, LUT_AMPL_WIDTH),
		6399 => to_signed(18865, LUT_AMPL_WIDTH),
		6400 => to_signed(18868, LUT_AMPL_WIDTH),
		6401 => to_signed(18870, LUT_AMPL_WIDTH),
		6402 => to_signed(18873, LUT_AMPL_WIDTH),
		6403 => to_signed(18875, LUT_AMPL_WIDTH),
		6404 => to_signed(18878, LUT_AMPL_WIDTH),
		6405 => to_signed(18880, LUT_AMPL_WIDTH),
		6406 => to_signed(18883, LUT_AMPL_WIDTH),
		6407 => to_signed(18885, LUT_AMPL_WIDTH),
		6408 => to_signed(18888, LUT_AMPL_WIDTH),
		6409 => to_signed(18891, LUT_AMPL_WIDTH),
		6410 => to_signed(18893, LUT_AMPL_WIDTH),
		6411 => to_signed(18896, LUT_AMPL_WIDTH),
		6412 => to_signed(18898, LUT_AMPL_WIDTH),
		6413 => to_signed(18901, LUT_AMPL_WIDTH),
		6414 => to_signed(18903, LUT_AMPL_WIDTH),
		6415 => to_signed(18906, LUT_AMPL_WIDTH),
		6416 => to_signed(18909, LUT_AMPL_WIDTH),
		6417 => to_signed(18911, LUT_AMPL_WIDTH),
		6418 => to_signed(18914, LUT_AMPL_WIDTH),
		6419 => to_signed(18916, LUT_AMPL_WIDTH),
		6420 => to_signed(18919, LUT_AMPL_WIDTH),
		6421 => to_signed(18921, LUT_AMPL_WIDTH),
		6422 => to_signed(18924, LUT_AMPL_WIDTH),
		6423 => to_signed(18927, LUT_AMPL_WIDTH),
		6424 => to_signed(18929, LUT_AMPL_WIDTH),
		6425 => to_signed(18932, LUT_AMPL_WIDTH),
		6426 => to_signed(18934, LUT_AMPL_WIDTH),
		6427 => to_signed(18937, LUT_AMPL_WIDTH),
		6428 => to_signed(18939, LUT_AMPL_WIDTH),
		6429 => to_signed(18942, LUT_AMPL_WIDTH),
		6430 => to_signed(18944, LUT_AMPL_WIDTH),
		6431 => to_signed(18947, LUT_AMPL_WIDTH),
		6432 => to_signed(18950, LUT_AMPL_WIDTH),
		6433 => to_signed(18952, LUT_AMPL_WIDTH),
		6434 => to_signed(18955, LUT_AMPL_WIDTH),
		6435 => to_signed(18957, LUT_AMPL_WIDTH),
		6436 => to_signed(18960, LUT_AMPL_WIDTH),
		6437 => to_signed(18962, LUT_AMPL_WIDTH),
		6438 => to_signed(18965, LUT_AMPL_WIDTH),
		6439 => to_signed(18968, LUT_AMPL_WIDTH),
		6440 => to_signed(18970, LUT_AMPL_WIDTH),
		6441 => to_signed(18973, LUT_AMPL_WIDTH),
		6442 => to_signed(18975, LUT_AMPL_WIDTH),
		6443 => to_signed(18978, LUT_AMPL_WIDTH),
		6444 => to_signed(18980, LUT_AMPL_WIDTH),
		6445 => to_signed(18983, LUT_AMPL_WIDTH),
		6446 => to_signed(18985, LUT_AMPL_WIDTH),
		6447 => to_signed(18988, LUT_AMPL_WIDTH),
		6448 => to_signed(18991, LUT_AMPL_WIDTH),
		6449 => to_signed(18993, LUT_AMPL_WIDTH),
		6450 => to_signed(18996, LUT_AMPL_WIDTH),
		6451 => to_signed(18998, LUT_AMPL_WIDTH),
		6452 => to_signed(19001, LUT_AMPL_WIDTH),
		6453 => to_signed(19003, LUT_AMPL_WIDTH),
		6454 => to_signed(19006, LUT_AMPL_WIDTH),
		6455 => to_signed(19009, LUT_AMPL_WIDTH),
		6456 => to_signed(19011, LUT_AMPL_WIDTH),
		6457 => to_signed(19014, LUT_AMPL_WIDTH),
		6458 => to_signed(19016, LUT_AMPL_WIDTH),
		6459 => to_signed(19019, LUT_AMPL_WIDTH),
		6460 => to_signed(19021, LUT_AMPL_WIDTH),
		6461 => to_signed(19024, LUT_AMPL_WIDTH),
		6462 => to_signed(19026, LUT_AMPL_WIDTH),
		6463 => to_signed(19029, LUT_AMPL_WIDTH),
		6464 => to_signed(19032, LUT_AMPL_WIDTH),
		6465 => to_signed(19034, LUT_AMPL_WIDTH),
		6466 => to_signed(19037, LUT_AMPL_WIDTH),
		6467 => to_signed(19039, LUT_AMPL_WIDTH),
		6468 => to_signed(19042, LUT_AMPL_WIDTH),
		6469 => to_signed(19044, LUT_AMPL_WIDTH),
		6470 => to_signed(19047, LUT_AMPL_WIDTH),
		6471 => to_signed(19049, LUT_AMPL_WIDTH),
		6472 => to_signed(19052, LUT_AMPL_WIDTH),
		6473 => to_signed(19055, LUT_AMPL_WIDTH),
		6474 => to_signed(19057, LUT_AMPL_WIDTH),
		6475 => to_signed(19060, LUT_AMPL_WIDTH),
		6476 => to_signed(19062, LUT_AMPL_WIDTH),
		6477 => to_signed(19065, LUT_AMPL_WIDTH),
		6478 => to_signed(19067, LUT_AMPL_WIDTH),
		6479 => to_signed(19070, LUT_AMPL_WIDTH),
		6480 => to_signed(19072, LUT_AMPL_WIDTH),
		6481 => to_signed(19075, LUT_AMPL_WIDTH),
		6482 => to_signed(19078, LUT_AMPL_WIDTH),
		6483 => to_signed(19080, LUT_AMPL_WIDTH),
		6484 => to_signed(19083, LUT_AMPL_WIDTH),
		6485 => to_signed(19085, LUT_AMPL_WIDTH),
		6486 => to_signed(19088, LUT_AMPL_WIDTH),
		6487 => to_signed(19090, LUT_AMPL_WIDTH),
		6488 => to_signed(19093, LUT_AMPL_WIDTH),
		6489 => to_signed(19095, LUT_AMPL_WIDTH),
		6490 => to_signed(19098, LUT_AMPL_WIDTH),
		6491 => to_signed(19101, LUT_AMPL_WIDTH),
		6492 => to_signed(19103, LUT_AMPL_WIDTH),
		6493 => to_signed(19106, LUT_AMPL_WIDTH),
		6494 => to_signed(19108, LUT_AMPL_WIDTH),
		6495 => to_signed(19111, LUT_AMPL_WIDTH),
		6496 => to_signed(19113, LUT_AMPL_WIDTH),
		6497 => to_signed(19116, LUT_AMPL_WIDTH),
		6498 => to_signed(19118, LUT_AMPL_WIDTH),
		6499 => to_signed(19121, LUT_AMPL_WIDTH),
		6500 => to_signed(19123, LUT_AMPL_WIDTH),
		6501 => to_signed(19126, LUT_AMPL_WIDTH),
		6502 => to_signed(19129, LUT_AMPL_WIDTH),
		6503 => to_signed(19131, LUT_AMPL_WIDTH),
		6504 => to_signed(19134, LUT_AMPL_WIDTH),
		6505 => to_signed(19136, LUT_AMPL_WIDTH),
		6506 => to_signed(19139, LUT_AMPL_WIDTH),
		6507 => to_signed(19141, LUT_AMPL_WIDTH),
		6508 => to_signed(19144, LUT_AMPL_WIDTH),
		6509 => to_signed(19146, LUT_AMPL_WIDTH),
		6510 => to_signed(19149, LUT_AMPL_WIDTH),
		6511 => to_signed(19152, LUT_AMPL_WIDTH),
		6512 => to_signed(19154, LUT_AMPL_WIDTH),
		6513 => to_signed(19157, LUT_AMPL_WIDTH),
		6514 => to_signed(19159, LUT_AMPL_WIDTH),
		6515 => to_signed(19162, LUT_AMPL_WIDTH),
		6516 => to_signed(19164, LUT_AMPL_WIDTH),
		6517 => to_signed(19167, LUT_AMPL_WIDTH),
		6518 => to_signed(19169, LUT_AMPL_WIDTH),
		6519 => to_signed(19172, LUT_AMPL_WIDTH),
		6520 => to_signed(19174, LUT_AMPL_WIDTH),
		6521 => to_signed(19177, LUT_AMPL_WIDTH),
		6522 => to_signed(19180, LUT_AMPL_WIDTH),
		6523 => to_signed(19182, LUT_AMPL_WIDTH),
		6524 => to_signed(19185, LUT_AMPL_WIDTH),
		6525 => to_signed(19187, LUT_AMPL_WIDTH),
		6526 => to_signed(19190, LUT_AMPL_WIDTH),
		6527 => to_signed(19192, LUT_AMPL_WIDTH),
		6528 => to_signed(19195, LUT_AMPL_WIDTH),
		6529 => to_signed(19197, LUT_AMPL_WIDTH),
		6530 => to_signed(19200, LUT_AMPL_WIDTH),
		6531 => to_signed(19202, LUT_AMPL_WIDTH),
		6532 => to_signed(19205, LUT_AMPL_WIDTH),
		6533 => to_signed(19208, LUT_AMPL_WIDTH),
		6534 => to_signed(19210, LUT_AMPL_WIDTH),
		6535 => to_signed(19213, LUT_AMPL_WIDTH),
		6536 => to_signed(19215, LUT_AMPL_WIDTH),
		6537 => to_signed(19218, LUT_AMPL_WIDTH),
		6538 => to_signed(19220, LUT_AMPL_WIDTH),
		6539 => to_signed(19223, LUT_AMPL_WIDTH),
		6540 => to_signed(19225, LUT_AMPL_WIDTH),
		6541 => to_signed(19228, LUT_AMPL_WIDTH),
		6542 => to_signed(19230, LUT_AMPL_WIDTH),
		6543 => to_signed(19233, LUT_AMPL_WIDTH),
		6544 => to_signed(19236, LUT_AMPL_WIDTH),
		6545 => to_signed(19238, LUT_AMPL_WIDTH),
		6546 => to_signed(19241, LUT_AMPL_WIDTH),
		6547 => to_signed(19243, LUT_AMPL_WIDTH),
		6548 => to_signed(19246, LUT_AMPL_WIDTH),
		6549 => to_signed(19248, LUT_AMPL_WIDTH),
		6550 => to_signed(19251, LUT_AMPL_WIDTH),
		6551 => to_signed(19253, LUT_AMPL_WIDTH),
		6552 => to_signed(19256, LUT_AMPL_WIDTH),
		6553 => to_signed(19258, LUT_AMPL_WIDTH),
		6554 => to_signed(19261, LUT_AMPL_WIDTH),
		6555 => to_signed(19264, LUT_AMPL_WIDTH),
		6556 => to_signed(19266, LUT_AMPL_WIDTH),
		6557 => to_signed(19269, LUT_AMPL_WIDTH),
		6558 => to_signed(19271, LUT_AMPL_WIDTH),
		6559 => to_signed(19274, LUT_AMPL_WIDTH),
		6560 => to_signed(19276, LUT_AMPL_WIDTH),
		6561 => to_signed(19279, LUT_AMPL_WIDTH),
		6562 => to_signed(19281, LUT_AMPL_WIDTH),
		6563 => to_signed(19284, LUT_AMPL_WIDTH),
		6564 => to_signed(19286, LUT_AMPL_WIDTH),
		6565 => to_signed(19289, LUT_AMPL_WIDTH),
		6566 => to_signed(19291, LUT_AMPL_WIDTH),
		6567 => to_signed(19294, LUT_AMPL_WIDTH),
		6568 => to_signed(19297, LUT_AMPL_WIDTH),
		6569 => to_signed(19299, LUT_AMPL_WIDTH),
		6570 => to_signed(19302, LUT_AMPL_WIDTH),
		6571 => to_signed(19304, LUT_AMPL_WIDTH),
		6572 => to_signed(19307, LUT_AMPL_WIDTH),
		6573 => to_signed(19309, LUT_AMPL_WIDTH),
		6574 => to_signed(19312, LUT_AMPL_WIDTH),
		6575 => to_signed(19314, LUT_AMPL_WIDTH),
		6576 => to_signed(19317, LUT_AMPL_WIDTH),
		6577 => to_signed(19319, LUT_AMPL_WIDTH),
		6578 => to_signed(19322, LUT_AMPL_WIDTH),
		6579 => to_signed(19324, LUT_AMPL_WIDTH),
		6580 => to_signed(19327, LUT_AMPL_WIDTH),
		6581 => to_signed(19330, LUT_AMPL_WIDTH),
		6582 => to_signed(19332, LUT_AMPL_WIDTH),
		6583 => to_signed(19335, LUT_AMPL_WIDTH),
		6584 => to_signed(19337, LUT_AMPL_WIDTH),
		6585 => to_signed(19340, LUT_AMPL_WIDTH),
		6586 => to_signed(19342, LUT_AMPL_WIDTH),
		6587 => to_signed(19345, LUT_AMPL_WIDTH),
		6588 => to_signed(19347, LUT_AMPL_WIDTH),
		6589 => to_signed(19350, LUT_AMPL_WIDTH),
		6590 => to_signed(19352, LUT_AMPL_WIDTH),
		6591 => to_signed(19355, LUT_AMPL_WIDTH),
		6592 => to_signed(19357, LUT_AMPL_WIDTH),
		6593 => to_signed(19360, LUT_AMPL_WIDTH),
		6594 => to_signed(19362, LUT_AMPL_WIDTH),
		6595 => to_signed(19365, LUT_AMPL_WIDTH),
		6596 => to_signed(19368, LUT_AMPL_WIDTH),
		6597 => to_signed(19370, LUT_AMPL_WIDTH),
		6598 => to_signed(19373, LUT_AMPL_WIDTH),
		6599 => to_signed(19375, LUT_AMPL_WIDTH),
		6600 => to_signed(19378, LUT_AMPL_WIDTH),
		6601 => to_signed(19380, LUT_AMPL_WIDTH),
		6602 => to_signed(19383, LUT_AMPL_WIDTH),
		6603 => to_signed(19385, LUT_AMPL_WIDTH),
		6604 => to_signed(19388, LUT_AMPL_WIDTH),
		6605 => to_signed(19390, LUT_AMPL_WIDTH),
		6606 => to_signed(19393, LUT_AMPL_WIDTH),
		6607 => to_signed(19395, LUT_AMPL_WIDTH),
		6608 => to_signed(19398, LUT_AMPL_WIDTH),
		6609 => to_signed(19400, LUT_AMPL_WIDTH),
		6610 => to_signed(19403, LUT_AMPL_WIDTH),
		6611 => to_signed(19406, LUT_AMPL_WIDTH),
		6612 => to_signed(19408, LUT_AMPL_WIDTH),
		6613 => to_signed(19411, LUT_AMPL_WIDTH),
		6614 => to_signed(19413, LUT_AMPL_WIDTH),
		6615 => to_signed(19416, LUT_AMPL_WIDTH),
		6616 => to_signed(19418, LUT_AMPL_WIDTH),
		6617 => to_signed(19421, LUT_AMPL_WIDTH),
		6618 => to_signed(19423, LUT_AMPL_WIDTH),
		6619 => to_signed(19426, LUT_AMPL_WIDTH),
		6620 => to_signed(19428, LUT_AMPL_WIDTH),
		6621 => to_signed(19431, LUT_AMPL_WIDTH),
		6622 => to_signed(19433, LUT_AMPL_WIDTH),
		6623 => to_signed(19436, LUT_AMPL_WIDTH),
		6624 => to_signed(19438, LUT_AMPL_WIDTH),
		6625 => to_signed(19441, LUT_AMPL_WIDTH),
		6626 => to_signed(19444, LUT_AMPL_WIDTH),
		6627 => to_signed(19446, LUT_AMPL_WIDTH),
		6628 => to_signed(19449, LUT_AMPL_WIDTH),
		6629 => to_signed(19451, LUT_AMPL_WIDTH),
		6630 => to_signed(19454, LUT_AMPL_WIDTH),
		6631 => to_signed(19456, LUT_AMPL_WIDTH),
		6632 => to_signed(19459, LUT_AMPL_WIDTH),
		6633 => to_signed(19461, LUT_AMPL_WIDTH),
		6634 => to_signed(19464, LUT_AMPL_WIDTH),
		6635 => to_signed(19466, LUT_AMPL_WIDTH),
		6636 => to_signed(19469, LUT_AMPL_WIDTH),
		6637 => to_signed(19471, LUT_AMPL_WIDTH),
		6638 => to_signed(19474, LUT_AMPL_WIDTH),
		6639 => to_signed(19476, LUT_AMPL_WIDTH),
		6640 => to_signed(19479, LUT_AMPL_WIDTH),
		6641 => to_signed(19481, LUT_AMPL_WIDTH),
		6642 => to_signed(19484, LUT_AMPL_WIDTH),
		6643 => to_signed(19486, LUT_AMPL_WIDTH),
		6644 => to_signed(19489, LUT_AMPL_WIDTH),
		6645 => to_signed(19492, LUT_AMPL_WIDTH),
		6646 => to_signed(19494, LUT_AMPL_WIDTH),
		6647 => to_signed(19497, LUT_AMPL_WIDTH),
		6648 => to_signed(19499, LUT_AMPL_WIDTH),
		6649 => to_signed(19502, LUT_AMPL_WIDTH),
		6650 => to_signed(19504, LUT_AMPL_WIDTH),
		6651 => to_signed(19507, LUT_AMPL_WIDTH),
		6652 => to_signed(19509, LUT_AMPL_WIDTH),
		6653 => to_signed(19512, LUT_AMPL_WIDTH),
		6654 => to_signed(19514, LUT_AMPL_WIDTH),
		6655 => to_signed(19517, LUT_AMPL_WIDTH),
		6656 => to_signed(19519, LUT_AMPL_WIDTH),
		6657 => to_signed(19522, LUT_AMPL_WIDTH),
		6658 => to_signed(19524, LUT_AMPL_WIDTH),
		6659 => to_signed(19527, LUT_AMPL_WIDTH),
		6660 => to_signed(19529, LUT_AMPL_WIDTH),
		6661 => to_signed(19532, LUT_AMPL_WIDTH),
		6662 => to_signed(19534, LUT_AMPL_WIDTH),
		6663 => to_signed(19537, LUT_AMPL_WIDTH),
		6664 => to_signed(19539, LUT_AMPL_WIDTH),
		6665 => to_signed(19542, LUT_AMPL_WIDTH),
		6666 => to_signed(19545, LUT_AMPL_WIDTH),
		6667 => to_signed(19547, LUT_AMPL_WIDTH),
		6668 => to_signed(19550, LUT_AMPL_WIDTH),
		6669 => to_signed(19552, LUT_AMPL_WIDTH),
		6670 => to_signed(19555, LUT_AMPL_WIDTH),
		6671 => to_signed(19557, LUT_AMPL_WIDTH),
		6672 => to_signed(19560, LUT_AMPL_WIDTH),
		6673 => to_signed(19562, LUT_AMPL_WIDTH),
		6674 => to_signed(19565, LUT_AMPL_WIDTH),
		6675 => to_signed(19567, LUT_AMPL_WIDTH),
		6676 => to_signed(19570, LUT_AMPL_WIDTH),
		6677 => to_signed(19572, LUT_AMPL_WIDTH),
		6678 => to_signed(19575, LUT_AMPL_WIDTH),
		6679 => to_signed(19577, LUT_AMPL_WIDTH),
		6680 => to_signed(19580, LUT_AMPL_WIDTH),
		6681 => to_signed(19582, LUT_AMPL_WIDTH),
		6682 => to_signed(19585, LUT_AMPL_WIDTH),
		6683 => to_signed(19587, LUT_AMPL_WIDTH),
		6684 => to_signed(19590, LUT_AMPL_WIDTH),
		6685 => to_signed(19592, LUT_AMPL_WIDTH),
		6686 => to_signed(19595, LUT_AMPL_WIDTH),
		6687 => to_signed(19597, LUT_AMPL_WIDTH),
		6688 => to_signed(19600, LUT_AMPL_WIDTH),
		6689 => to_signed(19602, LUT_AMPL_WIDTH),
		6690 => to_signed(19605, LUT_AMPL_WIDTH),
		6691 => to_signed(19607, LUT_AMPL_WIDTH),
		6692 => to_signed(19610, LUT_AMPL_WIDTH),
		6693 => to_signed(19613, LUT_AMPL_WIDTH),
		6694 => to_signed(19615, LUT_AMPL_WIDTH),
		6695 => to_signed(19618, LUT_AMPL_WIDTH),
		6696 => to_signed(19620, LUT_AMPL_WIDTH),
		6697 => to_signed(19623, LUT_AMPL_WIDTH),
		6698 => to_signed(19625, LUT_AMPL_WIDTH),
		6699 => to_signed(19628, LUT_AMPL_WIDTH),
		6700 => to_signed(19630, LUT_AMPL_WIDTH),
		6701 => to_signed(19633, LUT_AMPL_WIDTH),
		6702 => to_signed(19635, LUT_AMPL_WIDTH),
		6703 => to_signed(19638, LUT_AMPL_WIDTH),
		6704 => to_signed(19640, LUT_AMPL_WIDTH),
		6705 => to_signed(19643, LUT_AMPL_WIDTH),
		6706 => to_signed(19645, LUT_AMPL_WIDTH),
		6707 => to_signed(19648, LUT_AMPL_WIDTH),
		6708 => to_signed(19650, LUT_AMPL_WIDTH),
		6709 => to_signed(19653, LUT_AMPL_WIDTH),
		6710 => to_signed(19655, LUT_AMPL_WIDTH),
		6711 => to_signed(19658, LUT_AMPL_WIDTH),
		6712 => to_signed(19660, LUT_AMPL_WIDTH),
		6713 => to_signed(19663, LUT_AMPL_WIDTH),
		6714 => to_signed(19665, LUT_AMPL_WIDTH),
		6715 => to_signed(19668, LUT_AMPL_WIDTH),
		6716 => to_signed(19670, LUT_AMPL_WIDTH),
		6717 => to_signed(19673, LUT_AMPL_WIDTH),
		6718 => to_signed(19675, LUT_AMPL_WIDTH),
		6719 => to_signed(19678, LUT_AMPL_WIDTH),
		6720 => to_signed(19680, LUT_AMPL_WIDTH),
		6721 => to_signed(19683, LUT_AMPL_WIDTH),
		6722 => to_signed(19685, LUT_AMPL_WIDTH),
		6723 => to_signed(19688, LUT_AMPL_WIDTH),
		6724 => to_signed(19690, LUT_AMPL_WIDTH),
		6725 => to_signed(19693, LUT_AMPL_WIDTH),
		6726 => to_signed(19695, LUT_AMPL_WIDTH),
		6727 => to_signed(19698, LUT_AMPL_WIDTH),
		6728 => to_signed(19700, LUT_AMPL_WIDTH),
		6729 => to_signed(19703, LUT_AMPL_WIDTH),
		6730 => to_signed(19706, LUT_AMPL_WIDTH),
		6731 => to_signed(19708, LUT_AMPL_WIDTH),
		6732 => to_signed(19711, LUT_AMPL_WIDTH),
		6733 => to_signed(19713, LUT_AMPL_WIDTH),
		6734 => to_signed(19716, LUT_AMPL_WIDTH),
		6735 => to_signed(19718, LUT_AMPL_WIDTH),
		6736 => to_signed(19721, LUT_AMPL_WIDTH),
		6737 => to_signed(19723, LUT_AMPL_WIDTH),
		6738 => to_signed(19726, LUT_AMPL_WIDTH),
		6739 => to_signed(19728, LUT_AMPL_WIDTH),
		6740 => to_signed(19731, LUT_AMPL_WIDTH),
		6741 => to_signed(19733, LUT_AMPL_WIDTH),
		6742 => to_signed(19736, LUT_AMPL_WIDTH),
		6743 => to_signed(19738, LUT_AMPL_WIDTH),
		6744 => to_signed(19741, LUT_AMPL_WIDTH),
		6745 => to_signed(19743, LUT_AMPL_WIDTH),
		6746 => to_signed(19746, LUT_AMPL_WIDTH),
		6747 => to_signed(19748, LUT_AMPL_WIDTH),
		6748 => to_signed(19751, LUT_AMPL_WIDTH),
		6749 => to_signed(19753, LUT_AMPL_WIDTH),
		6750 => to_signed(19756, LUT_AMPL_WIDTH),
		6751 => to_signed(19758, LUT_AMPL_WIDTH),
		6752 => to_signed(19761, LUT_AMPL_WIDTH),
		6753 => to_signed(19763, LUT_AMPL_WIDTH),
		6754 => to_signed(19766, LUT_AMPL_WIDTH),
		6755 => to_signed(19768, LUT_AMPL_WIDTH),
		6756 => to_signed(19771, LUT_AMPL_WIDTH),
		6757 => to_signed(19773, LUT_AMPL_WIDTH),
		6758 => to_signed(19776, LUT_AMPL_WIDTH),
		6759 => to_signed(19778, LUT_AMPL_WIDTH),
		6760 => to_signed(19781, LUT_AMPL_WIDTH),
		6761 => to_signed(19783, LUT_AMPL_WIDTH),
		6762 => to_signed(19786, LUT_AMPL_WIDTH),
		6763 => to_signed(19788, LUT_AMPL_WIDTH),
		6764 => to_signed(19791, LUT_AMPL_WIDTH),
		6765 => to_signed(19793, LUT_AMPL_WIDTH),
		6766 => to_signed(19796, LUT_AMPL_WIDTH),
		6767 => to_signed(19798, LUT_AMPL_WIDTH),
		6768 => to_signed(19801, LUT_AMPL_WIDTH),
		6769 => to_signed(19803, LUT_AMPL_WIDTH),
		6770 => to_signed(19806, LUT_AMPL_WIDTH),
		6771 => to_signed(19808, LUT_AMPL_WIDTH),
		6772 => to_signed(19811, LUT_AMPL_WIDTH),
		6773 => to_signed(19813, LUT_AMPL_WIDTH),
		6774 => to_signed(19816, LUT_AMPL_WIDTH),
		6775 => to_signed(19818, LUT_AMPL_WIDTH),
		6776 => to_signed(19821, LUT_AMPL_WIDTH),
		6777 => to_signed(19823, LUT_AMPL_WIDTH),
		6778 => to_signed(19826, LUT_AMPL_WIDTH),
		6779 => to_signed(19828, LUT_AMPL_WIDTH),
		6780 => to_signed(19831, LUT_AMPL_WIDTH),
		6781 => to_signed(19833, LUT_AMPL_WIDTH),
		6782 => to_signed(19836, LUT_AMPL_WIDTH),
		6783 => to_signed(19838, LUT_AMPL_WIDTH),
		6784 => to_signed(19841, LUT_AMPL_WIDTH),
		6785 => to_signed(19843, LUT_AMPL_WIDTH),
		6786 => to_signed(19846, LUT_AMPL_WIDTH),
		6787 => to_signed(19848, LUT_AMPL_WIDTH),
		6788 => to_signed(19851, LUT_AMPL_WIDTH),
		6789 => to_signed(19853, LUT_AMPL_WIDTH),
		6790 => to_signed(19856, LUT_AMPL_WIDTH),
		6791 => to_signed(19858, LUT_AMPL_WIDTH),
		6792 => to_signed(19861, LUT_AMPL_WIDTH),
		6793 => to_signed(19863, LUT_AMPL_WIDTH),
		6794 => to_signed(19866, LUT_AMPL_WIDTH),
		6795 => to_signed(19868, LUT_AMPL_WIDTH),
		6796 => to_signed(19871, LUT_AMPL_WIDTH),
		6797 => to_signed(19873, LUT_AMPL_WIDTH),
		6798 => to_signed(19876, LUT_AMPL_WIDTH),
		6799 => to_signed(19878, LUT_AMPL_WIDTH),
		6800 => to_signed(19881, LUT_AMPL_WIDTH),
		6801 => to_signed(19883, LUT_AMPL_WIDTH),
		6802 => to_signed(19886, LUT_AMPL_WIDTH),
		6803 => to_signed(19888, LUT_AMPL_WIDTH),
		6804 => to_signed(19891, LUT_AMPL_WIDTH),
		6805 => to_signed(19893, LUT_AMPL_WIDTH),
		6806 => to_signed(19896, LUT_AMPL_WIDTH),
		6807 => to_signed(19898, LUT_AMPL_WIDTH),
		6808 => to_signed(19901, LUT_AMPL_WIDTH),
		6809 => to_signed(19903, LUT_AMPL_WIDTH),
		6810 => to_signed(19906, LUT_AMPL_WIDTH),
		6811 => to_signed(19908, LUT_AMPL_WIDTH),
		6812 => to_signed(19911, LUT_AMPL_WIDTH),
		6813 => to_signed(19913, LUT_AMPL_WIDTH),
		6814 => to_signed(19916, LUT_AMPL_WIDTH),
		6815 => to_signed(19918, LUT_AMPL_WIDTH),
		6816 => to_signed(19921, LUT_AMPL_WIDTH),
		6817 => to_signed(19923, LUT_AMPL_WIDTH),
		6818 => to_signed(19926, LUT_AMPL_WIDTH),
		6819 => to_signed(19928, LUT_AMPL_WIDTH),
		6820 => to_signed(19931, LUT_AMPL_WIDTH),
		6821 => to_signed(19933, LUT_AMPL_WIDTH),
		6822 => to_signed(19936, LUT_AMPL_WIDTH),
		6823 => to_signed(19938, LUT_AMPL_WIDTH),
		6824 => to_signed(19941, LUT_AMPL_WIDTH),
		6825 => to_signed(19943, LUT_AMPL_WIDTH),
		6826 => to_signed(19946, LUT_AMPL_WIDTH),
		6827 => to_signed(19948, LUT_AMPL_WIDTH),
		6828 => to_signed(19951, LUT_AMPL_WIDTH),
		6829 => to_signed(19953, LUT_AMPL_WIDTH),
		6830 => to_signed(19956, LUT_AMPL_WIDTH),
		6831 => to_signed(19958, LUT_AMPL_WIDTH),
		6832 => to_signed(19961, LUT_AMPL_WIDTH),
		6833 => to_signed(19963, LUT_AMPL_WIDTH),
		6834 => to_signed(19966, LUT_AMPL_WIDTH),
		6835 => to_signed(19968, LUT_AMPL_WIDTH),
		6836 => to_signed(19971, LUT_AMPL_WIDTH),
		6837 => to_signed(19973, LUT_AMPL_WIDTH),
		6838 => to_signed(19976, LUT_AMPL_WIDTH),
		6839 => to_signed(19978, LUT_AMPL_WIDTH),
		6840 => to_signed(19981, LUT_AMPL_WIDTH),
		6841 => to_signed(19983, LUT_AMPL_WIDTH),
		6842 => to_signed(19985, LUT_AMPL_WIDTH),
		6843 => to_signed(19988, LUT_AMPL_WIDTH),
		6844 => to_signed(19990, LUT_AMPL_WIDTH),
		6845 => to_signed(19993, LUT_AMPL_WIDTH),
		6846 => to_signed(19995, LUT_AMPL_WIDTH),
		6847 => to_signed(19998, LUT_AMPL_WIDTH),
		6848 => to_signed(20000, LUT_AMPL_WIDTH),
		6849 => to_signed(20003, LUT_AMPL_WIDTH),
		6850 => to_signed(20005, LUT_AMPL_WIDTH),
		6851 => to_signed(20008, LUT_AMPL_WIDTH),
		6852 => to_signed(20010, LUT_AMPL_WIDTH),
		6853 => to_signed(20013, LUT_AMPL_WIDTH),
		6854 => to_signed(20015, LUT_AMPL_WIDTH),
		6855 => to_signed(20018, LUT_AMPL_WIDTH),
		6856 => to_signed(20020, LUT_AMPL_WIDTH),
		6857 => to_signed(20023, LUT_AMPL_WIDTH),
		6858 => to_signed(20025, LUT_AMPL_WIDTH),
		6859 => to_signed(20028, LUT_AMPL_WIDTH),
		6860 => to_signed(20030, LUT_AMPL_WIDTH),
		6861 => to_signed(20033, LUT_AMPL_WIDTH),
		6862 => to_signed(20035, LUT_AMPL_WIDTH),
		6863 => to_signed(20038, LUT_AMPL_WIDTH),
		6864 => to_signed(20040, LUT_AMPL_WIDTH),
		6865 => to_signed(20043, LUT_AMPL_WIDTH),
		6866 => to_signed(20045, LUT_AMPL_WIDTH),
		6867 => to_signed(20048, LUT_AMPL_WIDTH),
		6868 => to_signed(20050, LUT_AMPL_WIDTH),
		6869 => to_signed(20053, LUT_AMPL_WIDTH),
		6870 => to_signed(20055, LUT_AMPL_WIDTH),
		6871 => to_signed(20058, LUT_AMPL_WIDTH),
		6872 => to_signed(20060, LUT_AMPL_WIDTH),
		6873 => to_signed(20063, LUT_AMPL_WIDTH),
		6874 => to_signed(20065, LUT_AMPL_WIDTH),
		6875 => to_signed(20068, LUT_AMPL_WIDTH),
		6876 => to_signed(20070, LUT_AMPL_WIDTH),
		6877 => to_signed(20072, LUT_AMPL_WIDTH),
		6878 => to_signed(20075, LUT_AMPL_WIDTH),
		6879 => to_signed(20077, LUT_AMPL_WIDTH),
		6880 => to_signed(20080, LUT_AMPL_WIDTH),
		6881 => to_signed(20082, LUT_AMPL_WIDTH),
		6882 => to_signed(20085, LUT_AMPL_WIDTH),
		6883 => to_signed(20087, LUT_AMPL_WIDTH),
		6884 => to_signed(20090, LUT_AMPL_WIDTH),
		6885 => to_signed(20092, LUT_AMPL_WIDTH),
		6886 => to_signed(20095, LUT_AMPL_WIDTH),
		6887 => to_signed(20097, LUT_AMPL_WIDTH),
		6888 => to_signed(20100, LUT_AMPL_WIDTH),
		6889 => to_signed(20102, LUT_AMPL_WIDTH),
		6890 => to_signed(20105, LUT_AMPL_WIDTH),
		6891 => to_signed(20107, LUT_AMPL_WIDTH),
		6892 => to_signed(20110, LUT_AMPL_WIDTH),
		6893 => to_signed(20112, LUT_AMPL_WIDTH),
		6894 => to_signed(20115, LUT_AMPL_WIDTH),
		6895 => to_signed(20117, LUT_AMPL_WIDTH),
		6896 => to_signed(20120, LUT_AMPL_WIDTH),
		6897 => to_signed(20122, LUT_AMPL_WIDTH),
		6898 => to_signed(20125, LUT_AMPL_WIDTH),
		6899 => to_signed(20127, LUT_AMPL_WIDTH),
		6900 => to_signed(20130, LUT_AMPL_WIDTH),
		6901 => to_signed(20132, LUT_AMPL_WIDTH),
		6902 => to_signed(20135, LUT_AMPL_WIDTH),
		6903 => to_signed(20137, LUT_AMPL_WIDTH),
		6904 => to_signed(20139, LUT_AMPL_WIDTH),
		6905 => to_signed(20142, LUT_AMPL_WIDTH),
		6906 => to_signed(20144, LUT_AMPL_WIDTH),
		6907 => to_signed(20147, LUT_AMPL_WIDTH),
		6908 => to_signed(20149, LUT_AMPL_WIDTH),
		6909 => to_signed(20152, LUT_AMPL_WIDTH),
		6910 => to_signed(20154, LUT_AMPL_WIDTH),
		6911 => to_signed(20157, LUT_AMPL_WIDTH),
		6912 => to_signed(20159, LUT_AMPL_WIDTH),
		6913 => to_signed(20162, LUT_AMPL_WIDTH),
		6914 => to_signed(20164, LUT_AMPL_WIDTH),
		6915 => to_signed(20167, LUT_AMPL_WIDTH),
		6916 => to_signed(20169, LUT_AMPL_WIDTH),
		6917 => to_signed(20172, LUT_AMPL_WIDTH),
		6918 => to_signed(20174, LUT_AMPL_WIDTH),
		6919 => to_signed(20177, LUT_AMPL_WIDTH),
		6920 => to_signed(20179, LUT_AMPL_WIDTH),
		6921 => to_signed(20182, LUT_AMPL_WIDTH),
		6922 => to_signed(20184, LUT_AMPL_WIDTH),
		6923 => to_signed(20187, LUT_AMPL_WIDTH),
		6924 => to_signed(20189, LUT_AMPL_WIDTH),
		6925 => to_signed(20191, LUT_AMPL_WIDTH),
		6926 => to_signed(20194, LUT_AMPL_WIDTH),
		6927 => to_signed(20196, LUT_AMPL_WIDTH),
		6928 => to_signed(20199, LUT_AMPL_WIDTH),
		6929 => to_signed(20201, LUT_AMPL_WIDTH),
		6930 => to_signed(20204, LUT_AMPL_WIDTH),
		6931 => to_signed(20206, LUT_AMPL_WIDTH),
		6932 => to_signed(20209, LUT_AMPL_WIDTH),
		6933 => to_signed(20211, LUT_AMPL_WIDTH),
		6934 => to_signed(20214, LUT_AMPL_WIDTH),
		6935 => to_signed(20216, LUT_AMPL_WIDTH),
		6936 => to_signed(20219, LUT_AMPL_WIDTH),
		6937 => to_signed(20221, LUT_AMPL_WIDTH),
		6938 => to_signed(20224, LUT_AMPL_WIDTH),
		6939 => to_signed(20226, LUT_AMPL_WIDTH),
		6940 => to_signed(20229, LUT_AMPL_WIDTH),
		6941 => to_signed(20231, LUT_AMPL_WIDTH),
		6942 => to_signed(20234, LUT_AMPL_WIDTH),
		6943 => to_signed(20236, LUT_AMPL_WIDTH),
		6944 => to_signed(20238, LUT_AMPL_WIDTH),
		6945 => to_signed(20241, LUT_AMPL_WIDTH),
		6946 => to_signed(20243, LUT_AMPL_WIDTH),
		6947 => to_signed(20246, LUT_AMPL_WIDTH),
		6948 => to_signed(20248, LUT_AMPL_WIDTH),
		6949 => to_signed(20251, LUT_AMPL_WIDTH),
		6950 => to_signed(20253, LUT_AMPL_WIDTH),
		6951 => to_signed(20256, LUT_AMPL_WIDTH),
		6952 => to_signed(20258, LUT_AMPL_WIDTH),
		6953 => to_signed(20261, LUT_AMPL_WIDTH),
		6954 => to_signed(20263, LUT_AMPL_WIDTH),
		6955 => to_signed(20266, LUT_AMPL_WIDTH),
		6956 => to_signed(20268, LUT_AMPL_WIDTH),
		6957 => to_signed(20271, LUT_AMPL_WIDTH),
		6958 => to_signed(20273, LUT_AMPL_WIDTH),
		6959 => to_signed(20275, LUT_AMPL_WIDTH),
		6960 => to_signed(20278, LUT_AMPL_WIDTH),
		6961 => to_signed(20280, LUT_AMPL_WIDTH),
		6962 => to_signed(20283, LUT_AMPL_WIDTH),
		6963 => to_signed(20285, LUT_AMPL_WIDTH),
		6964 => to_signed(20288, LUT_AMPL_WIDTH),
		6965 => to_signed(20290, LUT_AMPL_WIDTH),
		6966 => to_signed(20293, LUT_AMPL_WIDTH),
		6967 => to_signed(20295, LUT_AMPL_WIDTH),
		6968 => to_signed(20298, LUT_AMPL_WIDTH),
		6969 => to_signed(20300, LUT_AMPL_WIDTH),
		6970 => to_signed(20303, LUT_AMPL_WIDTH),
		6971 => to_signed(20305, LUT_AMPL_WIDTH),
		6972 => to_signed(20308, LUT_AMPL_WIDTH),
		6973 => to_signed(20310, LUT_AMPL_WIDTH),
		6974 => to_signed(20312, LUT_AMPL_WIDTH),
		6975 => to_signed(20315, LUT_AMPL_WIDTH),
		6976 => to_signed(20317, LUT_AMPL_WIDTH),
		6977 => to_signed(20320, LUT_AMPL_WIDTH),
		6978 => to_signed(20322, LUT_AMPL_WIDTH),
		6979 => to_signed(20325, LUT_AMPL_WIDTH),
		6980 => to_signed(20327, LUT_AMPL_WIDTH),
		6981 => to_signed(20330, LUT_AMPL_WIDTH),
		6982 => to_signed(20332, LUT_AMPL_WIDTH),
		6983 => to_signed(20335, LUT_AMPL_WIDTH),
		6984 => to_signed(20337, LUT_AMPL_WIDTH),
		6985 => to_signed(20340, LUT_AMPL_WIDTH),
		6986 => to_signed(20342, LUT_AMPL_WIDTH),
		6987 => to_signed(20345, LUT_AMPL_WIDTH),
		6988 => to_signed(20347, LUT_AMPL_WIDTH),
		6989 => to_signed(20349, LUT_AMPL_WIDTH),
		6990 => to_signed(20352, LUT_AMPL_WIDTH),
		6991 => to_signed(20354, LUT_AMPL_WIDTH),
		6992 => to_signed(20357, LUT_AMPL_WIDTH),
		6993 => to_signed(20359, LUT_AMPL_WIDTH),
		6994 => to_signed(20362, LUT_AMPL_WIDTH),
		6995 => to_signed(20364, LUT_AMPL_WIDTH),
		6996 => to_signed(20367, LUT_AMPL_WIDTH),
		6997 => to_signed(20369, LUT_AMPL_WIDTH),
		6998 => to_signed(20372, LUT_AMPL_WIDTH),
		6999 => to_signed(20374, LUT_AMPL_WIDTH),
		7000 => to_signed(20377, LUT_AMPL_WIDTH),
		7001 => to_signed(20379, LUT_AMPL_WIDTH),
		7002 => to_signed(20381, LUT_AMPL_WIDTH),
		7003 => to_signed(20384, LUT_AMPL_WIDTH),
		7004 => to_signed(20386, LUT_AMPL_WIDTH),
		7005 => to_signed(20389, LUT_AMPL_WIDTH),
		7006 => to_signed(20391, LUT_AMPL_WIDTH),
		7007 => to_signed(20394, LUT_AMPL_WIDTH),
		7008 => to_signed(20396, LUT_AMPL_WIDTH),
		7009 => to_signed(20399, LUT_AMPL_WIDTH),
		7010 => to_signed(20401, LUT_AMPL_WIDTH),
		7011 => to_signed(20404, LUT_AMPL_WIDTH),
		7012 => to_signed(20406, LUT_AMPL_WIDTH),
		7013 => to_signed(20408, LUT_AMPL_WIDTH),
		7014 => to_signed(20411, LUT_AMPL_WIDTH),
		7015 => to_signed(20413, LUT_AMPL_WIDTH),
		7016 => to_signed(20416, LUT_AMPL_WIDTH),
		7017 => to_signed(20418, LUT_AMPL_WIDTH),
		7018 => to_signed(20421, LUT_AMPL_WIDTH),
		7019 => to_signed(20423, LUT_AMPL_WIDTH),
		7020 => to_signed(20426, LUT_AMPL_WIDTH),
		7021 => to_signed(20428, LUT_AMPL_WIDTH),
		7022 => to_signed(20431, LUT_AMPL_WIDTH),
		7023 => to_signed(20433, LUT_AMPL_WIDTH),
		7024 => to_signed(20436, LUT_AMPL_WIDTH),
		7025 => to_signed(20438, LUT_AMPL_WIDTH),
		7026 => to_signed(20440, LUT_AMPL_WIDTH),
		7027 => to_signed(20443, LUT_AMPL_WIDTH),
		7028 => to_signed(20445, LUT_AMPL_WIDTH),
		7029 => to_signed(20448, LUT_AMPL_WIDTH),
		7030 => to_signed(20450, LUT_AMPL_WIDTH),
		7031 => to_signed(20453, LUT_AMPL_WIDTH),
		7032 => to_signed(20455, LUT_AMPL_WIDTH),
		7033 => to_signed(20458, LUT_AMPL_WIDTH),
		7034 => to_signed(20460, LUT_AMPL_WIDTH),
		7035 => to_signed(20463, LUT_AMPL_WIDTH),
		7036 => to_signed(20465, LUT_AMPL_WIDTH),
		7037 => to_signed(20467, LUT_AMPL_WIDTH),
		7038 => to_signed(20470, LUT_AMPL_WIDTH),
		7039 => to_signed(20472, LUT_AMPL_WIDTH),
		7040 => to_signed(20475, LUT_AMPL_WIDTH),
		7041 => to_signed(20477, LUT_AMPL_WIDTH),
		7042 => to_signed(20480, LUT_AMPL_WIDTH),
		7043 => to_signed(20482, LUT_AMPL_WIDTH),
		7044 => to_signed(20485, LUT_AMPL_WIDTH),
		7045 => to_signed(20487, LUT_AMPL_WIDTH),
		7046 => to_signed(20489, LUT_AMPL_WIDTH),
		7047 => to_signed(20492, LUT_AMPL_WIDTH),
		7048 => to_signed(20494, LUT_AMPL_WIDTH),
		7049 => to_signed(20497, LUT_AMPL_WIDTH),
		7050 => to_signed(20499, LUT_AMPL_WIDTH),
		7051 => to_signed(20502, LUT_AMPL_WIDTH),
		7052 => to_signed(20504, LUT_AMPL_WIDTH),
		7053 => to_signed(20507, LUT_AMPL_WIDTH),
		7054 => to_signed(20509, LUT_AMPL_WIDTH),
		7055 => to_signed(20512, LUT_AMPL_WIDTH),
		7056 => to_signed(20514, LUT_AMPL_WIDTH),
		7057 => to_signed(20516, LUT_AMPL_WIDTH),
		7058 => to_signed(20519, LUT_AMPL_WIDTH),
		7059 => to_signed(20521, LUT_AMPL_WIDTH),
		7060 => to_signed(20524, LUT_AMPL_WIDTH),
		7061 => to_signed(20526, LUT_AMPL_WIDTH),
		7062 => to_signed(20529, LUT_AMPL_WIDTH),
		7063 => to_signed(20531, LUT_AMPL_WIDTH),
		7064 => to_signed(20534, LUT_AMPL_WIDTH),
		7065 => to_signed(20536, LUT_AMPL_WIDTH),
		7066 => to_signed(20538, LUT_AMPL_WIDTH),
		7067 => to_signed(20541, LUT_AMPL_WIDTH),
		7068 => to_signed(20543, LUT_AMPL_WIDTH),
		7069 => to_signed(20546, LUT_AMPL_WIDTH),
		7070 => to_signed(20548, LUT_AMPL_WIDTH),
		7071 => to_signed(20551, LUT_AMPL_WIDTH),
		7072 => to_signed(20553, LUT_AMPL_WIDTH),
		7073 => to_signed(20556, LUT_AMPL_WIDTH),
		7074 => to_signed(20558, LUT_AMPL_WIDTH),
		7075 => to_signed(20560, LUT_AMPL_WIDTH),
		7076 => to_signed(20563, LUT_AMPL_WIDTH),
		7077 => to_signed(20565, LUT_AMPL_WIDTH),
		7078 => to_signed(20568, LUT_AMPL_WIDTH),
		7079 => to_signed(20570, LUT_AMPL_WIDTH),
		7080 => to_signed(20573, LUT_AMPL_WIDTH),
		7081 => to_signed(20575, LUT_AMPL_WIDTH),
		7082 => to_signed(20578, LUT_AMPL_WIDTH),
		7083 => to_signed(20580, LUT_AMPL_WIDTH),
		7084 => to_signed(20583, LUT_AMPL_WIDTH),
		7085 => to_signed(20585, LUT_AMPL_WIDTH),
		7086 => to_signed(20587, LUT_AMPL_WIDTH),
		7087 => to_signed(20590, LUT_AMPL_WIDTH),
		7088 => to_signed(20592, LUT_AMPL_WIDTH),
		7089 => to_signed(20595, LUT_AMPL_WIDTH),
		7090 => to_signed(20597, LUT_AMPL_WIDTH),
		7091 => to_signed(20600, LUT_AMPL_WIDTH),
		7092 => to_signed(20602, LUT_AMPL_WIDTH),
		7093 => to_signed(20604, LUT_AMPL_WIDTH),
		7094 => to_signed(20607, LUT_AMPL_WIDTH),
		7095 => to_signed(20609, LUT_AMPL_WIDTH),
		7096 => to_signed(20612, LUT_AMPL_WIDTH),
		7097 => to_signed(20614, LUT_AMPL_WIDTH),
		7098 => to_signed(20617, LUT_AMPL_WIDTH),
		7099 => to_signed(20619, LUT_AMPL_WIDTH),
		7100 => to_signed(20622, LUT_AMPL_WIDTH),
		7101 => to_signed(20624, LUT_AMPL_WIDTH),
		7102 => to_signed(20626, LUT_AMPL_WIDTH),
		7103 => to_signed(20629, LUT_AMPL_WIDTH),
		7104 => to_signed(20631, LUT_AMPL_WIDTH),
		7105 => to_signed(20634, LUT_AMPL_WIDTH),
		7106 => to_signed(20636, LUT_AMPL_WIDTH),
		7107 => to_signed(20639, LUT_AMPL_WIDTH),
		7108 => to_signed(20641, LUT_AMPL_WIDTH),
		7109 => to_signed(20644, LUT_AMPL_WIDTH),
		7110 => to_signed(20646, LUT_AMPL_WIDTH),
		7111 => to_signed(20648, LUT_AMPL_WIDTH),
		7112 => to_signed(20651, LUT_AMPL_WIDTH),
		7113 => to_signed(20653, LUT_AMPL_WIDTH),
		7114 => to_signed(20656, LUT_AMPL_WIDTH),
		7115 => to_signed(20658, LUT_AMPL_WIDTH),
		7116 => to_signed(20661, LUT_AMPL_WIDTH),
		7117 => to_signed(20663, LUT_AMPL_WIDTH),
		7118 => to_signed(20666, LUT_AMPL_WIDTH),
		7119 => to_signed(20668, LUT_AMPL_WIDTH),
		7120 => to_signed(20670, LUT_AMPL_WIDTH),
		7121 => to_signed(20673, LUT_AMPL_WIDTH),
		7122 => to_signed(20675, LUT_AMPL_WIDTH),
		7123 => to_signed(20678, LUT_AMPL_WIDTH),
		7124 => to_signed(20680, LUT_AMPL_WIDTH),
		7125 => to_signed(20683, LUT_AMPL_WIDTH),
		7126 => to_signed(20685, LUT_AMPL_WIDTH),
		7127 => to_signed(20687, LUT_AMPL_WIDTH),
		7128 => to_signed(20690, LUT_AMPL_WIDTH),
		7129 => to_signed(20692, LUT_AMPL_WIDTH),
		7130 => to_signed(20695, LUT_AMPL_WIDTH),
		7131 => to_signed(20697, LUT_AMPL_WIDTH),
		7132 => to_signed(20700, LUT_AMPL_WIDTH),
		7133 => to_signed(20702, LUT_AMPL_WIDTH),
		7134 => to_signed(20704, LUT_AMPL_WIDTH),
		7135 => to_signed(20707, LUT_AMPL_WIDTH),
		7136 => to_signed(20709, LUT_AMPL_WIDTH),
		7137 => to_signed(20712, LUT_AMPL_WIDTH),
		7138 => to_signed(20714, LUT_AMPL_WIDTH),
		7139 => to_signed(20717, LUT_AMPL_WIDTH),
		7140 => to_signed(20719, LUT_AMPL_WIDTH),
		7141 => to_signed(20722, LUT_AMPL_WIDTH),
		7142 => to_signed(20724, LUT_AMPL_WIDTH),
		7143 => to_signed(20726, LUT_AMPL_WIDTH),
		7144 => to_signed(20729, LUT_AMPL_WIDTH),
		7145 => to_signed(20731, LUT_AMPL_WIDTH),
		7146 => to_signed(20734, LUT_AMPL_WIDTH),
		7147 => to_signed(20736, LUT_AMPL_WIDTH),
		7148 => to_signed(20739, LUT_AMPL_WIDTH),
		7149 => to_signed(20741, LUT_AMPL_WIDTH),
		7150 => to_signed(20743, LUT_AMPL_WIDTH),
		7151 => to_signed(20746, LUT_AMPL_WIDTH),
		7152 => to_signed(20748, LUT_AMPL_WIDTH),
		7153 => to_signed(20751, LUT_AMPL_WIDTH),
		7154 => to_signed(20753, LUT_AMPL_WIDTH),
		7155 => to_signed(20756, LUT_AMPL_WIDTH),
		7156 => to_signed(20758, LUT_AMPL_WIDTH),
		7157 => to_signed(20760, LUT_AMPL_WIDTH),
		7158 => to_signed(20763, LUT_AMPL_WIDTH),
		7159 => to_signed(20765, LUT_AMPL_WIDTH),
		7160 => to_signed(20768, LUT_AMPL_WIDTH),
		7161 => to_signed(20770, LUT_AMPL_WIDTH),
		7162 => to_signed(20773, LUT_AMPL_WIDTH),
		7163 => to_signed(20775, LUT_AMPL_WIDTH),
		7164 => to_signed(20777, LUT_AMPL_WIDTH),
		7165 => to_signed(20780, LUT_AMPL_WIDTH),
		7166 => to_signed(20782, LUT_AMPL_WIDTH),
		7167 => to_signed(20785, LUT_AMPL_WIDTH),
		7168 => to_signed(20787, LUT_AMPL_WIDTH),
		7169 => to_signed(20790, LUT_AMPL_WIDTH),
		7170 => to_signed(20792, LUT_AMPL_WIDTH),
		7171 => to_signed(20794, LUT_AMPL_WIDTH),
		7172 => to_signed(20797, LUT_AMPL_WIDTH),
		7173 => to_signed(20799, LUT_AMPL_WIDTH),
		7174 => to_signed(20802, LUT_AMPL_WIDTH),
		7175 => to_signed(20804, LUT_AMPL_WIDTH),
		7176 => to_signed(20807, LUT_AMPL_WIDTH),
		7177 => to_signed(20809, LUT_AMPL_WIDTH),
		7178 => to_signed(20811, LUT_AMPL_WIDTH),
		7179 => to_signed(20814, LUT_AMPL_WIDTH),
		7180 => to_signed(20816, LUT_AMPL_WIDTH),
		7181 => to_signed(20819, LUT_AMPL_WIDTH),
		7182 => to_signed(20821, LUT_AMPL_WIDTH),
		7183 => to_signed(20824, LUT_AMPL_WIDTH),
		7184 => to_signed(20826, LUT_AMPL_WIDTH),
		7185 => to_signed(20828, LUT_AMPL_WIDTH),
		7186 => to_signed(20831, LUT_AMPL_WIDTH),
		7187 => to_signed(20833, LUT_AMPL_WIDTH),
		7188 => to_signed(20836, LUT_AMPL_WIDTH),
		7189 => to_signed(20838, LUT_AMPL_WIDTH),
		7190 => to_signed(20841, LUT_AMPL_WIDTH),
		7191 => to_signed(20843, LUT_AMPL_WIDTH),
		7192 => to_signed(20845, LUT_AMPL_WIDTH),
		7193 => to_signed(20848, LUT_AMPL_WIDTH),
		7194 => to_signed(20850, LUT_AMPL_WIDTH),
		7195 => to_signed(20853, LUT_AMPL_WIDTH),
		7196 => to_signed(20855, LUT_AMPL_WIDTH),
		7197 => to_signed(20858, LUT_AMPL_WIDTH),
		7198 => to_signed(20860, LUT_AMPL_WIDTH),
		7199 => to_signed(20862, LUT_AMPL_WIDTH),
		7200 => to_signed(20865, LUT_AMPL_WIDTH),
		7201 => to_signed(20867, LUT_AMPL_WIDTH),
		7202 => to_signed(20870, LUT_AMPL_WIDTH),
		7203 => to_signed(20872, LUT_AMPL_WIDTH),
		7204 => to_signed(20874, LUT_AMPL_WIDTH),
		7205 => to_signed(20877, LUT_AMPL_WIDTH),
		7206 => to_signed(20879, LUT_AMPL_WIDTH),
		7207 => to_signed(20882, LUT_AMPL_WIDTH),
		7208 => to_signed(20884, LUT_AMPL_WIDTH),
		7209 => to_signed(20887, LUT_AMPL_WIDTH),
		7210 => to_signed(20889, LUT_AMPL_WIDTH),
		7211 => to_signed(20891, LUT_AMPL_WIDTH),
		7212 => to_signed(20894, LUT_AMPL_WIDTH),
		7213 => to_signed(20896, LUT_AMPL_WIDTH),
		7214 => to_signed(20899, LUT_AMPL_WIDTH),
		7215 => to_signed(20901, LUT_AMPL_WIDTH),
		7216 => to_signed(20904, LUT_AMPL_WIDTH),
		7217 => to_signed(20906, LUT_AMPL_WIDTH),
		7218 => to_signed(20908, LUT_AMPL_WIDTH),
		7219 => to_signed(20911, LUT_AMPL_WIDTH),
		7220 => to_signed(20913, LUT_AMPL_WIDTH),
		7221 => to_signed(20916, LUT_AMPL_WIDTH),
		7222 => to_signed(20918, LUT_AMPL_WIDTH),
		7223 => to_signed(20920, LUT_AMPL_WIDTH),
		7224 => to_signed(20923, LUT_AMPL_WIDTH),
		7225 => to_signed(20925, LUT_AMPL_WIDTH),
		7226 => to_signed(20928, LUT_AMPL_WIDTH),
		7227 => to_signed(20930, LUT_AMPL_WIDTH),
		7228 => to_signed(20933, LUT_AMPL_WIDTH),
		7229 => to_signed(20935, LUT_AMPL_WIDTH),
		7230 => to_signed(20937, LUT_AMPL_WIDTH),
		7231 => to_signed(20940, LUT_AMPL_WIDTH),
		7232 => to_signed(20942, LUT_AMPL_WIDTH),
		7233 => to_signed(20945, LUT_AMPL_WIDTH),
		7234 => to_signed(20947, LUT_AMPL_WIDTH),
		7235 => to_signed(20949, LUT_AMPL_WIDTH),
		7236 => to_signed(20952, LUT_AMPL_WIDTH),
		7237 => to_signed(20954, LUT_AMPL_WIDTH),
		7238 => to_signed(20957, LUT_AMPL_WIDTH),
		7239 => to_signed(20959, LUT_AMPL_WIDTH),
		7240 => to_signed(20962, LUT_AMPL_WIDTH),
		7241 => to_signed(20964, LUT_AMPL_WIDTH),
		7242 => to_signed(20966, LUT_AMPL_WIDTH),
		7243 => to_signed(20969, LUT_AMPL_WIDTH),
		7244 => to_signed(20971, LUT_AMPL_WIDTH),
		7245 => to_signed(20974, LUT_AMPL_WIDTH),
		7246 => to_signed(20976, LUT_AMPL_WIDTH),
		7247 => to_signed(20978, LUT_AMPL_WIDTH),
		7248 => to_signed(20981, LUT_AMPL_WIDTH),
		7249 => to_signed(20983, LUT_AMPL_WIDTH),
		7250 => to_signed(20986, LUT_AMPL_WIDTH),
		7251 => to_signed(20988, LUT_AMPL_WIDTH),
		7252 => to_signed(20990, LUT_AMPL_WIDTH),
		7253 => to_signed(20993, LUT_AMPL_WIDTH),
		7254 => to_signed(20995, LUT_AMPL_WIDTH),
		7255 => to_signed(20998, LUT_AMPL_WIDTH),
		7256 => to_signed(21000, LUT_AMPL_WIDTH),
		7257 => to_signed(21003, LUT_AMPL_WIDTH),
		7258 => to_signed(21005, LUT_AMPL_WIDTH),
		7259 => to_signed(21007, LUT_AMPL_WIDTH),
		7260 => to_signed(21010, LUT_AMPL_WIDTH),
		7261 => to_signed(21012, LUT_AMPL_WIDTH),
		7262 => to_signed(21015, LUT_AMPL_WIDTH),
		7263 => to_signed(21017, LUT_AMPL_WIDTH),
		7264 => to_signed(21019, LUT_AMPL_WIDTH),
		7265 => to_signed(21022, LUT_AMPL_WIDTH),
		7266 => to_signed(21024, LUT_AMPL_WIDTH),
		7267 => to_signed(21027, LUT_AMPL_WIDTH),
		7268 => to_signed(21029, LUT_AMPL_WIDTH),
		7269 => to_signed(21031, LUT_AMPL_WIDTH),
		7270 => to_signed(21034, LUT_AMPL_WIDTH),
		7271 => to_signed(21036, LUT_AMPL_WIDTH),
		7272 => to_signed(21039, LUT_AMPL_WIDTH),
		7273 => to_signed(21041, LUT_AMPL_WIDTH),
		7274 => to_signed(21043, LUT_AMPL_WIDTH),
		7275 => to_signed(21046, LUT_AMPL_WIDTH),
		7276 => to_signed(21048, LUT_AMPL_WIDTH),
		7277 => to_signed(21051, LUT_AMPL_WIDTH),
		7278 => to_signed(21053, LUT_AMPL_WIDTH),
		7279 => to_signed(21056, LUT_AMPL_WIDTH),
		7280 => to_signed(21058, LUT_AMPL_WIDTH),
		7281 => to_signed(21060, LUT_AMPL_WIDTH),
		7282 => to_signed(21063, LUT_AMPL_WIDTH),
		7283 => to_signed(21065, LUT_AMPL_WIDTH),
		7284 => to_signed(21068, LUT_AMPL_WIDTH),
		7285 => to_signed(21070, LUT_AMPL_WIDTH),
		7286 => to_signed(21072, LUT_AMPL_WIDTH),
		7287 => to_signed(21075, LUT_AMPL_WIDTH),
		7288 => to_signed(21077, LUT_AMPL_WIDTH),
		7289 => to_signed(21080, LUT_AMPL_WIDTH),
		7290 => to_signed(21082, LUT_AMPL_WIDTH),
		7291 => to_signed(21084, LUT_AMPL_WIDTH),
		7292 => to_signed(21087, LUT_AMPL_WIDTH),
		7293 => to_signed(21089, LUT_AMPL_WIDTH),
		7294 => to_signed(21092, LUT_AMPL_WIDTH),
		7295 => to_signed(21094, LUT_AMPL_WIDTH),
		7296 => to_signed(21096, LUT_AMPL_WIDTH),
		7297 => to_signed(21099, LUT_AMPL_WIDTH),
		7298 => to_signed(21101, LUT_AMPL_WIDTH),
		7299 => to_signed(21104, LUT_AMPL_WIDTH),
		7300 => to_signed(21106, LUT_AMPL_WIDTH),
		7301 => to_signed(21108, LUT_AMPL_WIDTH),
		7302 => to_signed(21111, LUT_AMPL_WIDTH),
		7303 => to_signed(21113, LUT_AMPL_WIDTH),
		7304 => to_signed(21116, LUT_AMPL_WIDTH),
		7305 => to_signed(21118, LUT_AMPL_WIDTH),
		7306 => to_signed(21120, LUT_AMPL_WIDTH),
		7307 => to_signed(21123, LUT_AMPL_WIDTH),
		7308 => to_signed(21125, LUT_AMPL_WIDTH),
		7309 => to_signed(21128, LUT_AMPL_WIDTH),
		7310 => to_signed(21130, LUT_AMPL_WIDTH),
		7311 => to_signed(21132, LUT_AMPL_WIDTH),
		7312 => to_signed(21135, LUT_AMPL_WIDTH),
		7313 => to_signed(21137, LUT_AMPL_WIDTH),
		7314 => to_signed(21140, LUT_AMPL_WIDTH),
		7315 => to_signed(21142, LUT_AMPL_WIDTH),
		7316 => to_signed(21144, LUT_AMPL_WIDTH),
		7317 => to_signed(21147, LUT_AMPL_WIDTH),
		7318 => to_signed(21149, LUT_AMPL_WIDTH),
		7319 => to_signed(21152, LUT_AMPL_WIDTH),
		7320 => to_signed(21154, LUT_AMPL_WIDTH),
		7321 => to_signed(21156, LUT_AMPL_WIDTH),
		7322 => to_signed(21159, LUT_AMPL_WIDTH),
		7323 => to_signed(21161, LUT_AMPL_WIDTH),
		7324 => to_signed(21164, LUT_AMPL_WIDTH),
		7325 => to_signed(21166, LUT_AMPL_WIDTH),
		7326 => to_signed(21168, LUT_AMPL_WIDTH),
		7327 => to_signed(21171, LUT_AMPL_WIDTH),
		7328 => to_signed(21173, LUT_AMPL_WIDTH),
		7329 => to_signed(21176, LUT_AMPL_WIDTH),
		7330 => to_signed(21178, LUT_AMPL_WIDTH),
		7331 => to_signed(21180, LUT_AMPL_WIDTH),
		7332 => to_signed(21183, LUT_AMPL_WIDTH),
		7333 => to_signed(21185, LUT_AMPL_WIDTH),
		7334 => to_signed(21188, LUT_AMPL_WIDTH),
		7335 => to_signed(21190, LUT_AMPL_WIDTH),
		7336 => to_signed(21192, LUT_AMPL_WIDTH),
		7337 => to_signed(21195, LUT_AMPL_WIDTH),
		7338 => to_signed(21197, LUT_AMPL_WIDTH),
		7339 => to_signed(21200, LUT_AMPL_WIDTH),
		7340 => to_signed(21202, LUT_AMPL_WIDTH),
		7341 => to_signed(21204, LUT_AMPL_WIDTH),
		7342 => to_signed(21207, LUT_AMPL_WIDTH),
		7343 => to_signed(21209, LUT_AMPL_WIDTH),
		7344 => to_signed(21212, LUT_AMPL_WIDTH),
		7345 => to_signed(21214, LUT_AMPL_WIDTH),
		7346 => to_signed(21216, LUT_AMPL_WIDTH),
		7347 => to_signed(21219, LUT_AMPL_WIDTH),
		7348 => to_signed(21221, LUT_AMPL_WIDTH),
		7349 => to_signed(21224, LUT_AMPL_WIDTH),
		7350 => to_signed(21226, LUT_AMPL_WIDTH),
		7351 => to_signed(21228, LUT_AMPL_WIDTH),
		7352 => to_signed(21231, LUT_AMPL_WIDTH),
		7353 => to_signed(21233, LUT_AMPL_WIDTH),
		7354 => to_signed(21236, LUT_AMPL_WIDTH),
		7355 => to_signed(21238, LUT_AMPL_WIDTH),
		7356 => to_signed(21240, LUT_AMPL_WIDTH),
		7357 => to_signed(21243, LUT_AMPL_WIDTH),
		7358 => to_signed(21245, LUT_AMPL_WIDTH),
		7359 => to_signed(21247, LUT_AMPL_WIDTH),
		7360 => to_signed(21250, LUT_AMPL_WIDTH),
		7361 => to_signed(21252, LUT_AMPL_WIDTH),
		7362 => to_signed(21255, LUT_AMPL_WIDTH),
		7363 => to_signed(21257, LUT_AMPL_WIDTH),
		7364 => to_signed(21259, LUT_AMPL_WIDTH),
		7365 => to_signed(21262, LUT_AMPL_WIDTH),
		7366 => to_signed(21264, LUT_AMPL_WIDTH),
		7367 => to_signed(21267, LUT_AMPL_WIDTH),
		7368 => to_signed(21269, LUT_AMPL_WIDTH),
		7369 => to_signed(21271, LUT_AMPL_WIDTH),
		7370 => to_signed(21274, LUT_AMPL_WIDTH),
		7371 => to_signed(21276, LUT_AMPL_WIDTH),
		7372 => to_signed(21279, LUT_AMPL_WIDTH),
		7373 => to_signed(21281, LUT_AMPL_WIDTH),
		7374 => to_signed(21283, LUT_AMPL_WIDTH),
		7375 => to_signed(21286, LUT_AMPL_WIDTH),
		7376 => to_signed(21288, LUT_AMPL_WIDTH),
		7377 => to_signed(21290, LUT_AMPL_WIDTH),
		7378 => to_signed(21293, LUT_AMPL_WIDTH),
		7379 => to_signed(21295, LUT_AMPL_WIDTH),
		7380 => to_signed(21298, LUT_AMPL_WIDTH),
		7381 => to_signed(21300, LUT_AMPL_WIDTH),
		7382 => to_signed(21302, LUT_AMPL_WIDTH),
		7383 => to_signed(21305, LUT_AMPL_WIDTH),
		7384 => to_signed(21307, LUT_AMPL_WIDTH),
		7385 => to_signed(21310, LUT_AMPL_WIDTH),
		7386 => to_signed(21312, LUT_AMPL_WIDTH),
		7387 => to_signed(21314, LUT_AMPL_WIDTH),
		7388 => to_signed(21317, LUT_AMPL_WIDTH),
		7389 => to_signed(21319, LUT_AMPL_WIDTH),
		7390 => to_signed(21322, LUT_AMPL_WIDTH),
		7391 => to_signed(21324, LUT_AMPL_WIDTH),
		7392 => to_signed(21326, LUT_AMPL_WIDTH),
		7393 => to_signed(21329, LUT_AMPL_WIDTH),
		7394 => to_signed(21331, LUT_AMPL_WIDTH),
		7395 => to_signed(21333, LUT_AMPL_WIDTH),
		7396 => to_signed(21336, LUT_AMPL_WIDTH),
		7397 => to_signed(21338, LUT_AMPL_WIDTH),
		7398 => to_signed(21341, LUT_AMPL_WIDTH),
		7399 => to_signed(21343, LUT_AMPL_WIDTH),
		7400 => to_signed(21345, LUT_AMPL_WIDTH),
		7401 => to_signed(21348, LUT_AMPL_WIDTH),
		7402 => to_signed(21350, LUT_AMPL_WIDTH),
		7403 => to_signed(21353, LUT_AMPL_WIDTH),
		7404 => to_signed(21355, LUT_AMPL_WIDTH),
		7405 => to_signed(21357, LUT_AMPL_WIDTH),
		7406 => to_signed(21360, LUT_AMPL_WIDTH),
		7407 => to_signed(21362, LUT_AMPL_WIDTH),
		7408 => to_signed(21364, LUT_AMPL_WIDTH),
		7409 => to_signed(21367, LUT_AMPL_WIDTH),
		7410 => to_signed(21369, LUT_AMPL_WIDTH),
		7411 => to_signed(21372, LUT_AMPL_WIDTH),
		7412 => to_signed(21374, LUT_AMPL_WIDTH),
		7413 => to_signed(21376, LUT_AMPL_WIDTH),
		7414 => to_signed(21379, LUT_AMPL_WIDTH),
		7415 => to_signed(21381, LUT_AMPL_WIDTH),
		7416 => to_signed(21383, LUT_AMPL_WIDTH),
		7417 => to_signed(21386, LUT_AMPL_WIDTH),
		7418 => to_signed(21388, LUT_AMPL_WIDTH),
		7419 => to_signed(21391, LUT_AMPL_WIDTH),
		7420 => to_signed(21393, LUT_AMPL_WIDTH),
		7421 => to_signed(21395, LUT_AMPL_WIDTH),
		7422 => to_signed(21398, LUT_AMPL_WIDTH),
		7423 => to_signed(21400, LUT_AMPL_WIDTH),
		7424 => to_signed(21403, LUT_AMPL_WIDTH),
		7425 => to_signed(21405, LUT_AMPL_WIDTH),
		7426 => to_signed(21407, LUT_AMPL_WIDTH),
		7427 => to_signed(21410, LUT_AMPL_WIDTH),
		7428 => to_signed(21412, LUT_AMPL_WIDTH),
		7429 => to_signed(21414, LUT_AMPL_WIDTH),
		7430 => to_signed(21417, LUT_AMPL_WIDTH),
		7431 => to_signed(21419, LUT_AMPL_WIDTH),
		7432 => to_signed(21422, LUT_AMPL_WIDTH),
		7433 => to_signed(21424, LUT_AMPL_WIDTH),
		7434 => to_signed(21426, LUT_AMPL_WIDTH),
		7435 => to_signed(21429, LUT_AMPL_WIDTH),
		7436 => to_signed(21431, LUT_AMPL_WIDTH),
		7437 => to_signed(21433, LUT_AMPL_WIDTH),
		7438 => to_signed(21436, LUT_AMPL_WIDTH),
		7439 => to_signed(21438, LUT_AMPL_WIDTH),
		7440 => to_signed(21441, LUT_AMPL_WIDTH),
		7441 => to_signed(21443, LUT_AMPL_WIDTH),
		7442 => to_signed(21445, LUT_AMPL_WIDTH),
		7443 => to_signed(21448, LUT_AMPL_WIDTH),
		7444 => to_signed(21450, LUT_AMPL_WIDTH),
		7445 => to_signed(21452, LUT_AMPL_WIDTH),
		7446 => to_signed(21455, LUT_AMPL_WIDTH),
		7447 => to_signed(21457, LUT_AMPL_WIDTH),
		7448 => to_signed(21460, LUT_AMPL_WIDTH),
		7449 => to_signed(21462, LUT_AMPL_WIDTH),
		7450 => to_signed(21464, LUT_AMPL_WIDTH),
		7451 => to_signed(21467, LUT_AMPL_WIDTH),
		7452 => to_signed(21469, LUT_AMPL_WIDTH),
		7453 => to_signed(21471, LUT_AMPL_WIDTH),
		7454 => to_signed(21474, LUT_AMPL_WIDTH),
		7455 => to_signed(21476, LUT_AMPL_WIDTH),
		7456 => to_signed(21479, LUT_AMPL_WIDTH),
		7457 => to_signed(21481, LUT_AMPL_WIDTH),
		7458 => to_signed(21483, LUT_AMPL_WIDTH),
		7459 => to_signed(21486, LUT_AMPL_WIDTH),
		7460 => to_signed(21488, LUT_AMPL_WIDTH),
		7461 => to_signed(21490, LUT_AMPL_WIDTH),
		7462 => to_signed(21493, LUT_AMPL_WIDTH),
		7463 => to_signed(21495, LUT_AMPL_WIDTH),
		7464 => to_signed(21498, LUT_AMPL_WIDTH),
		7465 => to_signed(21500, LUT_AMPL_WIDTH),
		7466 => to_signed(21502, LUT_AMPL_WIDTH),
		7467 => to_signed(21505, LUT_AMPL_WIDTH),
		7468 => to_signed(21507, LUT_AMPL_WIDTH),
		7469 => to_signed(21509, LUT_AMPL_WIDTH),
		7470 => to_signed(21512, LUT_AMPL_WIDTH),
		7471 => to_signed(21514, LUT_AMPL_WIDTH),
		7472 => to_signed(21516, LUT_AMPL_WIDTH),
		7473 => to_signed(21519, LUT_AMPL_WIDTH),
		7474 => to_signed(21521, LUT_AMPL_WIDTH),
		7475 => to_signed(21524, LUT_AMPL_WIDTH),
		7476 => to_signed(21526, LUT_AMPL_WIDTH),
		7477 => to_signed(21528, LUT_AMPL_WIDTH),
		7478 => to_signed(21531, LUT_AMPL_WIDTH),
		7479 => to_signed(21533, LUT_AMPL_WIDTH),
		7480 => to_signed(21535, LUT_AMPL_WIDTH),
		7481 => to_signed(21538, LUT_AMPL_WIDTH),
		7482 => to_signed(21540, LUT_AMPL_WIDTH),
		7483 => to_signed(21543, LUT_AMPL_WIDTH),
		7484 => to_signed(21545, LUT_AMPL_WIDTH),
		7485 => to_signed(21547, LUT_AMPL_WIDTH),
		7486 => to_signed(21550, LUT_AMPL_WIDTH),
		7487 => to_signed(21552, LUT_AMPL_WIDTH),
		7488 => to_signed(21554, LUT_AMPL_WIDTH),
		7489 => to_signed(21557, LUT_AMPL_WIDTH),
		7490 => to_signed(21559, LUT_AMPL_WIDTH),
		7491 => to_signed(21561, LUT_AMPL_WIDTH),
		7492 => to_signed(21564, LUT_AMPL_WIDTH),
		7493 => to_signed(21566, LUT_AMPL_WIDTH),
		7494 => to_signed(21569, LUT_AMPL_WIDTH),
		7495 => to_signed(21571, LUT_AMPL_WIDTH),
		7496 => to_signed(21573, LUT_AMPL_WIDTH),
		7497 => to_signed(21576, LUT_AMPL_WIDTH),
		7498 => to_signed(21578, LUT_AMPL_WIDTH),
		7499 => to_signed(21580, LUT_AMPL_WIDTH),
		7500 => to_signed(21583, LUT_AMPL_WIDTH),
		7501 => to_signed(21585, LUT_AMPL_WIDTH),
		7502 => to_signed(21587, LUT_AMPL_WIDTH),
		7503 => to_signed(21590, LUT_AMPL_WIDTH),
		7504 => to_signed(21592, LUT_AMPL_WIDTH),
		7505 => to_signed(21595, LUT_AMPL_WIDTH),
		7506 => to_signed(21597, LUT_AMPL_WIDTH),
		7507 => to_signed(21599, LUT_AMPL_WIDTH),
		7508 => to_signed(21602, LUT_AMPL_WIDTH),
		7509 => to_signed(21604, LUT_AMPL_WIDTH),
		7510 => to_signed(21606, LUT_AMPL_WIDTH),
		7511 => to_signed(21609, LUT_AMPL_WIDTH),
		7512 => to_signed(21611, LUT_AMPL_WIDTH),
		7513 => to_signed(21613, LUT_AMPL_WIDTH),
		7514 => to_signed(21616, LUT_AMPL_WIDTH),
		7515 => to_signed(21618, LUT_AMPL_WIDTH),
		7516 => to_signed(21621, LUT_AMPL_WIDTH),
		7517 => to_signed(21623, LUT_AMPL_WIDTH),
		7518 => to_signed(21625, LUT_AMPL_WIDTH),
		7519 => to_signed(21628, LUT_AMPL_WIDTH),
		7520 => to_signed(21630, LUT_AMPL_WIDTH),
		7521 => to_signed(21632, LUT_AMPL_WIDTH),
		7522 => to_signed(21635, LUT_AMPL_WIDTH),
		7523 => to_signed(21637, LUT_AMPL_WIDTH),
		7524 => to_signed(21639, LUT_AMPL_WIDTH),
		7525 => to_signed(21642, LUT_AMPL_WIDTH),
		7526 => to_signed(21644, LUT_AMPL_WIDTH),
		7527 => to_signed(21646, LUT_AMPL_WIDTH),
		7528 => to_signed(21649, LUT_AMPL_WIDTH),
		7529 => to_signed(21651, LUT_AMPL_WIDTH),
		7530 => to_signed(21654, LUT_AMPL_WIDTH),
		7531 => to_signed(21656, LUT_AMPL_WIDTH),
		7532 => to_signed(21658, LUT_AMPL_WIDTH),
		7533 => to_signed(21661, LUT_AMPL_WIDTH),
		7534 => to_signed(21663, LUT_AMPL_WIDTH),
		7535 => to_signed(21665, LUT_AMPL_WIDTH),
		7536 => to_signed(21668, LUT_AMPL_WIDTH),
		7537 => to_signed(21670, LUT_AMPL_WIDTH),
		7538 => to_signed(21672, LUT_AMPL_WIDTH),
		7539 => to_signed(21675, LUT_AMPL_WIDTH),
		7540 => to_signed(21677, LUT_AMPL_WIDTH),
		7541 => to_signed(21679, LUT_AMPL_WIDTH),
		7542 => to_signed(21682, LUT_AMPL_WIDTH),
		7543 => to_signed(21684, LUT_AMPL_WIDTH),
		7544 => to_signed(21687, LUT_AMPL_WIDTH),
		7545 => to_signed(21689, LUT_AMPL_WIDTH),
		7546 => to_signed(21691, LUT_AMPL_WIDTH),
		7547 => to_signed(21694, LUT_AMPL_WIDTH),
		7548 => to_signed(21696, LUT_AMPL_WIDTH),
		7549 => to_signed(21698, LUT_AMPL_WIDTH),
		7550 => to_signed(21701, LUT_AMPL_WIDTH),
		7551 => to_signed(21703, LUT_AMPL_WIDTH),
		7552 => to_signed(21705, LUT_AMPL_WIDTH),
		7553 => to_signed(21708, LUT_AMPL_WIDTH),
		7554 => to_signed(21710, LUT_AMPL_WIDTH),
		7555 => to_signed(21712, LUT_AMPL_WIDTH),
		7556 => to_signed(21715, LUT_AMPL_WIDTH),
		7557 => to_signed(21717, LUT_AMPL_WIDTH),
		7558 => to_signed(21719, LUT_AMPL_WIDTH),
		7559 => to_signed(21722, LUT_AMPL_WIDTH),
		7560 => to_signed(21724, LUT_AMPL_WIDTH),
		7561 => to_signed(21727, LUT_AMPL_WIDTH),
		7562 => to_signed(21729, LUT_AMPL_WIDTH),
		7563 => to_signed(21731, LUT_AMPL_WIDTH),
		7564 => to_signed(21734, LUT_AMPL_WIDTH),
		7565 => to_signed(21736, LUT_AMPL_WIDTH),
		7566 => to_signed(21738, LUT_AMPL_WIDTH),
		7567 => to_signed(21741, LUT_AMPL_WIDTH),
		7568 => to_signed(21743, LUT_AMPL_WIDTH),
		7569 => to_signed(21745, LUT_AMPL_WIDTH),
		7570 => to_signed(21748, LUT_AMPL_WIDTH),
		7571 => to_signed(21750, LUT_AMPL_WIDTH),
		7572 => to_signed(21752, LUT_AMPL_WIDTH),
		7573 => to_signed(21755, LUT_AMPL_WIDTH),
		7574 => to_signed(21757, LUT_AMPL_WIDTH),
		7575 => to_signed(21759, LUT_AMPL_WIDTH),
		7576 => to_signed(21762, LUT_AMPL_WIDTH),
		7577 => to_signed(21764, LUT_AMPL_WIDTH),
		7578 => to_signed(21766, LUT_AMPL_WIDTH),
		7579 => to_signed(21769, LUT_AMPL_WIDTH),
		7580 => to_signed(21771, LUT_AMPL_WIDTH),
		7581 => to_signed(21774, LUT_AMPL_WIDTH),
		7582 => to_signed(21776, LUT_AMPL_WIDTH),
		7583 => to_signed(21778, LUT_AMPL_WIDTH),
		7584 => to_signed(21781, LUT_AMPL_WIDTH),
		7585 => to_signed(21783, LUT_AMPL_WIDTH),
		7586 => to_signed(21785, LUT_AMPL_WIDTH),
		7587 => to_signed(21788, LUT_AMPL_WIDTH),
		7588 => to_signed(21790, LUT_AMPL_WIDTH),
		7589 => to_signed(21792, LUT_AMPL_WIDTH),
		7590 => to_signed(21795, LUT_AMPL_WIDTH),
		7591 => to_signed(21797, LUT_AMPL_WIDTH),
		7592 => to_signed(21799, LUT_AMPL_WIDTH),
		7593 => to_signed(21802, LUT_AMPL_WIDTH),
		7594 => to_signed(21804, LUT_AMPL_WIDTH),
		7595 => to_signed(21806, LUT_AMPL_WIDTH),
		7596 => to_signed(21809, LUT_AMPL_WIDTH),
		7597 => to_signed(21811, LUT_AMPL_WIDTH),
		7598 => to_signed(21813, LUT_AMPL_WIDTH),
		7599 => to_signed(21816, LUT_AMPL_WIDTH),
		7600 => to_signed(21818, LUT_AMPL_WIDTH),
		7601 => to_signed(21820, LUT_AMPL_WIDTH),
		7602 => to_signed(21823, LUT_AMPL_WIDTH),
		7603 => to_signed(21825, LUT_AMPL_WIDTH),
		7604 => to_signed(21827, LUT_AMPL_WIDTH),
		7605 => to_signed(21830, LUT_AMPL_WIDTH),
		7606 => to_signed(21832, LUT_AMPL_WIDTH),
		7607 => to_signed(21835, LUT_AMPL_WIDTH),
		7608 => to_signed(21837, LUT_AMPL_WIDTH),
		7609 => to_signed(21839, LUT_AMPL_WIDTH),
		7610 => to_signed(21842, LUT_AMPL_WIDTH),
		7611 => to_signed(21844, LUT_AMPL_WIDTH),
		7612 => to_signed(21846, LUT_AMPL_WIDTH),
		7613 => to_signed(21849, LUT_AMPL_WIDTH),
		7614 => to_signed(21851, LUT_AMPL_WIDTH),
		7615 => to_signed(21853, LUT_AMPL_WIDTH),
		7616 => to_signed(21856, LUT_AMPL_WIDTH),
		7617 => to_signed(21858, LUT_AMPL_WIDTH),
		7618 => to_signed(21860, LUT_AMPL_WIDTH),
		7619 => to_signed(21863, LUT_AMPL_WIDTH),
		7620 => to_signed(21865, LUT_AMPL_WIDTH),
		7621 => to_signed(21867, LUT_AMPL_WIDTH),
		7622 => to_signed(21870, LUT_AMPL_WIDTH),
		7623 => to_signed(21872, LUT_AMPL_WIDTH),
		7624 => to_signed(21874, LUT_AMPL_WIDTH),
		7625 => to_signed(21877, LUT_AMPL_WIDTH),
		7626 => to_signed(21879, LUT_AMPL_WIDTH),
		7627 => to_signed(21881, LUT_AMPL_WIDTH),
		7628 => to_signed(21884, LUT_AMPL_WIDTH),
		7629 => to_signed(21886, LUT_AMPL_WIDTH),
		7630 => to_signed(21888, LUT_AMPL_WIDTH),
		7631 => to_signed(21891, LUT_AMPL_WIDTH),
		7632 => to_signed(21893, LUT_AMPL_WIDTH),
		7633 => to_signed(21895, LUT_AMPL_WIDTH),
		7634 => to_signed(21898, LUT_AMPL_WIDTH),
		7635 => to_signed(21900, LUT_AMPL_WIDTH),
		7636 => to_signed(21902, LUT_AMPL_WIDTH),
		7637 => to_signed(21905, LUT_AMPL_WIDTH),
		7638 => to_signed(21907, LUT_AMPL_WIDTH),
		7639 => to_signed(21909, LUT_AMPL_WIDTH),
		7640 => to_signed(21912, LUT_AMPL_WIDTH),
		7641 => to_signed(21914, LUT_AMPL_WIDTH),
		7642 => to_signed(21916, LUT_AMPL_WIDTH),
		7643 => to_signed(21919, LUT_AMPL_WIDTH),
		7644 => to_signed(21921, LUT_AMPL_WIDTH),
		7645 => to_signed(21923, LUT_AMPL_WIDTH),
		7646 => to_signed(21926, LUT_AMPL_WIDTH),
		7647 => to_signed(21928, LUT_AMPL_WIDTH),
		7648 => to_signed(21930, LUT_AMPL_WIDTH),
		7649 => to_signed(21933, LUT_AMPL_WIDTH),
		7650 => to_signed(21935, LUT_AMPL_WIDTH),
		7651 => to_signed(21937, LUT_AMPL_WIDTH),
		7652 => to_signed(21940, LUT_AMPL_WIDTH),
		7653 => to_signed(21942, LUT_AMPL_WIDTH),
		7654 => to_signed(21944, LUT_AMPL_WIDTH),
		7655 => to_signed(21947, LUT_AMPL_WIDTH),
		7656 => to_signed(21949, LUT_AMPL_WIDTH),
		7657 => to_signed(21951, LUT_AMPL_WIDTH),
		7658 => to_signed(21954, LUT_AMPL_WIDTH),
		7659 => to_signed(21956, LUT_AMPL_WIDTH),
		7660 => to_signed(21958, LUT_AMPL_WIDTH),
		7661 => to_signed(21961, LUT_AMPL_WIDTH),
		7662 => to_signed(21963, LUT_AMPL_WIDTH),
		7663 => to_signed(21965, LUT_AMPL_WIDTH),
		7664 => to_signed(21968, LUT_AMPL_WIDTH),
		7665 => to_signed(21970, LUT_AMPL_WIDTH),
		7666 => to_signed(21972, LUT_AMPL_WIDTH),
		7667 => to_signed(21975, LUT_AMPL_WIDTH),
		7668 => to_signed(21977, LUT_AMPL_WIDTH),
		7669 => to_signed(21979, LUT_AMPL_WIDTH),
		7670 => to_signed(21982, LUT_AMPL_WIDTH),
		7671 => to_signed(21984, LUT_AMPL_WIDTH),
		7672 => to_signed(21986, LUT_AMPL_WIDTH),
		7673 => to_signed(21989, LUT_AMPL_WIDTH),
		7674 => to_signed(21991, LUT_AMPL_WIDTH),
		7675 => to_signed(21993, LUT_AMPL_WIDTH),
		7676 => to_signed(21996, LUT_AMPL_WIDTH),
		7677 => to_signed(21998, LUT_AMPL_WIDTH),
		7678 => to_signed(22000, LUT_AMPL_WIDTH),
		7679 => to_signed(22003, LUT_AMPL_WIDTH),
		7680 => to_signed(22005, LUT_AMPL_WIDTH),
		7681 => to_signed(22007, LUT_AMPL_WIDTH),
		7682 => to_signed(22010, LUT_AMPL_WIDTH),
		7683 => to_signed(22012, LUT_AMPL_WIDTH),
		7684 => to_signed(22014, LUT_AMPL_WIDTH),
		7685 => to_signed(22017, LUT_AMPL_WIDTH),
		7686 => to_signed(22019, LUT_AMPL_WIDTH),
		7687 => to_signed(22021, LUT_AMPL_WIDTH),
		7688 => to_signed(22024, LUT_AMPL_WIDTH),
		7689 => to_signed(22026, LUT_AMPL_WIDTH),
		7690 => to_signed(22028, LUT_AMPL_WIDTH),
		7691 => to_signed(22031, LUT_AMPL_WIDTH),
		7692 => to_signed(22033, LUT_AMPL_WIDTH),
		7693 => to_signed(22035, LUT_AMPL_WIDTH),
		7694 => to_signed(22038, LUT_AMPL_WIDTH),
		7695 => to_signed(22040, LUT_AMPL_WIDTH),
		7696 => to_signed(22042, LUT_AMPL_WIDTH),
		7697 => to_signed(22045, LUT_AMPL_WIDTH),
		7698 => to_signed(22047, LUT_AMPL_WIDTH),
		7699 => to_signed(22049, LUT_AMPL_WIDTH),
		7700 => to_signed(22051, LUT_AMPL_WIDTH),
		7701 => to_signed(22054, LUT_AMPL_WIDTH),
		7702 => to_signed(22056, LUT_AMPL_WIDTH),
		7703 => to_signed(22058, LUT_AMPL_WIDTH),
		7704 => to_signed(22061, LUT_AMPL_WIDTH),
		7705 => to_signed(22063, LUT_AMPL_WIDTH),
		7706 => to_signed(22065, LUT_AMPL_WIDTH),
		7707 => to_signed(22068, LUT_AMPL_WIDTH),
		7708 => to_signed(22070, LUT_AMPL_WIDTH),
		7709 => to_signed(22072, LUT_AMPL_WIDTH),
		7710 => to_signed(22075, LUT_AMPL_WIDTH),
		7711 => to_signed(22077, LUT_AMPL_WIDTH),
		7712 => to_signed(22079, LUT_AMPL_WIDTH),
		7713 => to_signed(22082, LUT_AMPL_WIDTH),
		7714 => to_signed(22084, LUT_AMPL_WIDTH),
		7715 => to_signed(22086, LUT_AMPL_WIDTH),
		7716 => to_signed(22089, LUT_AMPL_WIDTH),
		7717 => to_signed(22091, LUT_AMPL_WIDTH),
		7718 => to_signed(22093, LUT_AMPL_WIDTH),
		7719 => to_signed(22096, LUT_AMPL_WIDTH),
		7720 => to_signed(22098, LUT_AMPL_WIDTH),
		7721 => to_signed(22100, LUT_AMPL_WIDTH),
		7722 => to_signed(22103, LUT_AMPL_WIDTH),
		7723 => to_signed(22105, LUT_AMPL_WIDTH),
		7724 => to_signed(22107, LUT_AMPL_WIDTH),
		7725 => to_signed(22110, LUT_AMPL_WIDTH),
		7726 => to_signed(22112, LUT_AMPL_WIDTH),
		7727 => to_signed(22114, LUT_AMPL_WIDTH),
		7728 => to_signed(22116, LUT_AMPL_WIDTH),
		7729 => to_signed(22119, LUT_AMPL_WIDTH),
		7730 => to_signed(22121, LUT_AMPL_WIDTH),
		7731 => to_signed(22123, LUT_AMPL_WIDTH),
		7732 => to_signed(22126, LUT_AMPL_WIDTH),
		7733 => to_signed(22128, LUT_AMPL_WIDTH),
		7734 => to_signed(22130, LUT_AMPL_WIDTH),
		7735 => to_signed(22133, LUT_AMPL_WIDTH),
		7736 => to_signed(22135, LUT_AMPL_WIDTH),
		7737 => to_signed(22137, LUT_AMPL_WIDTH),
		7738 => to_signed(22140, LUT_AMPL_WIDTH),
		7739 => to_signed(22142, LUT_AMPL_WIDTH),
		7740 => to_signed(22144, LUT_AMPL_WIDTH),
		7741 => to_signed(22147, LUT_AMPL_WIDTH),
		7742 => to_signed(22149, LUT_AMPL_WIDTH),
		7743 => to_signed(22151, LUT_AMPL_WIDTH),
		7744 => to_signed(22154, LUT_AMPL_WIDTH),
		7745 => to_signed(22156, LUT_AMPL_WIDTH),
		7746 => to_signed(22158, LUT_AMPL_WIDTH),
		7747 => to_signed(22160, LUT_AMPL_WIDTH),
		7748 => to_signed(22163, LUT_AMPL_WIDTH),
		7749 => to_signed(22165, LUT_AMPL_WIDTH),
		7750 => to_signed(22167, LUT_AMPL_WIDTH),
		7751 => to_signed(22170, LUT_AMPL_WIDTH),
		7752 => to_signed(22172, LUT_AMPL_WIDTH),
		7753 => to_signed(22174, LUT_AMPL_WIDTH),
		7754 => to_signed(22177, LUT_AMPL_WIDTH),
		7755 => to_signed(22179, LUT_AMPL_WIDTH),
		7756 => to_signed(22181, LUT_AMPL_WIDTH),
		7757 => to_signed(22184, LUT_AMPL_WIDTH),
		7758 => to_signed(22186, LUT_AMPL_WIDTH),
		7759 => to_signed(22188, LUT_AMPL_WIDTH),
		7760 => to_signed(22191, LUT_AMPL_WIDTH),
		7761 => to_signed(22193, LUT_AMPL_WIDTH),
		7762 => to_signed(22195, LUT_AMPL_WIDTH),
		7763 => to_signed(22197, LUT_AMPL_WIDTH),
		7764 => to_signed(22200, LUT_AMPL_WIDTH),
		7765 => to_signed(22202, LUT_AMPL_WIDTH),
		7766 => to_signed(22204, LUT_AMPL_WIDTH),
		7767 => to_signed(22207, LUT_AMPL_WIDTH),
		7768 => to_signed(22209, LUT_AMPL_WIDTH),
		7769 => to_signed(22211, LUT_AMPL_WIDTH),
		7770 => to_signed(22214, LUT_AMPL_WIDTH),
		7771 => to_signed(22216, LUT_AMPL_WIDTH),
		7772 => to_signed(22218, LUT_AMPL_WIDTH),
		7773 => to_signed(22221, LUT_AMPL_WIDTH),
		7774 => to_signed(22223, LUT_AMPL_WIDTH),
		7775 => to_signed(22225, LUT_AMPL_WIDTH),
		7776 => to_signed(22227, LUT_AMPL_WIDTH),
		7777 => to_signed(22230, LUT_AMPL_WIDTH),
		7778 => to_signed(22232, LUT_AMPL_WIDTH),
		7779 => to_signed(22234, LUT_AMPL_WIDTH),
		7780 => to_signed(22237, LUT_AMPL_WIDTH),
		7781 => to_signed(22239, LUT_AMPL_WIDTH),
		7782 => to_signed(22241, LUT_AMPL_WIDTH),
		7783 => to_signed(22244, LUT_AMPL_WIDTH),
		7784 => to_signed(22246, LUT_AMPL_WIDTH),
		7785 => to_signed(22248, LUT_AMPL_WIDTH),
		7786 => to_signed(22251, LUT_AMPL_WIDTH),
		7787 => to_signed(22253, LUT_AMPL_WIDTH),
		7788 => to_signed(22255, LUT_AMPL_WIDTH),
		7789 => to_signed(22257, LUT_AMPL_WIDTH),
		7790 => to_signed(22260, LUT_AMPL_WIDTH),
		7791 => to_signed(22262, LUT_AMPL_WIDTH),
		7792 => to_signed(22264, LUT_AMPL_WIDTH),
		7793 => to_signed(22267, LUT_AMPL_WIDTH),
		7794 => to_signed(22269, LUT_AMPL_WIDTH),
		7795 => to_signed(22271, LUT_AMPL_WIDTH),
		7796 => to_signed(22274, LUT_AMPL_WIDTH),
		7797 => to_signed(22276, LUT_AMPL_WIDTH),
		7798 => to_signed(22278, LUT_AMPL_WIDTH),
		7799 => to_signed(22281, LUT_AMPL_WIDTH),
		7800 => to_signed(22283, LUT_AMPL_WIDTH),
		7801 => to_signed(22285, LUT_AMPL_WIDTH),
		7802 => to_signed(22287, LUT_AMPL_WIDTH),
		7803 => to_signed(22290, LUT_AMPL_WIDTH),
		7804 => to_signed(22292, LUT_AMPL_WIDTH),
		7805 => to_signed(22294, LUT_AMPL_WIDTH),
		7806 => to_signed(22297, LUT_AMPL_WIDTH),
		7807 => to_signed(22299, LUT_AMPL_WIDTH),
		7808 => to_signed(22301, LUT_AMPL_WIDTH),
		7809 => to_signed(22304, LUT_AMPL_WIDTH),
		7810 => to_signed(22306, LUT_AMPL_WIDTH),
		7811 => to_signed(22308, LUT_AMPL_WIDTH),
		7812 => to_signed(22310, LUT_AMPL_WIDTH),
		7813 => to_signed(22313, LUT_AMPL_WIDTH),
		7814 => to_signed(22315, LUT_AMPL_WIDTH),
		7815 => to_signed(22317, LUT_AMPL_WIDTH),
		7816 => to_signed(22320, LUT_AMPL_WIDTH),
		7817 => to_signed(22322, LUT_AMPL_WIDTH),
		7818 => to_signed(22324, LUT_AMPL_WIDTH),
		7819 => to_signed(22327, LUT_AMPL_WIDTH),
		7820 => to_signed(22329, LUT_AMPL_WIDTH),
		7821 => to_signed(22331, LUT_AMPL_WIDTH),
		7822 => to_signed(22333, LUT_AMPL_WIDTH),
		7823 => to_signed(22336, LUT_AMPL_WIDTH),
		7824 => to_signed(22338, LUT_AMPL_WIDTH),
		7825 => to_signed(22340, LUT_AMPL_WIDTH),
		7826 => to_signed(22343, LUT_AMPL_WIDTH),
		7827 => to_signed(22345, LUT_AMPL_WIDTH),
		7828 => to_signed(22347, LUT_AMPL_WIDTH),
		7829 => to_signed(22350, LUT_AMPL_WIDTH),
		7830 => to_signed(22352, LUT_AMPL_WIDTH),
		7831 => to_signed(22354, LUT_AMPL_WIDTH),
		7832 => to_signed(22356, LUT_AMPL_WIDTH),
		7833 => to_signed(22359, LUT_AMPL_WIDTH),
		7834 => to_signed(22361, LUT_AMPL_WIDTH),
		7835 => to_signed(22363, LUT_AMPL_WIDTH),
		7836 => to_signed(22366, LUT_AMPL_WIDTH),
		7837 => to_signed(22368, LUT_AMPL_WIDTH),
		7838 => to_signed(22370, LUT_AMPL_WIDTH),
		7839 => to_signed(22373, LUT_AMPL_WIDTH),
		7840 => to_signed(22375, LUT_AMPL_WIDTH),
		7841 => to_signed(22377, LUT_AMPL_WIDTH),
		7842 => to_signed(22379, LUT_AMPL_WIDTH),
		7843 => to_signed(22382, LUT_AMPL_WIDTH),
		7844 => to_signed(22384, LUT_AMPL_WIDTH),
		7845 => to_signed(22386, LUT_AMPL_WIDTH),
		7846 => to_signed(22389, LUT_AMPL_WIDTH),
		7847 => to_signed(22391, LUT_AMPL_WIDTH),
		7848 => to_signed(22393, LUT_AMPL_WIDTH),
		7849 => to_signed(22395, LUT_AMPL_WIDTH),
		7850 => to_signed(22398, LUT_AMPL_WIDTH),
		7851 => to_signed(22400, LUT_AMPL_WIDTH),
		7852 => to_signed(22402, LUT_AMPL_WIDTH),
		7853 => to_signed(22405, LUT_AMPL_WIDTH),
		7854 => to_signed(22407, LUT_AMPL_WIDTH),
		7855 => to_signed(22409, LUT_AMPL_WIDTH),
		7856 => to_signed(22411, LUT_AMPL_WIDTH),
		7857 => to_signed(22414, LUT_AMPL_WIDTH),
		7858 => to_signed(22416, LUT_AMPL_WIDTH),
		7859 => to_signed(22418, LUT_AMPL_WIDTH),
		7860 => to_signed(22421, LUT_AMPL_WIDTH),
		7861 => to_signed(22423, LUT_AMPL_WIDTH),
		7862 => to_signed(22425, LUT_AMPL_WIDTH),
		7863 => to_signed(22428, LUT_AMPL_WIDTH),
		7864 => to_signed(22430, LUT_AMPL_WIDTH),
		7865 => to_signed(22432, LUT_AMPL_WIDTH),
		7866 => to_signed(22434, LUT_AMPL_WIDTH),
		7867 => to_signed(22437, LUT_AMPL_WIDTH),
		7868 => to_signed(22439, LUT_AMPL_WIDTH),
		7869 => to_signed(22441, LUT_AMPL_WIDTH),
		7870 => to_signed(22444, LUT_AMPL_WIDTH),
		7871 => to_signed(22446, LUT_AMPL_WIDTH),
		7872 => to_signed(22448, LUT_AMPL_WIDTH),
		7873 => to_signed(22450, LUT_AMPL_WIDTH),
		7874 => to_signed(22453, LUT_AMPL_WIDTH),
		7875 => to_signed(22455, LUT_AMPL_WIDTH),
		7876 => to_signed(22457, LUT_AMPL_WIDTH),
		7877 => to_signed(22460, LUT_AMPL_WIDTH),
		7878 => to_signed(22462, LUT_AMPL_WIDTH),
		7879 => to_signed(22464, LUT_AMPL_WIDTH),
		7880 => to_signed(22466, LUT_AMPL_WIDTH),
		7881 => to_signed(22469, LUT_AMPL_WIDTH),
		7882 => to_signed(22471, LUT_AMPL_WIDTH),
		7883 => to_signed(22473, LUT_AMPL_WIDTH),
		7884 => to_signed(22476, LUT_AMPL_WIDTH),
		7885 => to_signed(22478, LUT_AMPL_WIDTH),
		7886 => to_signed(22480, LUT_AMPL_WIDTH),
		7887 => to_signed(22482, LUT_AMPL_WIDTH),
		7888 => to_signed(22485, LUT_AMPL_WIDTH),
		7889 => to_signed(22487, LUT_AMPL_WIDTH),
		7890 => to_signed(22489, LUT_AMPL_WIDTH),
		7891 => to_signed(22492, LUT_AMPL_WIDTH),
		7892 => to_signed(22494, LUT_AMPL_WIDTH),
		7893 => to_signed(22496, LUT_AMPL_WIDTH),
		7894 => to_signed(22498, LUT_AMPL_WIDTH),
		7895 => to_signed(22501, LUT_AMPL_WIDTH),
		7896 => to_signed(22503, LUT_AMPL_WIDTH),
		7897 => to_signed(22505, LUT_AMPL_WIDTH),
		7898 => to_signed(22508, LUT_AMPL_WIDTH),
		7899 => to_signed(22510, LUT_AMPL_WIDTH),
		7900 => to_signed(22512, LUT_AMPL_WIDTH),
		7901 => to_signed(22514, LUT_AMPL_WIDTH),
		7902 => to_signed(22517, LUT_AMPL_WIDTH),
		7903 => to_signed(22519, LUT_AMPL_WIDTH),
		7904 => to_signed(22521, LUT_AMPL_WIDTH),
		7905 => to_signed(22524, LUT_AMPL_WIDTH),
		7906 => to_signed(22526, LUT_AMPL_WIDTH),
		7907 => to_signed(22528, LUT_AMPL_WIDTH),
		7908 => to_signed(22530, LUT_AMPL_WIDTH),
		7909 => to_signed(22533, LUT_AMPL_WIDTH),
		7910 => to_signed(22535, LUT_AMPL_WIDTH),
		7911 => to_signed(22537, LUT_AMPL_WIDTH),
		7912 => to_signed(22540, LUT_AMPL_WIDTH),
		7913 => to_signed(22542, LUT_AMPL_WIDTH),
		7914 => to_signed(22544, LUT_AMPL_WIDTH),
		7915 => to_signed(22546, LUT_AMPL_WIDTH),
		7916 => to_signed(22549, LUT_AMPL_WIDTH),
		7917 => to_signed(22551, LUT_AMPL_WIDTH),
		7918 => to_signed(22553, LUT_AMPL_WIDTH),
		7919 => to_signed(22555, LUT_AMPL_WIDTH),
		7920 => to_signed(22558, LUT_AMPL_WIDTH),
		7921 => to_signed(22560, LUT_AMPL_WIDTH),
		7922 => to_signed(22562, LUT_AMPL_WIDTH),
		7923 => to_signed(22565, LUT_AMPL_WIDTH),
		7924 => to_signed(22567, LUT_AMPL_WIDTH),
		7925 => to_signed(22569, LUT_AMPL_WIDTH),
		7926 => to_signed(22571, LUT_AMPL_WIDTH),
		7927 => to_signed(22574, LUT_AMPL_WIDTH),
		7928 => to_signed(22576, LUT_AMPL_WIDTH),
		7929 => to_signed(22578, LUT_AMPL_WIDTH),
		7930 => to_signed(22581, LUT_AMPL_WIDTH),
		7931 => to_signed(22583, LUT_AMPL_WIDTH),
		7932 => to_signed(22585, LUT_AMPL_WIDTH),
		7933 => to_signed(22587, LUT_AMPL_WIDTH),
		7934 => to_signed(22590, LUT_AMPL_WIDTH),
		7935 => to_signed(22592, LUT_AMPL_WIDTH),
		7936 => to_signed(22594, LUT_AMPL_WIDTH),
		7937 => to_signed(22596, LUT_AMPL_WIDTH),
		7938 => to_signed(22599, LUT_AMPL_WIDTH),
		7939 => to_signed(22601, LUT_AMPL_WIDTH),
		7940 => to_signed(22603, LUT_AMPL_WIDTH),
		7941 => to_signed(22606, LUT_AMPL_WIDTH),
		7942 => to_signed(22608, LUT_AMPL_WIDTH),
		7943 => to_signed(22610, LUT_AMPL_WIDTH),
		7944 => to_signed(22612, LUT_AMPL_WIDTH),
		7945 => to_signed(22615, LUT_AMPL_WIDTH),
		7946 => to_signed(22617, LUT_AMPL_WIDTH),
		7947 => to_signed(22619, LUT_AMPL_WIDTH),
		7948 => to_signed(22621, LUT_AMPL_WIDTH),
		7949 => to_signed(22624, LUT_AMPL_WIDTH),
		7950 => to_signed(22626, LUT_AMPL_WIDTH),
		7951 => to_signed(22628, LUT_AMPL_WIDTH),
		7952 => to_signed(22631, LUT_AMPL_WIDTH),
		7953 => to_signed(22633, LUT_AMPL_WIDTH),
		7954 => to_signed(22635, LUT_AMPL_WIDTH),
		7955 => to_signed(22637, LUT_AMPL_WIDTH),
		7956 => to_signed(22640, LUT_AMPL_WIDTH),
		7957 => to_signed(22642, LUT_AMPL_WIDTH),
		7958 => to_signed(22644, LUT_AMPL_WIDTH),
		7959 => to_signed(22646, LUT_AMPL_WIDTH),
		7960 => to_signed(22649, LUT_AMPL_WIDTH),
		7961 => to_signed(22651, LUT_AMPL_WIDTH),
		7962 => to_signed(22653, LUT_AMPL_WIDTH),
		7963 => to_signed(22656, LUT_AMPL_WIDTH),
		7964 => to_signed(22658, LUT_AMPL_WIDTH),
		7965 => to_signed(22660, LUT_AMPL_WIDTH),
		7966 => to_signed(22662, LUT_AMPL_WIDTH),
		7967 => to_signed(22665, LUT_AMPL_WIDTH),
		7968 => to_signed(22667, LUT_AMPL_WIDTH),
		7969 => to_signed(22669, LUT_AMPL_WIDTH),
		7970 => to_signed(22671, LUT_AMPL_WIDTH),
		7971 => to_signed(22674, LUT_AMPL_WIDTH),
		7972 => to_signed(22676, LUT_AMPL_WIDTH),
		7973 => to_signed(22678, LUT_AMPL_WIDTH),
		7974 => to_signed(22680, LUT_AMPL_WIDTH),
		7975 => to_signed(22683, LUT_AMPL_WIDTH),
		7976 => to_signed(22685, LUT_AMPL_WIDTH),
		7977 => to_signed(22687, LUT_AMPL_WIDTH),
		7978 => to_signed(22690, LUT_AMPL_WIDTH),
		7979 => to_signed(22692, LUT_AMPL_WIDTH),
		7980 => to_signed(22694, LUT_AMPL_WIDTH),
		7981 => to_signed(22696, LUT_AMPL_WIDTH),
		7982 => to_signed(22699, LUT_AMPL_WIDTH),
		7983 => to_signed(22701, LUT_AMPL_WIDTH),
		7984 => to_signed(22703, LUT_AMPL_WIDTH),
		7985 => to_signed(22705, LUT_AMPL_WIDTH),
		7986 => to_signed(22708, LUT_AMPL_WIDTH),
		7987 => to_signed(22710, LUT_AMPL_WIDTH),
		7988 => to_signed(22712, LUT_AMPL_WIDTH),
		7989 => to_signed(22714, LUT_AMPL_WIDTH),
		7990 => to_signed(22717, LUT_AMPL_WIDTH),
		7991 => to_signed(22719, LUT_AMPL_WIDTH),
		7992 => to_signed(22721, LUT_AMPL_WIDTH),
		7993 => to_signed(22724, LUT_AMPL_WIDTH),
		7994 => to_signed(22726, LUT_AMPL_WIDTH),
		7995 => to_signed(22728, LUT_AMPL_WIDTH),
		7996 => to_signed(22730, LUT_AMPL_WIDTH),
		7997 => to_signed(22733, LUT_AMPL_WIDTH),
		7998 => to_signed(22735, LUT_AMPL_WIDTH),
		7999 => to_signed(22737, LUT_AMPL_WIDTH),
		8000 => to_signed(22739, LUT_AMPL_WIDTH),
		8001 => to_signed(22742, LUT_AMPL_WIDTH),
		8002 => to_signed(22744, LUT_AMPL_WIDTH),
		8003 => to_signed(22746, LUT_AMPL_WIDTH),
		8004 => to_signed(22748, LUT_AMPL_WIDTH),
		8005 => to_signed(22751, LUT_AMPL_WIDTH),
		8006 => to_signed(22753, LUT_AMPL_WIDTH),
		8007 => to_signed(22755, LUT_AMPL_WIDTH),
		8008 => to_signed(22757, LUT_AMPL_WIDTH),
		8009 => to_signed(22760, LUT_AMPL_WIDTH),
		8010 => to_signed(22762, LUT_AMPL_WIDTH),
		8011 => to_signed(22764, LUT_AMPL_WIDTH),
		8012 => to_signed(22766, LUT_AMPL_WIDTH),
		8013 => to_signed(22769, LUT_AMPL_WIDTH),
		8014 => to_signed(22771, LUT_AMPL_WIDTH),
		8015 => to_signed(22773, LUT_AMPL_WIDTH),
		8016 => to_signed(22776, LUT_AMPL_WIDTH),
		8017 => to_signed(22778, LUT_AMPL_WIDTH),
		8018 => to_signed(22780, LUT_AMPL_WIDTH),
		8019 => to_signed(22782, LUT_AMPL_WIDTH),
		8020 => to_signed(22785, LUT_AMPL_WIDTH),
		8021 => to_signed(22787, LUT_AMPL_WIDTH),
		8022 => to_signed(22789, LUT_AMPL_WIDTH),
		8023 => to_signed(22791, LUT_AMPL_WIDTH),
		8024 => to_signed(22794, LUT_AMPL_WIDTH),
		8025 => to_signed(22796, LUT_AMPL_WIDTH),
		8026 => to_signed(22798, LUT_AMPL_WIDTH),
		8027 => to_signed(22800, LUT_AMPL_WIDTH),
		8028 => to_signed(22803, LUT_AMPL_WIDTH),
		8029 => to_signed(22805, LUT_AMPL_WIDTH),
		8030 => to_signed(22807, LUT_AMPL_WIDTH),
		8031 => to_signed(22809, LUT_AMPL_WIDTH),
		8032 => to_signed(22812, LUT_AMPL_WIDTH),
		8033 => to_signed(22814, LUT_AMPL_WIDTH),
		8034 => to_signed(22816, LUT_AMPL_WIDTH),
		8035 => to_signed(22818, LUT_AMPL_WIDTH),
		8036 => to_signed(22821, LUT_AMPL_WIDTH),
		8037 => to_signed(22823, LUT_AMPL_WIDTH),
		8038 => to_signed(22825, LUT_AMPL_WIDTH),
		8039 => to_signed(22827, LUT_AMPL_WIDTH),
		8040 => to_signed(22830, LUT_AMPL_WIDTH),
		8041 => to_signed(22832, LUT_AMPL_WIDTH),
		8042 => to_signed(22834, LUT_AMPL_WIDTH),
		8043 => to_signed(22836, LUT_AMPL_WIDTH),
		8044 => to_signed(22839, LUT_AMPL_WIDTH),
		8045 => to_signed(22841, LUT_AMPL_WIDTH),
		8046 => to_signed(22843, LUT_AMPL_WIDTH),
		8047 => to_signed(22845, LUT_AMPL_WIDTH),
		8048 => to_signed(22848, LUT_AMPL_WIDTH),
		8049 => to_signed(22850, LUT_AMPL_WIDTH),
		8050 => to_signed(22852, LUT_AMPL_WIDTH),
		8051 => to_signed(22854, LUT_AMPL_WIDTH),
		8052 => to_signed(22857, LUT_AMPL_WIDTH),
		8053 => to_signed(22859, LUT_AMPL_WIDTH),
		8054 => to_signed(22861, LUT_AMPL_WIDTH),
		8055 => to_signed(22863, LUT_AMPL_WIDTH),
		8056 => to_signed(22866, LUT_AMPL_WIDTH),
		8057 => to_signed(22868, LUT_AMPL_WIDTH),
		8058 => to_signed(22870, LUT_AMPL_WIDTH),
		8059 => to_signed(22872, LUT_AMPL_WIDTH),
		8060 => to_signed(22875, LUT_AMPL_WIDTH),
		8061 => to_signed(22877, LUT_AMPL_WIDTH),
		8062 => to_signed(22879, LUT_AMPL_WIDTH),
		8063 => to_signed(22881, LUT_AMPL_WIDTH),
		8064 => to_signed(22884, LUT_AMPL_WIDTH),
		8065 => to_signed(22886, LUT_AMPL_WIDTH),
		8066 => to_signed(22888, LUT_AMPL_WIDTH),
		8067 => to_signed(22890, LUT_AMPL_WIDTH),
		8068 => to_signed(22893, LUT_AMPL_WIDTH),
		8069 => to_signed(22895, LUT_AMPL_WIDTH),
		8070 => to_signed(22897, LUT_AMPL_WIDTH),
		8071 => to_signed(22899, LUT_AMPL_WIDTH),
		8072 => to_signed(22902, LUT_AMPL_WIDTH),
		8073 => to_signed(22904, LUT_AMPL_WIDTH),
		8074 => to_signed(22906, LUT_AMPL_WIDTH),
		8075 => to_signed(22908, LUT_AMPL_WIDTH),
		8076 => to_signed(22911, LUT_AMPL_WIDTH),
		8077 => to_signed(22913, LUT_AMPL_WIDTH),
		8078 => to_signed(22915, LUT_AMPL_WIDTH),
		8079 => to_signed(22917, LUT_AMPL_WIDTH),
		8080 => to_signed(22920, LUT_AMPL_WIDTH),
		8081 => to_signed(22922, LUT_AMPL_WIDTH),
		8082 => to_signed(22924, LUT_AMPL_WIDTH),
		8083 => to_signed(22926, LUT_AMPL_WIDTH),
		8084 => to_signed(22929, LUT_AMPL_WIDTH),
		8085 => to_signed(22931, LUT_AMPL_WIDTH),
		8086 => to_signed(22933, LUT_AMPL_WIDTH),
		8087 => to_signed(22935, LUT_AMPL_WIDTH),
		8088 => to_signed(22938, LUT_AMPL_WIDTH),
		8089 => to_signed(22940, LUT_AMPL_WIDTH),
		8090 => to_signed(22942, LUT_AMPL_WIDTH),
		8091 => to_signed(22944, LUT_AMPL_WIDTH),
		8092 => to_signed(22947, LUT_AMPL_WIDTH),
		8093 => to_signed(22949, LUT_AMPL_WIDTH),
		8094 => to_signed(22951, LUT_AMPL_WIDTH),
		8095 => to_signed(22953, LUT_AMPL_WIDTH),
		8096 => to_signed(22956, LUT_AMPL_WIDTH),
		8097 => to_signed(22958, LUT_AMPL_WIDTH),
		8098 => to_signed(22960, LUT_AMPL_WIDTH),
		8099 => to_signed(22962, LUT_AMPL_WIDTH),
		8100 => to_signed(22965, LUT_AMPL_WIDTH),
		8101 => to_signed(22967, LUT_AMPL_WIDTH),
		8102 => to_signed(22969, LUT_AMPL_WIDTH),
		8103 => to_signed(22971, LUT_AMPL_WIDTH),
		8104 => to_signed(22973, LUT_AMPL_WIDTH),
		8105 => to_signed(22976, LUT_AMPL_WIDTH),
		8106 => to_signed(22978, LUT_AMPL_WIDTH),
		8107 => to_signed(22980, LUT_AMPL_WIDTH),
		8108 => to_signed(22982, LUT_AMPL_WIDTH),
		8109 => to_signed(22985, LUT_AMPL_WIDTH),
		8110 => to_signed(22987, LUT_AMPL_WIDTH),
		8111 => to_signed(22989, LUT_AMPL_WIDTH),
		8112 => to_signed(22991, LUT_AMPL_WIDTH),
		8113 => to_signed(22994, LUT_AMPL_WIDTH),
		8114 => to_signed(22996, LUT_AMPL_WIDTH),
		8115 => to_signed(22998, LUT_AMPL_WIDTH),
		8116 => to_signed(23000, LUT_AMPL_WIDTH),
		8117 => to_signed(23003, LUT_AMPL_WIDTH),
		8118 => to_signed(23005, LUT_AMPL_WIDTH),
		8119 => to_signed(23007, LUT_AMPL_WIDTH),
		8120 => to_signed(23009, LUT_AMPL_WIDTH),
		8121 => to_signed(23012, LUT_AMPL_WIDTH),
		8122 => to_signed(23014, LUT_AMPL_WIDTH),
		8123 => to_signed(23016, LUT_AMPL_WIDTH),
		8124 => to_signed(23018, LUT_AMPL_WIDTH),
		8125 => to_signed(23020, LUT_AMPL_WIDTH),
		8126 => to_signed(23023, LUT_AMPL_WIDTH),
		8127 => to_signed(23025, LUT_AMPL_WIDTH),
		8128 => to_signed(23027, LUT_AMPL_WIDTH),
		8129 => to_signed(23029, LUT_AMPL_WIDTH),
		8130 => to_signed(23032, LUT_AMPL_WIDTH),
		8131 => to_signed(23034, LUT_AMPL_WIDTH),
		8132 => to_signed(23036, LUT_AMPL_WIDTH),
		8133 => to_signed(23038, LUT_AMPL_WIDTH),
		8134 => to_signed(23041, LUT_AMPL_WIDTH),
		8135 => to_signed(23043, LUT_AMPL_WIDTH),
		8136 => to_signed(23045, LUT_AMPL_WIDTH),
		8137 => to_signed(23047, LUT_AMPL_WIDTH),
		8138 => to_signed(23050, LUT_AMPL_WIDTH),
		8139 => to_signed(23052, LUT_AMPL_WIDTH),
		8140 => to_signed(23054, LUT_AMPL_WIDTH),
		8141 => to_signed(23056, LUT_AMPL_WIDTH),
		8142 => to_signed(23058, LUT_AMPL_WIDTH),
		8143 => to_signed(23061, LUT_AMPL_WIDTH),
		8144 => to_signed(23063, LUT_AMPL_WIDTH),
		8145 => to_signed(23065, LUT_AMPL_WIDTH),
		8146 => to_signed(23067, LUT_AMPL_WIDTH),
		8147 => to_signed(23070, LUT_AMPL_WIDTH),
		8148 => to_signed(23072, LUT_AMPL_WIDTH),
		8149 => to_signed(23074, LUT_AMPL_WIDTH),
		8150 => to_signed(23076, LUT_AMPL_WIDTH),
		8151 => to_signed(23079, LUT_AMPL_WIDTH),
		8152 => to_signed(23081, LUT_AMPL_WIDTH),
		8153 => to_signed(23083, LUT_AMPL_WIDTH),
		8154 => to_signed(23085, LUT_AMPL_WIDTH),
		8155 => to_signed(23087, LUT_AMPL_WIDTH),
		8156 => to_signed(23090, LUT_AMPL_WIDTH),
		8157 => to_signed(23092, LUT_AMPL_WIDTH),
		8158 => to_signed(23094, LUT_AMPL_WIDTH),
		8159 => to_signed(23096, LUT_AMPL_WIDTH),
		8160 => to_signed(23099, LUT_AMPL_WIDTH),
		8161 => to_signed(23101, LUT_AMPL_WIDTH),
		8162 => to_signed(23103, LUT_AMPL_WIDTH),
		8163 => to_signed(23105, LUT_AMPL_WIDTH),
		8164 => to_signed(23107, LUT_AMPL_WIDTH),
		8165 => to_signed(23110, LUT_AMPL_WIDTH),
		8166 => to_signed(23112, LUT_AMPL_WIDTH),
		8167 => to_signed(23114, LUT_AMPL_WIDTH),
		8168 => to_signed(23116, LUT_AMPL_WIDTH),
		8169 => to_signed(23119, LUT_AMPL_WIDTH),
		8170 => to_signed(23121, LUT_AMPL_WIDTH),
		8171 => to_signed(23123, LUT_AMPL_WIDTH),
		8172 => to_signed(23125, LUT_AMPL_WIDTH),
		8173 => to_signed(23128, LUT_AMPL_WIDTH),
		8174 => to_signed(23130, LUT_AMPL_WIDTH),
		8175 => to_signed(23132, LUT_AMPL_WIDTH),
		8176 => to_signed(23134, LUT_AMPL_WIDTH),
		8177 => to_signed(23136, LUT_AMPL_WIDTH),
		8178 => to_signed(23139, LUT_AMPL_WIDTH),
		8179 => to_signed(23141, LUT_AMPL_WIDTH),
		8180 => to_signed(23143, LUT_AMPL_WIDTH),
		8181 => to_signed(23145, LUT_AMPL_WIDTH),
		8182 => to_signed(23148, LUT_AMPL_WIDTH),
		8183 => to_signed(23150, LUT_AMPL_WIDTH),
		8184 => to_signed(23152, LUT_AMPL_WIDTH),
		8185 => to_signed(23154, LUT_AMPL_WIDTH),
		8186 => to_signed(23156, LUT_AMPL_WIDTH),
		8187 => to_signed(23159, LUT_AMPL_WIDTH),
		8188 => to_signed(23161, LUT_AMPL_WIDTH),
		8189 => to_signed(23163, LUT_AMPL_WIDTH),
		8190 => to_signed(23165, LUT_AMPL_WIDTH),
		8191 => to_signed(23168, LUT_AMPL_WIDTH),
		8192 => to_signed(23170, LUT_AMPL_WIDTH),
		8193 => to_signed(23172, LUT_AMPL_WIDTH),
		8194 => to_signed(23174, LUT_AMPL_WIDTH),
		8195 => to_signed(23176, LUT_AMPL_WIDTH),
		8196 => to_signed(23179, LUT_AMPL_WIDTH),
		8197 => to_signed(23181, LUT_AMPL_WIDTH),
		8198 => to_signed(23183, LUT_AMPL_WIDTH),
		8199 => to_signed(23185, LUT_AMPL_WIDTH),
		8200 => to_signed(23188, LUT_AMPL_WIDTH),
		8201 => to_signed(23190, LUT_AMPL_WIDTH),
		8202 => to_signed(23192, LUT_AMPL_WIDTH),
		8203 => to_signed(23194, LUT_AMPL_WIDTH),
		8204 => to_signed(23196, LUT_AMPL_WIDTH),
		8205 => to_signed(23199, LUT_AMPL_WIDTH),
		8206 => to_signed(23201, LUT_AMPL_WIDTH),
		8207 => to_signed(23203, LUT_AMPL_WIDTH),
		8208 => to_signed(23205, LUT_AMPL_WIDTH),
		8209 => to_signed(23208, LUT_AMPL_WIDTH),
		8210 => to_signed(23210, LUT_AMPL_WIDTH),
		8211 => to_signed(23212, LUT_AMPL_WIDTH),
		8212 => to_signed(23214, LUT_AMPL_WIDTH),
		8213 => to_signed(23216, LUT_AMPL_WIDTH),
		8214 => to_signed(23219, LUT_AMPL_WIDTH),
		8215 => to_signed(23221, LUT_AMPL_WIDTH),
		8216 => to_signed(23223, LUT_AMPL_WIDTH),
		8217 => to_signed(23225, LUT_AMPL_WIDTH),
		8218 => to_signed(23227, LUT_AMPL_WIDTH),
		8219 => to_signed(23230, LUT_AMPL_WIDTH),
		8220 => to_signed(23232, LUT_AMPL_WIDTH),
		8221 => to_signed(23234, LUT_AMPL_WIDTH),
		8222 => to_signed(23236, LUT_AMPL_WIDTH),
		8223 => to_signed(23239, LUT_AMPL_WIDTH),
		8224 => to_signed(23241, LUT_AMPL_WIDTH),
		8225 => to_signed(23243, LUT_AMPL_WIDTH),
		8226 => to_signed(23245, LUT_AMPL_WIDTH),
		8227 => to_signed(23247, LUT_AMPL_WIDTH),
		8228 => to_signed(23250, LUT_AMPL_WIDTH),
		8229 => to_signed(23252, LUT_AMPL_WIDTH),
		8230 => to_signed(23254, LUT_AMPL_WIDTH),
		8231 => to_signed(23256, LUT_AMPL_WIDTH),
		8232 => to_signed(23258, LUT_AMPL_WIDTH),
		8233 => to_signed(23261, LUT_AMPL_WIDTH),
		8234 => to_signed(23263, LUT_AMPL_WIDTH),
		8235 => to_signed(23265, LUT_AMPL_WIDTH),
		8236 => to_signed(23267, LUT_AMPL_WIDTH),
		8237 => to_signed(23270, LUT_AMPL_WIDTH),
		8238 => to_signed(23272, LUT_AMPL_WIDTH),
		8239 => to_signed(23274, LUT_AMPL_WIDTH),
		8240 => to_signed(23276, LUT_AMPL_WIDTH),
		8241 => to_signed(23278, LUT_AMPL_WIDTH),
		8242 => to_signed(23281, LUT_AMPL_WIDTH),
		8243 => to_signed(23283, LUT_AMPL_WIDTH),
		8244 => to_signed(23285, LUT_AMPL_WIDTH),
		8245 => to_signed(23287, LUT_AMPL_WIDTH),
		8246 => to_signed(23289, LUT_AMPL_WIDTH),
		8247 => to_signed(23292, LUT_AMPL_WIDTH),
		8248 => to_signed(23294, LUT_AMPL_WIDTH),
		8249 => to_signed(23296, LUT_AMPL_WIDTH),
		8250 => to_signed(23298, LUT_AMPL_WIDTH),
		8251 => to_signed(23300, LUT_AMPL_WIDTH),
		8252 => to_signed(23303, LUT_AMPL_WIDTH),
		8253 => to_signed(23305, LUT_AMPL_WIDTH),
		8254 => to_signed(23307, LUT_AMPL_WIDTH),
		8255 => to_signed(23309, LUT_AMPL_WIDTH),
		8256 => to_signed(23311, LUT_AMPL_WIDTH),
		8257 => to_signed(23314, LUT_AMPL_WIDTH),
		8258 => to_signed(23316, LUT_AMPL_WIDTH),
		8259 => to_signed(23318, LUT_AMPL_WIDTH),
		8260 => to_signed(23320, LUT_AMPL_WIDTH),
		8261 => to_signed(23323, LUT_AMPL_WIDTH),
		8262 => to_signed(23325, LUT_AMPL_WIDTH),
		8263 => to_signed(23327, LUT_AMPL_WIDTH),
		8264 => to_signed(23329, LUT_AMPL_WIDTH),
		8265 => to_signed(23331, LUT_AMPL_WIDTH),
		8266 => to_signed(23334, LUT_AMPL_WIDTH),
		8267 => to_signed(23336, LUT_AMPL_WIDTH),
		8268 => to_signed(23338, LUT_AMPL_WIDTH),
		8269 => to_signed(23340, LUT_AMPL_WIDTH),
		8270 => to_signed(23342, LUT_AMPL_WIDTH),
		8271 => to_signed(23345, LUT_AMPL_WIDTH),
		8272 => to_signed(23347, LUT_AMPL_WIDTH),
		8273 => to_signed(23349, LUT_AMPL_WIDTH),
		8274 => to_signed(23351, LUT_AMPL_WIDTH),
		8275 => to_signed(23353, LUT_AMPL_WIDTH),
		8276 => to_signed(23356, LUT_AMPL_WIDTH),
		8277 => to_signed(23358, LUT_AMPL_WIDTH),
		8278 => to_signed(23360, LUT_AMPL_WIDTH),
		8279 => to_signed(23362, LUT_AMPL_WIDTH),
		8280 => to_signed(23364, LUT_AMPL_WIDTH),
		8281 => to_signed(23367, LUT_AMPL_WIDTH),
		8282 => to_signed(23369, LUT_AMPL_WIDTH),
		8283 => to_signed(23371, LUT_AMPL_WIDTH),
		8284 => to_signed(23373, LUT_AMPL_WIDTH),
		8285 => to_signed(23375, LUT_AMPL_WIDTH),
		8286 => to_signed(23378, LUT_AMPL_WIDTH),
		8287 => to_signed(23380, LUT_AMPL_WIDTH),
		8288 => to_signed(23382, LUT_AMPL_WIDTH),
		8289 => to_signed(23384, LUT_AMPL_WIDTH),
		8290 => to_signed(23386, LUT_AMPL_WIDTH),
		8291 => to_signed(23389, LUT_AMPL_WIDTH),
		8292 => to_signed(23391, LUT_AMPL_WIDTH),
		8293 => to_signed(23393, LUT_AMPL_WIDTH),
		8294 => to_signed(23395, LUT_AMPL_WIDTH),
		8295 => to_signed(23397, LUT_AMPL_WIDTH),
		8296 => to_signed(23400, LUT_AMPL_WIDTH),
		8297 => to_signed(23402, LUT_AMPL_WIDTH),
		8298 => to_signed(23404, LUT_AMPL_WIDTH),
		8299 => to_signed(23406, LUT_AMPL_WIDTH),
		8300 => to_signed(23408, LUT_AMPL_WIDTH),
		8301 => to_signed(23411, LUT_AMPL_WIDTH),
		8302 => to_signed(23413, LUT_AMPL_WIDTH),
		8303 => to_signed(23415, LUT_AMPL_WIDTH),
		8304 => to_signed(23417, LUT_AMPL_WIDTH),
		8305 => to_signed(23419, LUT_AMPL_WIDTH),
		8306 => to_signed(23422, LUT_AMPL_WIDTH),
		8307 => to_signed(23424, LUT_AMPL_WIDTH),
		8308 => to_signed(23426, LUT_AMPL_WIDTH),
		8309 => to_signed(23428, LUT_AMPL_WIDTH),
		8310 => to_signed(23430, LUT_AMPL_WIDTH),
		8311 => to_signed(23433, LUT_AMPL_WIDTH),
		8312 => to_signed(23435, LUT_AMPL_WIDTH),
		8313 => to_signed(23437, LUT_AMPL_WIDTH),
		8314 => to_signed(23439, LUT_AMPL_WIDTH),
		8315 => to_signed(23441, LUT_AMPL_WIDTH),
		8316 => to_signed(23444, LUT_AMPL_WIDTH),
		8317 => to_signed(23446, LUT_AMPL_WIDTH),
		8318 => to_signed(23448, LUT_AMPL_WIDTH),
		8319 => to_signed(23450, LUT_AMPL_WIDTH),
		8320 => to_signed(23452, LUT_AMPL_WIDTH),
		8321 => to_signed(23455, LUT_AMPL_WIDTH),
		8322 => to_signed(23457, LUT_AMPL_WIDTH),
		8323 => to_signed(23459, LUT_AMPL_WIDTH),
		8324 => to_signed(23461, LUT_AMPL_WIDTH),
		8325 => to_signed(23463, LUT_AMPL_WIDTH),
		8326 => to_signed(23466, LUT_AMPL_WIDTH),
		8327 => to_signed(23468, LUT_AMPL_WIDTH),
		8328 => to_signed(23470, LUT_AMPL_WIDTH),
		8329 => to_signed(23472, LUT_AMPL_WIDTH),
		8330 => to_signed(23474, LUT_AMPL_WIDTH),
		8331 => to_signed(23476, LUT_AMPL_WIDTH),
		8332 => to_signed(23479, LUT_AMPL_WIDTH),
		8333 => to_signed(23481, LUT_AMPL_WIDTH),
		8334 => to_signed(23483, LUT_AMPL_WIDTH),
		8335 => to_signed(23485, LUT_AMPL_WIDTH),
		8336 => to_signed(23487, LUT_AMPL_WIDTH),
		8337 => to_signed(23490, LUT_AMPL_WIDTH),
		8338 => to_signed(23492, LUT_AMPL_WIDTH),
		8339 => to_signed(23494, LUT_AMPL_WIDTH),
		8340 => to_signed(23496, LUT_AMPL_WIDTH),
		8341 => to_signed(23498, LUT_AMPL_WIDTH),
		8342 => to_signed(23501, LUT_AMPL_WIDTH),
		8343 => to_signed(23503, LUT_AMPL_WIDTH),
		8344 => to_signed(23505, LUT_AMPL_WIDTH),
		8345 => to_signed(23507, LUT_AMPL_WIDTH),
		8346 => to_signed(23509, LUT_AMPL_WIDTH),
		8347 => to_signed(23512, LUT_AMPL_WIDTH),
		8348 => to_signed(23514, LUT_AMPL_WIDTH),
		8349 => to_signed(23516, LUT_AMPL_WIDTH),
		8350 => to_signed(23518, LUT_AMPL_WIDTH),
		8351 => to_signed(23520, LUT_AMPL_WIDTH),
		8352 => to_signed(23522, LUT_AMPL_WIDTH),
		8353 => to_signed(23525, LUT_AMPL_WIDTH),
		8354 => to_signed(23527, LUT_AMPL_WIDTH),
		8355 => to_signed(23529, LUT_AMPL_WIDTH),
		8356 => to_signed(23531, LUT_AMPL_WIDTH),
		8357 => to_signed(23533, LUT_AMPL_WIDTH),
		8358 => to_signed(23536, LUT_AMPL_WIDTH),
		8359 => to_signed(23538, LUT_AMPL_WIDTH),
		8360 => to_signed(23540, LUT_AMPL_WIDTH),
		8361 => to_signed(23542, LUT_AMPL_WIDTH),
		8362 => to_signed(23544, LUT_AMPL_WIDTH),
		8363 => to_signed(23546, LUT_AMPL_WIDTH),
		8364 => to_signed(23549, LUT_AMPL_WIDTH),
		8365 => to_signed(23551, LUT_AMPL_WIDTH),
		8366 => to_signed(23553, LUT_AMPL_WIDTH),
		8367 => to_signed(23555, LUT_AMPL_WIDTH),
		8368 => to_signed(23557, LUT_AMPL_WIDTH),
		8369 => to_signed(23560, LUT_AMPL_WIDTH),
		8370 => to_signed(23562, LUT_AMPL_WIDTH),
		8371 => to_signed(23564, LUT_AMPL_WIDTH),
		8372 => to_signed(23566, LUT_AMPL_WIDTH),
		8373 => to_signed(23568, LUT_AMPL_WIDTH),
		8374 => to_signed(23571, LUT_AMPL_WIDTH),
		8375 => to_signed(23573, LUT_AMPL_WIDTH),
		8376 => to_signed(23575, LUT_AMPL_WIDTH),
		8377 => to_signed(23577, LUT_AMPL_WIDTH),
		8378 => to_signed(23579, LUT_AMPL_WIDTH),
		8379 => to_signed(23581, LUT_AMPL_WIDTH),
		8380 => to_signed(23584, LUT_AMPL_WIDTH),
		8381 => to_signed(23586, LUT_AMPL_WIDTH),
		8382 => to_signed(23588, LUT_AMPL_WIDTH),
		8383 => to_signed(23590, LUT_AMPL_WIDTH),
		8384 => to_signed(23592, LUT_AMPL_WIDTH),
		8385 => to_signed(23595, LUT_AMPL_WIDTH),
		8386 => to_signed(23597, LUT_AMPL_WIDTH),
		8387 => to_signed(23599, LUT_AMPL_WIDTH),
		8388 => to_signed(23601, LUT_AMPL_WIDTH),
		8389 => to_signed(23603, LUT_AMPL_WIDTH),
		8390 => to_signed(23605, LUT_AMPL_WIDTH),
		8391 => to_signed(23608, LUT_AMPL_WIDTH),
		8392 => to_signed(23610, LUT_AMPL_WIDTH),
		8393 => to_signed(23612, LUT_AMPL_WIDTH),
		8394 => to_signed(23614, LUT_AMPL_WIDTH),
		8395 => to_signed(23616, LUT_AMPL_WIDTH),
		8396 => to_signed(23618, LUT_AMPL_WIDTH),
		8397 => to_signed(23621, LUT_AMPL_WIDTH),
		8398 => to_signed(23623, LUT_AMPL_WIDTH),
		8399 => to_signed(23625, LUT_AMPL_WIDTH),
		8400 => to_signed(23627, LUT_AMPL_WIDTH),
		8401 => to_signed(23629, LUT_AMPL_WIDTH),
		8402 => to_signed(23632, LUT_AMPL_WIDTH),
		8403 => to_signed(23634, LUT_AMPL_WIDTH),
		8404 => to_signed(23636, LUT_AMPL_WIDTH),
		8405 => to_signed(23638, LUT_AMPL_WIDTH),
		8406 => to_signed(23640, LUT_AMPL_WIDTH),
		8407 => to_signed(23642, LUT_AMPL_WIDTH),
		8408 => to_signed(23645, LUT_AMPL_WIDTH),
		8409 => to_signed(23647, LUT_AMPL_WIDTH),
		8410 => to_signed(23649, LUT_AMPL_WIDTH),
		8411 => to_signed(23651, LUT_AMPL_WIDTH),
		8412 => to_signed(23653, LUT_AMPL_WIDTH),
		8413 => to_signed(23655, LUT_AMPL_WIDTH),
		8414 => to_signed(23658, LUT_AMPL_WIDTH),
		8415 => to_signed(23660, LUT_AMPL_WIDTH),
		8416 => to_signed(23662, LUT_AMPL_WIDTH),
		8417 => to_signed(23664, LUT_AMPL_WIDTH),
		8418 => to_signed(23666, LUT_AMPL_WIDTH),
		8419 => to_signed(23668, LUT_AMPL_WIDTH),
		8420 => to_signed(23671, LUT_AMPL_WIDTH),
		8421 => to_signed(23673, LUT_AMPL_WIDTH),
		8422 => to_signed(23675, LUT_AMPL_WIDTH),
		8423 => to_signed(23677, LUT_AMPL_WIDTH),
		8424 => to_signed(23679, LUT_AMPL_WIDTH),
		8425 => to_signed(23682, LUT_AMPL_WIDTH),
		8426 => to_signed(23684, LUT_AMPL_WIDTH),
		8427 => to_signed(23686, LUT_AMPL_WIDTH),
		8428 => to_signed(23688, LUT_AMPL_WIDTH),
		8429 => to_signed(23690, LUT_AMPL_WIDTH),
		8430 => to_signed(23692, LUT_AMPL_WIDTH),
		8431 => to_signed(23695, LUT_AMPL_WIDTH),
		8432 => to_signed(23697, LUT_AMPL_WIDTH),
		8433 => to_signed(23699, LUT_AMPL_WIDTH),
		8434 => to_signed(23701, LUT_AMPL_WIDTH),
		8435 => to_signed(23703, LUT_AMPL_WIDTH),
		8436 => to_signed(23705, LUT_AMPL_WIDTH),
		8437 => to_signed(23708, LUT_AMPL_WIDTH),
		8438 => to_signed(23710, LUT_AMPL_WIDTH),
		8439 => to_signed(23712, LUT_AMPL_WIDTH),
		8440 => to_signed(23714, LUT_AMPL_WIDTH),
		8441 => to_signed(23716, LUT_AMPL_WIDTH),
		8442 => to_signed(23718, LUT_AMPL_WIDTH),
		8443 => to_signed(23721, LUT_AMPL_WIDTH),
		8444 => to_signed(23723, LUT_AMPL_WIDTH),
		8445 => to_signed(23725, LUT_AMPL_WIDTH),
		8446 => to_signed(23727, LUT_AMPL_WIDTH),
		8447 => to_signed(23729, LUT_AMPL_WIDTH),
		8448 => to_signed(23731, LUT_AMPL_WIDTH),
		8449 => to_signed(23734, LUT_AMPL_WIDTH),
		8450 => to_signed(23736, LUT_AMPL_WIDTH),
		8451 => to_signed(23738, LUT_AMPL_WIDTH),
		8452 => to_signed(23740, LUT_AMPL_WIDTH),
		8453 => to_signed(23742, LUT_AMPL_WIDTH),
		8454 => to_signed(23744, LUT_AMPL_WIDTH),
		8455 => to_signed(23747, LUT_AMPL_WIDTH),
		8456 => to_signed(23749, LUT_AMPL_WIDTH),
		8457 => to_signed(23751, LUT_AMPL_WIDTH),
		8458 => to_signed(23753, LUT_AMPL_WIDTH),
		8459 => to_signed(23755, LUT_AMPL_WIDTH),
		8460 => to_signed(23757, LUT_AMPL_WIDTH),
		8461 => to_signed(23760, LUT_AMPL_WIDTH),
		8462 => to_signed(23762, LUT_AMPL_WIDTH),
		8463 => to_signed(23764, LUT_AMPL_WIDTH),
		8464 => to_signed(23766, LUT_AMPL_WIDTH),
		8465 => to_signed(23768, LUT_AMPL_WIDTH),
		8466 => to_signed(23770, LUT_AMPL_WIDTH),
		8467 => to_signed(23773, LUT_AMPL_WIDTH),
		8468 => to_signed(23775, LUT_AMPL_WIDTH),
		8469 => to_signed(23777, LUT_AMPL_WIDTH),
		8470 => to_signed(23779, LUT_AMPL_WIDTH),
		8471 => to_signed(23781, LUT_AMPL_WIDTH),
		8472 => to_signed(23783, LUT_AMPL_WIDTH),
		8473 => to_signed(23785, LUT_AMPL_WIDTH),
		8474 => to_signed(23788, LUT_AMPL_WIDTH),
		8475 => to_signed(23790, LUT_AMPL_WIDTH),
		8476 => to_signed(23792, LUT_AMPL_WIDTH),
		8477 => to_signed(23794, LUT_AMPL_WIDTH),
		8478 => to_signed(23796, LUT_AMPL_WIDTH),
		8479 => to_signed(23798, LUT_AMPL_WIDTH),
		8480 => to_signed(23801, LUT_AMPL_WIDTH),
		8481 => to_signed(23803, LUT_AMPL_WIDTH),
		8482 => to_signed(23805, LUT_AMPL_WIDTH),
		8483 => to_signed(23807, LUT_AMPL_WIDTH),
		8484 => to_signed(23809, LUT_AMPL_WIDTH),
		8485 => to_signed(23811, LUT_AMPL_WIDTH),
		8486 => to_signed(23814, LUT_AMPL_WIDTH),
		8487 => to_signed(23816, LUT_AMPL_WIDTH),
		8488 => to_signed(23818, LUT_AMPL_WIDTH),
		8489 => to_signed(23820, LUT_AMPL_WIDTH),
		8490 => to_signed(23822, LUT_AMPL_WIDTH),
		8491 => to_signed(23824, LUT_AMPL_WIDTH),
		8492 => to_signed(23827, LUT_AMPL_WIDTH),
		8493 => to_signed(23829, LUT_AMPL_WIDTH),
		8494 => to_signed(23831, LUT_AMPL_WIDTH),
		8495 => to_signed(23833, LUT_AMPL_WIDTH),
		8496 => to_signed(23835, LUT_AMPL_WIDTH),
		8497 => to_signed(23837, LUT_AMPL_WIDTH),
		8498 => to_signed(23839, LUT_AMPL_WIDTH),
		8499 => to_signed(23842, LUT_AMPL_WIDTH),
		8500 => to_signed(23844, LUT_AMPL_WIDTH),
		8501 => to_signed(23846, LUT_AMPL_WIDTH),
		8502 => to_signed(23848, LUT_AMPL_WIDTH),
		8503 => to_signed(23850, LUT_AMPL_WIDTH),
		8504 => to_signed(23852, LUT_AMPL_WIDTH),
		8505 => to_signed(23855, LUT_AMPL_WIDTH),
		8506 => to_signed(23857, LUT_AMPL_WIDTH),
		8507 => to_signed(23859, LUT_AMPL_WIDTH),
		8508 => to_signed(23861, LUT_AMPL_WIDTH),
		8509 => to_signed(23863, LUT_AMPL_WIDTH),
		8510 => to_signed(23865, LUT_AMPL_WIDTH),
		8511 => to_signed(23867, LUT_AMPL_WIDTH),
		8512 => to_signed(23870, LUT_AMPL_WIDTH),
		8513 => to_signed(23872, LUT_AMPL_WIDTH),
		8514 => to_signed(23874, LUT_AMPL_WIDTH),
		8515 => to_signed(23876, LUT_AMPL_WIDTH),
		8516 => to_signed(23878, LUT_AMPL_WIDTH),
		8517 => to_signed(23880, LUT_AMPL_WIDTH),
		8518 => to_signed(23883, LUT_AMPL_WIDTH),
		8519 => to_signed(23885, LUT_AMPL_WIDTH),
		8520 => to_signed(23887, LUT_AMPL_WIDTH),
		8521 => to_signed(23889, LUT_AMPL_WIDTH),
		8522 => to_signed(23891, LUT_AMPL_WIDTH),
		8523 => to_signed(23893, LUT_AMPL_WIDTH),
		8524 => to_signed(23895, LUT_AMPL_WIDTH),
		8525 => to_signed(23898, LUT_AMPL_WIDTH),
		8526 => to_signed(23900, LUT_AMPL_WIDTH),
		8527 => to_signed(23902, LUT_AMPL_WIDTH),
		8528 => to_signed(23904, LUT_AMPL_WIDTH),
		8529 => to_signed(23906, LUT_AMPL_WIDTH),
		8530 => to_signed(23908, LUT_AMPL_WIDTH),
		8531 => to_signed(23910, LUT_AMPL_WIDTH),
		8532 => to_signed(23913, LUT_AMPL_WIDTH),
		8533 => to_signed(23915, LUT_AMPL_WIDTH),
		8534 => to_signed(23917, LUT_AMPL_WIDTH),
		8535 => to_signed(23919, LUT_AMPL_WIDTH),
		8536 => to_signed(23921, LUT_AMPL_WIDTH),
		8537 => to_signed(23923, LUT_AMPL_WIDTH),
		8538 => to_signed(23925, LUT_AMPL_WIDTH),
		8539 => to_signed(23928, LUT_AMPL_WIDTH),
		8540 => to_signed(23930, LUT_AMPL_WIDTH),
		8541 => to_signed(23932, LUT_AMPL_WIDTH),
		8542 => to_signed(23934, LUT_AMPL_WIDTH),
		8543 => to_signed(23936, LUT_AMPL_WIDTH),
		8544 => to_signed(23938, LUT_AMPL_WIDTH),
		8545 => to_signed(23940, LUT_AMPL_WIDTH),
		8546 => to_signed(23943, LUT_AMPL_WIDTH),
		8547 => to_signed(23945, LUT_AMPL_WIDTH),
		8548 => to_signed(23947, LUT_AMPL_WIDTH),
		8549 => to_signed(23949, LUT_AMPL_WIDTH),
		8550 => to_signed(23951, LUT_AMPL_WIDTH),
		8551 => to_signed(23953, LUT_AMPL_WIDTH),
		8552 => to_signed(23956, LUT_AMPL_WIDTH),
		8553 => to_signed(23958, LUT_AMPL_WIDTH),
		8554 => to_signed(23960, LUT_AMPL_WIDTH),
		8555 => to_signed(23962, LUT_AMPL_WIDTH),
		8556 => to_signed(23964, LUT_AMPL_WIDTH),
		8557 => to_signed(23966, LUT_AMPL_WIDTH),
		8558 => to_signed(23968, LUT_AMPL_WIDTH),
		8559 => to_signed(23971, LUT_AMPL_WIDTH),
		8560 => to_signed(23973, LUT_AMPL_WIDTH),
		8561 => to_signed(23975, LUT_AMPL_WIDTH),
		8562 => to_signed(23977, LUT_AMPL_WIDTH),
		8563 => to_signed(23979, LUT_AMPL_WIDTH),
		8564 => to_signed(23981, LUT_AMPL_WIDTH),
		8565 => to_signed(23983, LUT_AMPL_WIDTH),
		8566 => to_signed(23985, LUT_AMPL_WIDTH),
		8567 => to_signed(23988, LUT_AMPL_WIDTH),
		8568 => to_signed(23990, LUT_AMPL_WIDTH),
		8569 => to_signed(23992, LUT_AMPL_WIDTH),
		8570 => to_signed(23994, LUT_AMPL_WIDTH),
		8571 => to_signed(23996, LUT_AMPL_WIDTH),
		8572 => to_signed(23998, LUT_AMPL_WIDTH),
		8573 => to_signed(24000, LUT_AMPL_WIDTH),
		8574 => to_signed(24003, LUT_AMPL_WIDTH),
		8575 => to_signed(24005, LUT_AMPL_WIDTH),
		8576 => to_signed(24007, LUT_AMPL_WIDTH),
		8577 => to_signed(24009, LUT_AMPL_WIDTH),
		8578 => to_signed(24011, LUT_AMPL_WIDTH),
		8579 => to_signed(24013, LUT_AMPL_WIDTH),
		8580 => to_signed(24015, LUT_AMPL_WIDTH),
		8581 => to_signed(24018, LUT_AMPL_WIDTH),
		8582 => to_signed(24020, LUT_AMPL_WIDTH),
		8583 => to_signed(24022, LUT_AMPL_WIDTH),
		8584 => to_signed(24024, LUT_AMPL_WIDTH),
		8585 => to_signed(24026, LUT_AMPL_WIDTH),
		8586 => to_signed(24028, LUT_AMPL_WIDTH),
		8587 => to_signed(24030, LUT_AMPL_WIDTH),
		8588 => to_signed(24033, LUT_AMPL_WIDTH),
		8589 => to_signed(24035, LUT_AMPL_WIDTH),
		8590 => to_signed(24037, LUT_AMPL_WIDTH),
		8591 => to_signed(24039, LUT_AMPL_WIDTH),
		8592 => to_signed(24041, LUT_AMPL_WIDTH),
		8593 => to_signed(24043, LUT_AMPL_WIDTH),
		8594 => to_signed(24045, LUT_AMPL_WIDTH),
		8595 => to_signed(24047, LUT_AMPL_WIDTH),
		8596 => to_signed(24050, LUT_AMPL_WIDTH),
		8597 => to_signed(24052, LUT_AMPL_WIDTH),
		8598 => to_signed(24054, LUT_AMPL_WIDTH),
		8599 => to_signed(24056, LUT_AMPL_WIDTH),
		8600 => to_signed(24058, LUT_AMPL_WIDTH),
		8601 => to_signed(24060, LUT_AMPL_WIDTH),
		8602 => to_signed(24062, LUT_AMPL_WIDTH),
		8603 => to_signed(24065, LUT_AMPL_WIDTH),
		8604 => to_signed(24067, LUT_AMPL_WIDTH),
		8605 => to_signed(24069, LUT_AMPL_WIDTH),
		8606 => to_signed(24071, LUT_AMPL_WIDTH),
		8607 => to_signed(24073, LUT_AMPL_WIDTH),
		8608 => to_signed(24075, LUT_AMPL_WIDTH),
		8609 => to_signed(24077, LUT_AMPL_WIDTH),
		8610 => to_signed(24079, LUT_AMPL_WIDTH),
		8611 => to_signed(24082, LUT_AMPL_WIDTH),
		8612 => to_signed(24084, LUT_AMPL_WIDTH),
		8613 => to_signed(24086, LUT_AMPL_WIDTH),
		8614 => to_signed(24088, LUT_AMPL_WIDTH),
		8615 => to_signed(24090, LUT_AMPL_WIDTH),
		8616 => to_signed(24092, LUT_AMPL_WIDTH),
		8617 => to_signed(24094, LUT_AMPL_WIDTH),
		8618 => to_signed(24096, LUT_AMPL_WIDTH),
		8619 => to_signed(24099, LUT_AMPL_WIDTH),
		8620 => to_signed(24101, LUT_AMPL_WIDTH),
		8621 => to_signed(24103, LUT_AMPL_WIDTH),
		8622 => to_signed(24105, LUT_AMPL_WIDTH),
		8623 => to_signed(24107, LUT_AMPL_WIDTH),
		8624 => to_signed(24109, LUT_AMPL_WIDTH),
		8625 => to_signed(24111, LUT_AMPL_WIDTH),
		8626 => to_signed(24114, LUT_AMPL_WIDTH),
		8627 => to_signed(24116, LUT_AMPL_WIDTH),
		8628 => to_signed(24118, LUT_AMPL_WIDTH),
		8629 => to_signed(24120, LUT_AMPL_WIDTH),
		8630 => to_signed(24122, LUT_AMPL_WIDTH),
		8631 => to_signed(24124, LUT_AMPL_WIDTH),
		8632 => to_signed(24126, LUT_AMPL_WIDTH),
		8633 => to_signed(24128, LUT_AMPL_WIDTH),
		8634 => to_signed(24131, LUT_AMPL_WIDTH),
		8635 => to_signed(24133, LUT_AMPL_WIDTH),
		8636 => to_signed(24135, LUT_AMPL_WIDTH),
		8637 => to_signed(24137, LUT_AMPL_WIDTH),
		8638 => to_signed(24139, LUT_AMPL_WIDTH),
		8639 => to_signed(24141, LUT_AMPL_WIDTH),
		8640 => to_signed(24143, LUT_AMPL_WIDTH),
		8641 => to_signed(24145, LUT_AMPL_WIDTH),
		8642 => to_signed(24148, LUT_AMPL_WIDTH),
		8643 => to_signed(24150, LUT_AMPL_WIDTH),
		8644 => to_signed(24152, LUT_AMPL_WIDTH),
		8645 => to_signed(24154, LUT_AMPL_WIDTH),
		8646 => to_signed(24156, LUT_AMPL_WIDTH),
		8647 => to_signed(24158, LUT_AMPL_WIDTH),
		8648 => to_signed(24160, LUT_AMPL_WIDTH),
		8649 => to_signed(24162, LUT_AMPL_WIDTH),
		8650 => to_signed(24164, LUT_AMPL_WIDTH),
		8651 => to_signed(24167, LUT_AMPL_WIDTH),
		8652 => to_signed(24169, LUT_AMPL_WIDTH),
		8653 => to_signed(24171, LUT_AMPL_WIDTH),
		8654 => to_signed(24173, LUT_AMPL_WIDTH),
		8655 => to_signed(24175, LUT_AMPL_WIDTH),
		8656 => to_signed(24177, LUT_AMPL_WIDTH),
		8657 => to_signed(24179, LUT_AMPL_WIDTH),
		8658 => to_signed(24181, LUT_AMPL_WIDTH),
		8659 => to_signed(24184, LUT_AMPL_WIDTH),
		8660 => to_signed(24186, LUT_AMPL_WIDTH),
		8661 => to_signed(24188, LUT_AMPL_WIDTH),
		8662 => to_signed(24190, LUT_AMPL_WIDTH),
		8663 => to_signed(24192, LUT_AMPL_WIDTH),
		8664 => to_signed(24194, LUT_AMPL_WIDTH),
		8665 => to_signed(24196, LUT_AMPL_WIDTH),
		8666 => to_signed(24198, LUT_AMPL_WIDTH),
		8667 => to_signed(24201, LUT_AMPL_WIDTH),
		8668 => to_signed(24203, LUT_AMPL_WIDTH),
		8669 => to_signed(24205, LUT_AMPL_WIDTH),
		8670 => to_signed(24207, LUT_AMPL_WIDTH),
		8671 => to_signed(24209, LUT_AMPL_WIDTH),
		8672 => to_signed(24211, LUT_AMPL_WIDTH),
		8673 => to_signed(24213, LUT_AMPL_WIDTH),
		8674 => to_signed(24215, LUT_AMPL_WIDTH),
		8675 => to_signed(24217, LUT_AMPL_WIDTH),
		8676 => to_signed(24220, LUT_AMPL_WIDTH),
		8677 => to_signed(24222, LUT_AMPL_WIDTH),
		8678 => to_signed(24224, LUT_AMPL_WIDTH),
		8679 => to_signed(24226, LUT_AMPL_WIDTH),
		8680 => to_signed(24228, LUT_AMPL_WIDTH),
		8681 => to_signed(24230, LUT_AMPL_WIDTH),
		8682 => to_signed(24232, LUT_AMPL_WIDTH),
		8683 => to_signed(24234, LUT_AMPL_WIDTH),
		8684 => to_signed(24237, LUT_AMPL_WIDTH),
		8685 => to_signed(24239, LUT_AMPL_WIDTH),
		8686 => to_signed(24241, LUT_AMPL_WIDTH),
		8687 => to_signed(24243, LUT_AMPL_WIDTH),
		8688 => to_signed(24245, LUT_AMPL_WIDTH),
		8689 => to_signed(24247, LUT_AMPL_WIDTH),
		8690 => to_signed(24249, LUT_AMPL_WIDTH),
		8691 => to_signed(24251, LUT_AMPL_WIDTH),
		8692 => to_signed(24253, LUT_AMPL_WIDTH),
		8693 => to_signed(24256, LUT_AMPL_WIDTH),
		8694 => to_signed(24258, LUT_AMPL_WIDTH),
		8695 => to_signed(24260, LUT_AMPL_WIDTH),
		8696 => to_signed(24262, LUT_AMPL_WIDTH),
		8697 => to_signed(24264, LUT_AMPL_WIDTH),
		8698 => to_signed(24266, LUT_AMPL_WIDTH),
		8699 => to_signed(24268, LUT_AMPL_WIDTH),
		8700 => to_signed(24270, LUT_AMPL_WIDTH),
		8701 => to_signed(24272, LUT_AMPL_WIDTH),
		8702 => to_signed(24275, LUT_AMPL_WIDTH),
		8703 => to_signed(24277, LUT_AMPL_WIDTH),
		8704 => to_signed(24279, LUT_AMPL_WIDTH),
		8705 => to_signed(24281, LUT_AMPL_WIDTH),
		8706 => to_signed(24283, LUT_AMPL_WIDTH),
		8707 => to_signed(24285, LUT_AMPL_WIDTH),
		8708 => to_signed(24287, LUT_AMPL_WIDTH),
		8709 => to_signed(24289, LUT_AMPL_WIDTH),
		8710 => to_signed(24291, LUT_AMPL_WIDTH),
		8711 => to_signed(24294, LUT_AMPL_WIDTH),
		8712 => to_signed(24296, LUT_AMPL_WIDTH),
		8713 => to_signed(24298, LUT_AMPL_WIDTH),
		8714 => to_signed(24300, LUT_AMPL_WIDTH),
		8715 => to_signed(24302, LUT_AMPL_WIDTH),
		8716 => to_signed(24304, LUT_AMPL_WIDTH),
		8717 => to_signed(24306, LUT_AMPL_WIDTH),
		8718 => to_signed(24308, LUT_AMPL_WIDTH),
		8719 => to_signed(24310, LUT_AMPL_WIDTH),
		8720 => to_signed(24312, LUT_AMPL_WIDTH),
		8721 => to_signed(24315, LUT_AMPL_WIDTH),
		8722 => to_signed(24317, LUT_AMPL_WIDTH),
		8723 => to_signed(24319, LUT_AMPL_WIDTH),
		8724 => to_signed(24321, LUT_AMPL_WIDTH),
		8725 => to_signed(24323, LUT_AMPL_WIDTH),
		8726 => to_signed(24325, LUT_AMPL_WIDTH),
		8727 => to_signed(24327, LUT_AMPL_WIDTH),
		8728 => to_signed(24329, LUT_AMPL_WIDTH),
		8729 => to_signed(24331, LUT_AMPL_WIDTH),
		8730 => to_signed(24334, LUT_AMPL_WIDTH),
		8731 => to_signed(24336, LUT_AMPL_WIDTH),
		8732 => to_signed(24338, LUT_AMPL_WIDTH),
		8733 => to_signed(24340, LUT_AMPL_WIDTH),
		8734 => to_signed(24342, LUT_AMPL_WIDTH),
		8735 => to_signed(24344, LUT_AMPL_WIDTH),
		8736 => to_signed(24346, LUT_AMPL_WIDTH),
		8737 => to_signed(24348, LUT_AMPL_WIDTH),
		8738 => to_signed(24350, LUT_AMPL_WIDTH),
		8739 => to_signed(24352, LUT_AMPL_WIDTH),
		8740 => to_signed(24355, LUT_AMPL_WIDTH),
		8741 => to_signed(24357, LUT_AMPL_WIDTH),
		8742 => to_signed(24359, LUT_AMPL_WIDTH),
		8743 => to_signed(24361, LUT_AMPL_WIDTH),
		8744 => to_signed(24363, LUT_AMPL_WIDTH),
		8745 => to_signed(24365, LUT_AMPL_WIDTH),
		8746 => to_signed(24367, LUT_AMPL_WIDTH),
		8747 => to_signed(24369, LUT_AMPL_WIDTH),
		8748 => to_signed(24371, LUT_AMPL_WIDTH),
		8749 => to_signed(24373, LUT_AMPL_WIDTH),
		8750 => to_signed(24376, LUT_AMPL_WIDTH),
		8751 => to_signed(24378, LUT_AMPL_WIDTH),
		8752 => to_signed(24380, LUT_AMPL_WIDTH),
		8753 => to_signed(24382, LUT_AMPL_WIDTH),
		8754 => to_signed(24384, LUT_AMPL_WIDTH),
		8755 => to_signed(24386, LUT_AMPL_WIDTH),
		8756 => to_signed(24388, LUT_AMPL_WIDTH),
		8757 => to_signed(24390, LUT_AMPL_WIDTH),
		8758 => to_signed(24392, LUT_AMPL_WIDTH),
		8759 => to_signed(24394, LUT_AMPL_WIDTH),
		8760 => to_signed(24397, LUT_AMPL_WIDTH),
		8761 => to_signed(24399, LUT_AMPL_WIDTH),
		8762 => to_signed(24401, LUT_AMPL_WIDTH),
		8763 => to_signed(24403, LUT_AMPL_WIDTH),
		8764 => to_signed(24405, LUT_AMPL_WIDTH),
		8765 => to_signed(24407, LUT_AMPL_WIDTH),
		8766 => to_signed(24409, LUT_AMPL_WIDTH),
		8767 => to_signed(24411, LUT_AMPL_WIDTH),
		8768 => to_signed(24413, LUT_AMPL_WIDTH),
		8769 => to_signed(24415, LUT_AMPL_WIDTH),
		8770 => to_signed(24417, LUT_AMPL_WIDTH),
		8771 => to_signed(24420, LUT_AMPL_WIDTH),
		8772 => to_signed(24422, LUT_AMPL_WIDTH),
		8773 => to_signed(24424, LUT_AMPL_WIDTH),
		8774 => to_signed(24426, LUT_AMPL_WIDTH),
		8775 => to_signed(24428, LUT_AMPL_WIDTH),
		8776 => to_signed(24430, LUT_AMPL_WIDTH),
		8777 => to_signed(24432, LUT_AMPL_WIDTH),
		8778 => to_signed(24434, LUT_AMPL_WIDTH),
		8779 => to_signed(24436, LUT_AMPL_WIDTH),
		8780 => to_signed(24438, LUT_AMPL_WIDTH),
		8781 => to_signed(24441, LUT_AMPL_WIDTH),
		8782 => to_signed(24443, LUT_AMPL_WIDTH),
		8783 => to_signed(24445, LUT_AMPL_WIDTH),
		8784 => to_signed(24447, LUT_AMPL_WIDTH),
		8785 => to_signed(24449, LUT_AMPL_WIDTH),
		8786 => to_signed(24451, LUT_AMPL_WIDTH),
		8787 => to_signed(24453, LUT_AMPL_WIDTH),
		8788 => to_signed(24455, LUT_AMPL_WIDTH),
		8789 => to_signed(24457, LUT_AMPL_WIDTH),
		8790 => to_signed(24459, LUT_AMPL_WIDTH),
		8791 => to_signed(24461, LUT_AMPL_WIDTH),
		8792 => to_signed(24464, LUT_AMPL_WIDTH),
		8793 => to_signed(24466, LUT_AMPL_WIDTH),
		8794 => to_signed(24468, LUT_AMPL_WIDTH),
		8795 => to_signed(24470, LUT_AMPL_WIDTH),
		8796 => to_signed(24472, LUT_AMPL_WIDTH),
		8797 => to_signed(24474, LUT_AMPL_WIDTH),
		8798 => to_signed(24476, LUT_AMPL_WIDTH),
		8799 => to_signed(24478, LUT_AMPL_WIDTH),
		8800 => to_signed(24480, LUT_AMPL_WIDTH),
		8801 => to_signed(24482, LUT_AMPL_WIDTH),
		8802 => to_signed(24484, LUT_AMPL_WIDTH),
		8803 => to_signed(24487, LUT_AMPL_WIDTH),
		8804 => to_signed(24489, LUT_AMPL_WIDTH),
		8805 => to_signed(24491, LUT_AMPL_WIDTH),
		8806 => to_signed(24493, LUT_AMPL_WIDTH),
		8807 => to_signed(24495, LUT_AMPL_WIDTH),
		8808 => to_signed(24497, LUT_AMPL_WIDTH),
		8809 => to_signed(24499, LUT_AMPL_WIDTH),
		8810 => to_signed(24501, LUT_AMPL_WIDTH),
		8811 => to_signed(24503, LUT_AMPL_WIDTH),
		8812 => to_signed(24505, LUT_AMPL_WIDTH),
		8813 => to_signed(24507, LUT_AMPL_WIDTH),
		8814 => to_signed(24509, LUT_AMPL_WIDTH),
		8815 => to_signed(24512, LUT_AMPL_WIDTH),
		8816 => to_signed(24514, LUT_AMPL_WIDTH),
		8817 => to_signed(24516, LUT_AMPL_WIDTH),
		8818 => to_signed(24518, LUT_AMPL_WIDTH),
		8819 => to_signed(24520, LUT_AMPL_WIDTH),
		8820 => to_signed(24522, LUT_AMPL_WIDTH),
		8821 => to_signed(24524, LUT_AMPL_WIDTH),
		8822 => to_signed(24526, LUT_AMPL_WIDTH),
		8823 => to_signed(24528, LUT_AMPL_WIDTH),
		8824 => to_signed(24530, LUT_AMPL_WIDTH),
		8825 => to_signed(24532, LUT_AMPL_WIDTH),
		8826 => to_signed(24534, LUT_AMPL_WIDTH),
		8827 => to_signed(24537, LUT_AMPL_WIDTH),
		8828 => to_signed(24539, LUT_AMPL_WIDTH),
		8829 => to_signed(24541, LUT_AMPL_WIDTH),
		8830 => to_signed(24543, LUT_AMPL_WIDTH),
		8831 => to_signed(24545, LUT_AMPL_WIDTH),
		8832 => to_signed(24547, LUT_AMPL_WIDTH),
		8833 => to_signed(24549, LUT_AMPL_WIDTH),
		8834 => to_signed(24551, LUT_AMPL_WIDTH),
		8835 => to_signed(24553, LUT_AMPL_WIDTH),
		8836 => to_signed(24555, LUT_AMPL_WIDTH),
		8837 => to_signed(24557, LUT_AMPL_WIDTH),
		8838 => to_signed(24559, LUT_AMPL_WIDTH),
		8839 => to_signed(24562, LUT_AMPL_WIDTH),
		8840 => to_signed(24564, LUT_AMPL_WIDTH),
		8841 => to_signed(24566, LUT_AMPL_WIDTH),
		8842 => to_signed(24568, LUT_AMPL_WIDTH),
		8843 => to_signed(24570, LUT_AMPL_WIDTH),
		8844 => to_signed(24572, LUT_AMPL_WIDTH),
		8845 => to_signed(24574, LUT_AMPL_WIDTH),
		8846 => to_signed(24576, LUT_AMPL_WIDTH),
		8847 => to_signed(24578, LUT_AMPL_WIDTH),
		8848 => to_signed(24580, LUT_AMPL_WIDTH),
		8849 => to_signed(24582, LUT_AMPL_WIDTH),
		8850 => to_signed(24584, LUT_AMPL_WIDTH),
		8851 => to_signed(24586, LUT_AMPL_WIDTH),
		8852 => to_signed(24589, LUT_AMPL_WIDTH),
		8853 => to_signed(24591, LUT_AMPL_WIDTH),
		8854 => to_signed(24593, LUT_AMPL_WIDTH),
		8855 => to_signed(24595, LUT_AMPL_WIDTH),
		8856 => to_signed(24597, LUT_AMPL_WIDTH),
		8857 => to_signed(24599, LUT_AMPL_WIDTH),
		8858 => to_signed(24601, LUT_AMPL_WIDTH),
		8859 => to_signed(24603, LUT_AMPL_WIDTH),
		8860 => to_signed(24605, LUT_AMPL_WIDTH),
		8861 => to_signed(24607, LUT_AMPL_WIDTH),
		8862 => to_signed(24609, LUT_AMPL_WIDTH),
		8863 => to_signed(24611, LUT_AMPL_WIDTH),
		8864 => to_signed(24613, LUT_AMPL_WIDTH),
		8865 => to_signed(24616, LUT_AMPL_WIDTH),
		8866 => to_signed(24618, LUT_AMPL_WIDTH),
		8867 => to_signed(24620, LUT_AMPL_WIDTH),
		8868 => to_signed(24622, LUT_AMPL_WIDTH),
		8869 => to_signed(24624, LUT_AMPL_WIDTH),
		8870 => to_signed(24626, LUT_AMPL_WIDTH),
		8871 => to_signed(24628, LUT_AMPL_WIDTH),
		8872 => to_signed(24630, LUT_AMPL_WIDTH),
		8873 => to_signed(24632, LUT_AMPL_WIDTH),
		8874 => to_signed(24634, LUT_AMPL_WIDTH),
		8875 => to_signed(24636, LUT_AMPL_WIDTH),
		8876 => to_signed(24638, LUT_AMPL_WIDTH),
		8877 => to_signed(24640, LUT_AMPL_WIDTH),
		8878 => to_signed(24642, LUT_AMPL_WIDTH),
		8879 => to_signed(24645, LUT_AMPL_WIDTH),
		8880 => to_signed(24647, LUT_AMPL_WIDTH),
		8881 => to_signed(24649, LUT_AMPL_WIDTH),
		8882 => to_signed(24651, LUT_AMPL_WIDTH),
		8883 => to_signed(24653, LUT_AMPL_WIDTH),
		8884 => to_signed(24655, LUT_AMPL_WIDTH),
		8885 => to_signed(24657, LUT_AMPL_WIDTH),
		8886 => to_signed(24659, LUT_AMPL_WIDTH),
		8887 => to_signed(24661, LUT_AMPL_WIDTH),
		8888 => to_signed(24663, LUT_AMPL_WIDTH),
		8889 => to_signed(24665, LUT_AMPL_WIDTH),
		8890 => to_signed(24667, LUT_AMPL_WIDTH),
		8891 => to_signed(24669, LUT_AMPL_WIDTH),
		8892 => to_signed(24671, LUT_AMPL_WIDTH),
		8893 => to_signed(24673, LUT_AMPL_WIDTH),
		8894 => to_signed(24676, LUT_AMPL_WIDTH),
		8895 => to_signed(24678, LUT_AMPL_WIDTH),
		8896 => to_signed(24680, LUT_AMPL_WIDTH),
		8897 => to_signed(24682, LUT_AMPL_WIDTH),
		8898 => to_signed(24684, LUT_AMPL_WIDTH),
		8899 => to_signed(24686, LUT_AMPL_WIDTH),
		8900 => to_signed(24688, LUT_AMPL_WIDTH),
		8901 => to_signed(24690, LUT_AMPL_WIDTH),
		8902 => to_signed(24692, LUT_AMPL_WIDTH),
		8903 => to_signed(24694, LUT_AMPL_WIDTH),
		8904 => to_signed(24696, LUT_AMPL_WIDTH),
		8905 => to_signed(24698, LUT_AMPL_WIDTH),
		8906 => to_signed(24700, LUT_AMPL_WIDTH),
		8907 => to_signed(24702, LUT_AMPL_WIDTH),
		8908 => to_signed(24704, LUT_AMPL_WIDTH),
		8909 => to_signed(24707, LUT_AMPL_WIDTH),
		8910 => to_signed(24709, LUT_AMPL_WIDTH),
		8911 => to_signed(24711, LUT_AMPL_WIDTH),
		8912 => to_signed(24713, LUT_AMPL_WIDTH),
		8913 => to_signed(24715, LUT_AMPL_WIDTH),
		8914 => to_signed(24717, LUT_AMPL_WIDTH),
		8915 => to_signed(24719, LUT_AMPL_WIDTH),
		8916 => to_signed(24721, LUT_AMPL_WIDTH),
		8917 => to_signed(24723, LUT_AMPL_WIDTH),
		8918 => to_signed(24725, LUT_AMPL_WIDTH),
		8919 => to_signed(24727, LUT_AMPL_WIDTH),
		8920 => to_signed(24729, LUT_AMPL_WIDTH),
		8921 => to_signed(24731, LUT_AMPL_WIDTH),
		8922 => to_signed(24733, LUT_AMPL_WIDTH),
		8923 => to_signed(24735, LUT_AMPL_WIDTH),
		8924 => to_signed(24737, LUT_AMPL_WIDTH),
		8925 => to_signed(24740, LUT_AMPL_WIDTH),
		8926 => to_signed(24742, LUT_AMPL_WIDTH),
		8927 => to_signed(24744, LUT_AMPL_WIDTH),
		8928 => to_signed(24746, LUT_AMPL_WIDTH),
		8929 => to_signed(24748, LUT_AMPL_WIDTH),
		8930 => to_signed(24750, LUT_AMPL_WIDTH),
		8931 => to_signed(24752, LUT_AMPL_WIDTH),
		8932 => to_signed(24754, LUT_AMPL_WIDTH),
		8933 => to_signed(24756, LUT_AMPL_WIDTH),
		8934 => to_signed(24758, LUT_AMPL_WIDTH),
		8935 => to_signed(24760, LUT_AMPL_WIDTH),
		8936 => to_signed(24762, LUT_AMPL_WIDTH),
		8937 => to_signed(24764, LUT_AMPL_WIDTH),
		8938 => to_signed(24766, LUT_AMPL_WIDTH),
		8939 => to_signed(24768, LUT_AMPL_WIDTH),
		8940 => to_signed(24770, LUT_AMPL_WIDTH),
		8941 => to_signed(24772, LUT_AMPL_WIDTH),
		8942 => to_signed(24774, LUT_AMPL_WIDTH),
		8943 => to_signed(24777, LUT_AMPL_WIDTH),
		8944 => to_signed(24779, LUT_AMPL_WIDTH),
		8945 => to_signed(24781, LUT_AMPL_WIDTH),
		8946 => to_signed(24783, LUT_AMPL_WIDTH),
		8947 => to_signed(24785, LUT_AMPL_WIDTH),
		8948 => to_signed(24787, LUT_AMPL_WIDTH),
		8949 => to_signed(24789, LUT_AMPL_WIDTH),
		8950 => to_signed(24791, LUT_AMPL_WIDTH),
		8951 => to_signed(24793, LUT_AMPL_WIDTH),
		8952 => to_signed(24795, LUT_AMPL_WIDTH),
		8953 => to_signed(24797, LUT_AMPL_WIDTH),
		8954 => to_signed(24799, LUT_AMPL_WIDTH),
		8955 => to_signed(24801, LUT_AMPL_WIDTH),
		8956 => to_signed(24803, LUT_AMPL_WIDTH),
		8957 => to_signed(24805, LUT_AMPL_WIDTH),
		8958 => to_signed(24807, LUT_AMPL_WIDTH),
		8959 => to_signed(24809, LUT_AMPL_WIDTH),
		8960 => to_signed(24811, LUT_AMPL_WIDTH),
		8961 => to_signed(24814, LUT_AMPL_WIDTH),
		8962 => to_signed(24816, LUT_AMPL_WIDTH),
		8963 => to_signed(24818, LUT_AMPL_WIDTH),
		8964 => to_signed(24820, LUT_AMPL_WIDTH),
		8965 => to_signed(24822, LUT_AMPL_WIDTH),
		8966 => to_signed(24824, LUT_AMPL_WIDTH),
		8967 => to_signed(24826, LUT_AMPL_WIDTH),
		8968 => to_signed(24828, LUT_AMPL_WIDTH),
		8969 => to_signed(24830, LUT_AMPL_WIDTH),
		8970 => to_signed(24832, LUT_AMPL_WIDTH),
		8971 => to_signed(24834, LUT_AMPL_WIDTH),
		8972 => to_signed(24836, LUT_AMPL_WIDTH),
		8973 => to_signed(24838, LUT_AMPL_WIDTH),
		8974 => to_signed(24840, LUT_AMPL_WIDTH),
		8975 => to_signed(24842, LUT_AMPL_WIDTH),
		8976 => to_signed(24844, LUT_AMPL_WIDTH),
		8977 => to_signed(24846, LUT_AMPL_WIDTH),
		8978 => to_signed(24848, LUT_AMPL_WIDTH),
		8979 => to_signed(24850, LUT_AMPL_WIDTH),
		8980 => to_signed(24852, LUT_AMPL_WIDTH),
		8981 => to_signed(24855, LUT_AMPL_WIDTH),
		8982 => to_signed(24857, LUT_AMPL_WIDTH),
		8983 => to_signed(24859, LUT_AMPL_WIDTH),
		8984 => to_signed(24861, LUT_AMPL_WIDTH),
		8985 => to_signed(24863, LUT_AMPL_WIDTH),
		8986 => to_signed(24865, LUT_AMPL_WIDTH),
		8987 => to_signed(24867, LUT_AMPL_WIDTH),
		8988 => to_signed(24869, LUT_AMPL_WIDTH),
		8989 => to_signed(24871, LUT_AMPL_WIDTH),
		8990 => to_signed(24873, LUT_AMPL_WIDTH),
		8991 => to_signed(24875, LUT_AMPL_WIDTH),
		8992 => to_signed(24877, LUT_AMPL_WIDTH),
		8993 => to_signed(24879, LUT_AMPL_WIDTH),
		8994 => to_signed(24881, LUT_AMPL_WIDTH),
		8995 => to_signed(24883, LUT_AMPL_WIDTH),
		8996 => to_signed(24885, LUT_AMPL_WIDTH),
		8997 => to_signed(24887, LUT_AMPL_WIDTH),
		8998 => to_signed(24889, LUT_AMPL_WIDTH),
		8999 => to_signed(24891, LUT_AMPL_WIDTH),
		9000 => to_signed(24893, LUT_AMPL_WIDTH),
		9001 => to_signed(24895, LUT_AMPL_WIDTH),
		9002 => to_signed(24897, LUT_AMPL_WIDTH),
		9003 => to_signed(24899, LUT_AMPL_WIDTH),
		9004 => to_signed(24902, LUT_AMPL_WIDTH),
		9005 => to_signed(24904, LUT_AMPL_WIDTH),
		9006 => to_signed(24906, LUT_AMPL_WIDTH),
		9007 => to_signed(24908, LUT_AMPL_WIDTH),
		9008 => to_signed(24910, LUT_AMPL_WIDTH),
		9009 => to_signed(24912, LUT_AMPL_WIDTH),
		9010 => to_signed(24914, LUT_AMPL_WIDTH),
		9011 => to_signed(24916, LUT_AMPL_WIDTH),
		9012 => to_signed(24918, LUT_AMPL_WIDTH),
		9013 => to_signed(24920, LUT_AMPL_WIDTH),
		9014 => to_signed(24922, LUT_AMPL_WIDTH),
		9015 => to_signed(24924, LUT_AMPL_WIDTH),
		9016 => to_signed(24926, LUT_AMPL_WIDTH),
		9017 => to_signed(24928, LUT_AMPL_WIDTH),
		9018 => to_signed(24930, LUT_AMPL_WIDTH),
		9019 => to_signed(24932, LUT_AMPL_WIDTH),
		9020 => to_signed(24934, LUT_AMPL_WIDTH),
		9021 => to_signed(24936, LUT_AMPL_WIDTH),
		9022 => to_signed(24938, LUT_AMPL_WIDTH),
		9023 => to_signed(24940, LUT_AMPL_WIDTH),
		9024 => to_signed(24942, LUT_AMPL_WIDTH),
		9025 => to_signed(24944, LUT_AMPL_WIDTH),
		9026 => to_signed(24946, LUT_AMPL_WIDTH),
		9027 => to_signed(24948, LUT_AMPL_WIDTH),
		9028 => to_signed(24950, LUT_AMPL_WIDTH),
		9029 => to_signed(24953, LUT_AMPL_WIDTH),
		9030 => to_signed(24955, LUT_AMPL_WIDTH),
		9031 => to_signed(24957, LUT_AMPL_WIDTH),
		9032 => to_signed(24959, LUT_AMPL_WIDTH),
		9033 => to_signed(24961, LUT_AMPL_WIDTH),
		9034 => to_signed(24963, LUT_AMPL_WIDTH),
		9035 => to_signed(24965, LUT_AMPL_WIDTH),
		9036 => to_signed(24967, LUT_AMPL_WIDTH),
		9037 => to_signed(24969, LUT_AMPL_WIDTH),
		9038 => to_signed(24971, LUT_AMPL_WIDTH),
		9039 => to_signed(24973, LUT_AMPL_WIDTH),
		9040 => to_signed(24975, LUT_AMPL_WIDTH),
		9041 => to_signed(24977, LUT_AMPL_WIDTH),
		9042 => to_signed(24979, LUT_AMPL_WIDTH),
		9043 => to_signed(24981, LUT_AMPL_WIDTH),
		9044 => to_signed(24983, LUT_AMPL_WIDTH),
		9045 => to_signed(24985, LUT_AMPL_WIDTH),
		9046 => to_signed(24987, LUT_AMPL_WIDTH),
		9047 => to_signed(24989, LUT_AMPL_WIDTH),
		9048 => to_signed(24991, LUT_AMPL_WIDTH),
		9049 => to_signed(24993, LUT_AMPL_WIDTH),
		9050 => to_signed(24995, LUT_AMPL_WIDTH),
		9051 => to_signed(24997, LUT_AMPL_WIDTH),
		9052 => to_signed(24999, LUT_AMPL_WIDTH),
		9053 => to_signed(25001, LUT_AMPL_WIDTH),
		9054 => to_signed(25003, LUT_AMPL_WIDTH),
		9055 => to_signed(25005, LUT_AMPL_WIDTH),
		9056 => to_signed(25007, LUT_AMPL_WIDTH),
		9057 => to_signed(25009, LUT_AMPL_WIDTH),
		9058 => to_signed(25011, LUT_AMPL_WIDTH),
		9059 => to_signed(25013, LUT_AMPL_WIDTH),
		9060 => to_signed(25016, LUT_AMPL_WIDTH),
		9061 => to_signed(25018, LUT_AMPL_WIDTH),
		9062 => to_signed(25020, LUT_AMPL_WIDTH),
		9063 => to_signed(25022, LUT_AMPL_WIDTH),
		9064 => to_signed(25024, LUT_AMPL_WIDTH),
		9065 => to_signed(25026, LUT_AMPL_WIDTH),
		9066 => to_signed(25028, LUT_AMPL_WIDTH),
		9067 => to_signed(25030, LUT_AMPL_WIDTH),
		9068 => to_signed(25032, LUT_AMPL_WIDTH),
		9069 => to_signed(25034, LUT_AMPL_WIDTH),
		9070 => to_signed(25036, LUT_AMPL_WIDTH),
		9071 => to_signed(25038, LUT_AMPL_WIDTH),
		9072 => to_signed(25040, LUT_AMPL_WIDTH),
		9073 => to_signed(25042, LUT_AMPL_WIDTH),
		9074 => to_signed(25044, LUT_AMPL_WIDTH),
		9075 => to_signed(25046, LUT_AMPL_WIDTH),
		9076 => to_signed(25048, LUT_AMPL_WIDTH),
		9077 => to_signed(25050, LUT_AMPL_WIDTH),
		9078 => to_signed(25052, LUT_AMPL_WIDTH),
		9079 => to_signed(25054, LUT_AMPL_WIDTH),
		9080 => to_signed(25056, LUT_AMPL_WIDTH),
		9081 => to_signed(25058, LUT_AMPL_WIDTH),
		9082 => to_signed(25060, LUT_AMPL_WIDTH),
		9083 => to_signed(25062, LUT_AMPL_WIDTH),
		9084 => to_signed(25064, LUT_AMPL_WIDTH),
		9085 => to_signed(25066, LUT_AMPL_WIDTH),
		9086 => to_signed(25068, LUT_AMPL_WIDTH),
		9087 => to_signed(25070, LUT_AMPL_WIDTH),
		9088 => to_signed(25072, LUT_AMPL_WIDTH),
		9089 => to_signed(25074, LUT_AMPL_WIDTH),
		9090 => to_signed(25076, LUT_AMPL_WIDTH),
		9091 => to_signed(25078, LUT_AMPL_WIDTH),
		9092 => to_signed(25080, LUT_AMPL_WIDTH),
		9093 => to_signed(25082, LUT_AMPL_WIDTH),
		9094 => to_signed(25084, LUT_AMPL_WIDTH),
		9095 => to_signed(25086, LUT_AMPL_WIDTH),
		9096 => to_signed(25088, LUT_AMPL_WIDTH),
		9097 => to_signed(25090, LUT_AMPL_WIDTH),
		9098 => to_signed(25092, LUT_AMPL_WIDTH),
		9099 => to_signed(25094, LUT_AMPL_WIDTH),
		9100 => to_signed(25096, LUT_AMPL_WIDTH),
		9101 => to_signed(25099, LUT_AMPL_WIDTH),
		9102 => to_signed(25101, LUT_AMPL_WIDTH),
		9103 => to_signed(25103, LUT_AMPL_WIDTH),
		9104 => to_signed(25105, LUT_AMPL_WIDTH),
		9105 => to_signed(25107, LUT_AMPL_WIDTH),
		9106 => to_signed(25109, LUT_AMPL_WIDTH),
		9107 => to_signed(25111, LUT_AMPL_WIDTH),
		9108 => to_signed(25113, LUT_AMPL_WIDTH),
		9109 => to_signed(25115, LUT_AMPL_WIDTH),
		9110 => to_signed(25117, LUT_AMPL_WIDTH),
		9111 => to_signed(25119, LUT_AMPL_WIDTH),
		9112 => to_signed(25121, LUT_AMPL_WIDTH),
		9113 => to_signed(25123, LUT_AMPL_WIDTH),
		9114 => to_signed(25125, LUT_AMPL_WIDTH),
		9115 => to_signed(25127, LUT_AMPL_WIDTH),
		9116 => to_signed(25129, LUT_AMPL_WIDTH),
		9117 => to_signed(25131, LUT_AMPL_WIDTH),
		9118 => to_signed(25133, LUT_AMPL_WIDTH),
		9119 => to_signed(25135, LUT_AMPL_WIDTH),
		9120 => to_signed(25137, LUT_AMPL_WIDTH),
		9121 => to_signed(25139, LUT_AMPL_WIDTH),
		9122 => to_signed(25141, LUT_AMPL_WIDTH),
		9123 => to_signed(25143, LUT_AMPL_WIDTH),
		9124 => to_signed(25145, LUT_AMPL_WIDTH),
		9125 => to_signed(25147, LUT_AMPL_WIDTH),
		9126 => to_signed(25149, LUT_AMPL_WIDTH),
		9127 => to_signed(25151, LUT_AMPL_WIDTH),
		9128 => to_signed(25153, LUT_AMPL_WIDTH),
		9129 => to_signed(25155, LUT_AMPL_WIDTH),
		9130 => to_signed(25157, LUT_AMPL_WIDTH),
		9131 => to_signed(25159, LUT_AMPL_WIDTH),
		9132 => to_signed(25161, LUT_AMPL_WIDTH),
		9133 => to_signed(25163, LUT_AMPL_WIDTH),
		9134 => to_signed(25165, LUT_AMPL_WIDTH),
		9135 => to_signed(25167, LUT_AMPL_WIDTH),
		9136 => to_signed(25169, LUT_AMPL_WIDTH),
		9137 => to_signed(25171, LUT_AMPL_WIDTH),
		9138 => to_signed(25173, LUT_AMPL_WIDTH),
		9139 => to_signed(25175, LUT_AMPL_WIDTH),
		9140 => to_signed(25177, LUT_AMPL_WIDTH),
		9141 => to_signed(25179, LUT_AMPL_WIDTH),
		9142 => to_signed(25181, LUT_AMPL_WIDTH),
		9143 => to_signed(25183, LUT_AMPL_WIDTH),
		9144 => to_signed(25185, LUT_AMPL_WIDTH),
		9145 => to_signed(25187, LUT_AMPL_WIDTH),
		9146 => to_signed(25189, LUT_AMPL_WIDTH),
		9147 => to_signed(25191, LUT_AMPL_WIDTH),
		9148 => to_signed(25193, LUT_AMPL_WIDTH),
		9149 => to_signed(25195, LUT_AMPL_WIDTH),
		9150 => to_signed(25197, LUT_AMPL_WIDTH),
		9151 => to_signed(25199, LUT_AMPL_WIDTH),
		9152 => to_signed(25201, LUT_AMPL_WIDTH),
		9153 => to_signed(25203, LUT_AMPL_WIDTH),
		9154 => to_signed(25205, LUT_AMPL_WIDTH),
		9155 => to_signed(25207, LUT_AMPL_WIDTH),
		9156 => to_signed(25209, LUT_AMPL_WIDTH),
		9157 => to_signed(25211, LUT_AMPL_WIDTH),
		9158 => to_signed(25213, LUT_AMPL_WIDTH),
		9159 => to_signed(25215, LUT_AMPL_WIDTH),
		9160 => to_signed(25217, LUT_AMPL_WIDTH),
		9161 => to_signed(25219, LUT_AMPL_WIDTH),
		9162 => to_signed(25221, LUT_AMPL_WIDTH),
		9163 => to_signed(25223, LUT_AMPL_WIDTH),
		9164 => to_signed(25225, LUT_AMPL_WIDTH),
		9165 => to_signed(25227, LUT_AMPL_WIDTH),
		9166 => to_signed(25229, LUT_AMPL_WIDTH),
		9167 => to_signed(25231, LUT_AMPL_WIDTH),
		9168 => to_signed(25233, LUT_AMPL_WIDTH),
		9169 => to_signed(25235, LUT_AMPL_WIDTH),
		9170 => to_signed(25237, LUT_AMPL_WIDTH),
		9171 => to_signed(25239, LUT_AMPL_WIDTH),
		9172 => to_signed(25241, LUT_AMPL_WIDTH),
		9173 => to_signed(25243, LUT_AMPL_WIDTH),
		9174 => to_signed(25245, LUT_AMPL_WIDTH),
		9175 => to_signed(25247, LUT_AMPL_WIDTH),
		9176 => to_signed(25249, LUT_AMPL_WIDTH),
		9177 => to_signed(25251, LUT_AMPL_WIDTH),
		9178 => to_signed(25253, LUT_AMPL_WIDTH),
		9179 => to_signed(25255, LUT_AMPL_WIDTH),
		9180 => to_signed(25257, LUT_AMPL_WIDTH),
		9181 => to_signed(25259, LUT_AMPL_WIDTH),
		9182 => to_signed(25261, LUT_AMPL_WIDTH),
		9183 => to_signed(25263, LUT_AMPL_WIDTH),
		9184 => to_signed(25265, LUT_AMPL_WIDTH),
		9185 => to_signed(25267, LUT_AMPL_WIDTH),
		9186 => to_signed(25269, LUT_AMPL_WIDTH),
		9187 => to_signed(25271, LUT_AMPL_WIDTH),
		9188 => to_signed(25273, LUT_AMPL_WIDTH),
		9189 => to_signed(25275, LUT_AMPL_WIDTH),
		9190 => to_signed(25277, LUT_AMPL_WIDTH),
		9191 => to_signed(25279, LUT_AMPL_WIDTH),
		9192 => to_signed(25281, LUT_AMPL_WIDTH),
		9193 => to_signed(25283, LUT_AMPL_WIDTH),
		9194 => to_signed(25285, LUT_AMPL_WIDTH),
		9195 => to_signed(25287, LUT_AMPL_WIDTH),
		9196 => to_signed(25289, LUT_AMPL_WIDTH),
		9197 => to_signed(25291, LUT_AMPL_WIDTH),
		9198 => to_signed(25293, LUT_AMPL_WIDTH),
		9199 => to_signed(25295, LUT_AMPL_WIDTH),
		9200 => to_signed(25297, LUT_AMPL_WIDTH),
		9201 => to_signed(25299, LUT_AMPL_WIDTH),
		9202 => to_signed(25301, LUT_AMPL_WIDTH),
		9203 => to_signed(25303, LUT_AMPL_WIDTH),
		9204 => to_signed(25305, LUT_AMPL_WIDTH),
		9205 => to_signed(25307, LUT_AMPL_WIDTH),
		9206 => to_signed(25309, LUT_AMPL_WIDTH),
		9207 => to_signed(25311, LUT_AMPL_WIDTH),
		9208 => to_signed(25313, LUT_AMPL_WIDTH),
		9209 => to_signed(25315, LUT_AMPL_WIDTH),
		9210 => to_signed(25317, LUT_AMPL_WIDTH),
		9211 => to_signed(25319, LUT_AMPL_WIDTH),
		9212 => to_signed(25321, LUT_AMPL_WIDTH),
		9213 => to_signed(25323, LUT_AMPL_WIDTH),
		9214 => to_signed(25325, LUT_AMPL_WIDTH),
		9215 => to_signed(25327, LUT_AMPL_WIDTH),
		9216 => to_signed(25329, LUT_AMPL_WIDTH),
		9217 => to_signed(25331, LUT_AMPL_WIDTH),
		9218 => to_signed(25333, LUT_AMPL_WIDTH),
		9219 => to_signed(25335, LUT_AMPL_WIDTH),
		9220 => to_signed(25337, LUT_AMPL_WIDTH),
		9221 => to_signed(25339, LUT_AMPL_WIDTH),
		9222 => to_signed(25341, LUT_AMPL_WIDTH),
		9223 => to_signed(25343, LUT_AMPL_WIDTH),
		9224 => to_signed(25345, LUT_AMPL_WIDTH),
		9225 => to_signed(25347, LUT_AMPL_WIDTH),
		9226 => to_signed(25349, LUT_AMPL_WIDTH),
		9227 => to_signed(25351, LUT_AMPL_WIDTH),
		9228 => to_signed(25353, LUT_AMPL_WIDTH),
		9229 => to_signed(25355, LUT_AMPL_WIDTH),
		9230 => to_signed(25357, LUT_AMPL_WIDTH),
		9231 => to_signed(25359, LUT_AMPL_WIDTH),
		9232 => to_signed(25361, LUT_AMPL_WIDTH),
		9233 => to_signed(25363, LUT_AMPL_WIDTH),
		9234 => to_signed(25365, LUT_AMPL_WIDTH),
		9235 => to_signed(25367, LUT_AMPL_WIDTH),
		9236 => to_signed(25369, LUT_AMPL_WIDTH),
		9237 => to_signed(25371, LUT_AMPL_WIDTH),
		9238 => to_signed(25373, LUT_AMPL_WIDTH),
		9239 => to_signed(25375, LUT_AMPL_WIDTH),
		9240 => to_signed(25377, LUT_AMPL_WIDTH),
		9241 => to_signed(25379, LUT_AMPL_WIDTH),
		9242 => to_signed(25381, LUT_AMPL_WIDTH),
		9243 => to_signed(25383, LUT_AMPL_WIDTH),
		9244 => to_signed(25385, LUT_AMPL_WIDTH),
		9245 => to_signed(25387, LUT_AMPL_WIDTH),
		9246 => to_signed(25389, LUT_AMPL_WIDTH),
		9247 => to_signed(25391, LUT_AMPL_WIDTH),
		9248 => to_signed(25393, LUT_AMPL_WIDTH),
		9249 => to_signed(25395, LUT_AMPL_WIDTH),
		9250 => to_signed(25397, LUT_AMPL_WIDTH),
		9251 => to_signed(25399, LUT_AMPL_WIDTH),
		9252 => to_signed(25401, LUT_AMPL_WIDTH),
		9253 => to_signed(25403, LUT_AMPL_WIDTH),
		9254 => to_signed(25405, LUT_AMPL_WIDTH),
		9255 => to_signed(25407, LUT_AMPL_WIDTH),
		9256 => to_signed(25409, LUT_AMPL_WIDTH),
		9257 => to_signed(25411, LUT_AMPL_WIDTH),
		9258 => to_signed(25413, LUT_AMPL_WIDTH),
		9259 => to_signed(25415, LUT_AMPL_WIDTH),
		9260 => to_signed(25417, LUT_AMPL_WIDTH),
		9261 => to_signed(25419, LUT_AMPL_WIDTH),
		9262 => to_signed(25421, LUT_AMPL_WIDTH),
		9263 => to_signed(25423, LUT_AMPL_WIDTH),
		9264 => to_signed(25425, LUT_AMPL_WIDTH),
		9265 => to_signed(25427, LUT_AMPL_WIDTH),
		9266 => to_signed(25429, LUT_AMPL_WIDTH),
		9267 => to_signed(25431, LUT_AMPL_WIDTH),
		9268 => to_signed(25433, LUT_AMPL_WIDTH),
		9269 => to_signed(25435, LUT_AMPL_WIDTH),
		9270 => to_signed(25437, LUT_AMPL_WIDTH),
		9271 => to_signed(25438, LUT_AMPL_WIDTH),
		9272 => to_signed(25440, LUT_AMPL_WIDTH),
		9273 => to_signed(25442, LUT_AMPL_WIDTH),
		9274 => to_signed(25444, LUT_AMPL_WIDTH),
		9275 => to_signed(25446, LUT_AMPL_WIDTH),
		9276 => to_signed(25448, LUT_AMPL_WIDTH),
		9277 => to_signed(25450, LUT_AMPL_WIDTH),
		9278 => to_signed(25452, LUT_AMPL_WIDTH),
		9279 => to_signed(25454, LUT_AMPL_WIDTH),
		9280 => to_signed(25456, LUT_AMPL_WIDTH),
		9281 => to_signed(25458, LUT_AMPL_WIDTH),
		9282 => to_signed(25460, LUT_AMPL_WIDTH),
		9283 => to_signed(25462, LUT_AMPL_WIDTH),
		9284 => to_signed(25464, LUT_AMPL_WIDTH),
		9285 => to_signed(25466, LUT_AMPL_WIDTH),
		9286 => to_signed(25468, LUT_AMPL_WIDTH),
		9287 => to_signed(25470, LUT_AMPL_WIDTH),
		9288 => to_signed(25472, LUT_AMPL_WIDTH),
		9289 => to_signed(25474, LUT_AMPL_WIDTH),
		9290 => to_signed(25476, LUT_AMPL_WIDTH),
		9291 => to_signed(25478, LUT_AMPL_WIDTH),
		9292 => to_signed(25480, LUT_AMPL_WIDTH),
		9293 => to_signed(25482, LUT_AMPL_WIDTH),
		9294 => to_signed(25484, LUT_AMPL_WIDTH),
		9295 => to_signed(25486, LUT_AMPL_WIDTH),
		9296 => to_signed(25488, LUT_AMPL_WIDTH),
		9297 => to_signed(25490, LUT_AMPL_WIDTH),
		9298 => to_signed(25492, LUT_AMPL_WIDTH),
		9299 => to_signed(25494, LUT_AMPL_WIDTH),
		9300 => to_signed(25496, LUT_AMPL_WIDTH),
		9301 => to_signed(25498, LUT_AMPL_WIDTH),
		9302 => to_signed(25500, LUT_AMPL_WIDTH),
		9303 => to_signed(25502, LUT_AMPL_WIDTH),
		9304 => to_signed(25504, LUT_AMPL_WIDTH),
		9305 => to_signed(25506, LUT_AMPL_WIDTH),
		9306 => to_signed(25508, LUT_AMPL_WIDTH),
		9307 => to_signed(25510, LUT_AMPL_WIDTH),
		9308 => to_signed(25512, LUT_AMPL_WIDTH),
		9309 => to_signed(25514, LUT_AMPL_WIDTH),
		9310 => to_signed(25516, LUT_AMPL_WIDTH),
		9311 => to_signed(25518, LUT_AMPL_WIDTH),
		9312 => to_signed(25519, LUT_AMPL_WIDTH),
		9313 => to_signed(25521, LUT_AMPL_WIDTH),
		9314 => to_signed(25523, LUT_AMPL_WIDTH),
		9315 => to_signed(25525, LUT_AMPL_WIDTH),
		9316 => to_signed(25527, LUT_AMPL_WIDTH),
		9317 => to_signed(25529, LUT_AMPL_WIDTH),
		9318 => to_signed(25531, LUT_AMPL_WIDTH),
		9319 => to_signed(25533, LUT_AMPL_WIDTH),
		9320 => to_signed(25535, LUT_AMPL_WIDTH),
		9321 => to_signed(25537, LUT_AMPL_WIDTH),
		9322 => to_signed(25539, LUT_AMPL_WIDTH),
		9323 => to_signed(25541, LUT_AMPL_WIDTH),
		9324 => to_signed(25543, LUT_AMPL_WIDTH),
		9325 => to_signed(25545, LUT_AMPL_WIDTH),
		9326 => to_signed(25547, LUT_AMPL_WIDTH),
		9327 => to_signed(25549, LUT_AMPL_WIDTH),
		9328 => to_signed(25551, LUT_AMPL_WIDTH),
		9329 => to_signed(25553, LUT_AMPL_WIDTH),
		9330 => to_signed(25555, LUT_AMPL_WIDTH),
		9331 => to_signed(25557, LUT_AMPL_WIDTH),
		9332 => to_signed(25559, LUT_AMPL_WIDTH),
		9333 => to_signed(25561, LUT_AMPL_WIDTH),
		9334 => to_signed(25563, LUT_AMPL_WIDTH),
		9335 => to_signed(25565, LUT_AMPL_WIDTH),
		9336 => to_signed(25567, LUT_AMPL_WIDTH),
		9337 => to_signed(25569, LUT_AMPL_WIDTH),
		9338 => to_signed(25571, LUT_AMPL_WIDTH),
		9339 => to_signed(25573, LUT_AMPL_WIDTH),
		9340 => to_signed(25575, LUT_AMPL_WIDTH),
		9341 => to_signed(25577, LUT_AMPL_WIDTH),
		9342 => to_signed(25578, LUT_AMPL_WIDTH),
		9343 => to_signed(25580, LUT_AMPL_WIDTH),
		9344 => to_signed(25582, LUT_AMPL_WIDTH),
		9345 => to_signed(25584, LUT_AMPL_WIDTH),
		9346 => to_signed(25586, LUT_AMPL_WIDTH),
		9347 => to_signed(25588, LUT_AMPL_WIDTH),
		9348 => to_signed(25590, LUT_AMPL_WIDTH),
		9349 => to_signed(25592, LUT_AMPL_WIDTH),
		9350 => to_signed(25594, LUT_AMPL_WIDTH),
		9351 => to_signed(25596, LUT_AMPL_WIDTH),
		9352 => to_signed(25598, LUT_AMPL_WIDTH),
		9353 => to_signed(25600, LUT_AMPL_WIDTH),
		9354 => to_signed(25602, LUT_AMPL_WIDTH),
		9355 => to_signed(25604, LUT_AMPL_WIDTH),
		9356 => to_signed(25606, LUT_AMPL_WIDTH),
		9357 => to_signed(25608, LUT_AMPL_WIDTH),
		9358 => to_signed(25610, LUT_AMPL_WIDTH),
		9359 => to_signed(25612, LUT_AMPL_WIDTH),
		9360 => to_signed(25614, LUT_AMPL_WIDTH),
		9361 => to_signed(25616, LUT_AMPL_WIDTH),
		9362 => to_signed(25618, LUT_AMPL_WIDTH),
		9363 => to_signed(25620, LUT_AMPL_WIDTH),
		9364 => to_signed(25622, LUT_AMPL_WIDTH),
		9365 => to_signed(25624, LUT_AMPL_WIDTH),
		9366 => to_signed(25626, LUT_AMPL_WIDTH),
		9367 => to_signed(25628, LUT_AMPL_WIDTH),
		9368 => to_signed(25629, LUT_AMPL_WIDTH),
		9369 => to_signed(25631, LUT_AMPL_WIDTH),
		9370 => to_signed(25633, LUT_AMPL_WIDTH),
		9371 => to_signed(25635, LUT_AMPL_WIDTH),
		9372 => to_signed(25637, LUT_AMPL_WIDTH),
		9373 => to_signed(25639, LUT_AMPL_WIDTH),
		9374 => to_signed(25641, LUT_AMPL_WIDTH),
		9375 => to_signed(25643, LUT_AMPL_WIDTH),
		9376 => to_signed(25645, LUT_AMPL_WIDTH),
		9377 => to_signed(25647, LUT_AMPL_WIDTH),
		9378 => to_signed(25649, LUT_AMPL_WIDTH),
		9379 => to_signed(25651, LUT_AMPL_WIDTH),
		9380 => to_signed(25653, LUT_AMPL_WIDTH),
		9381 => to_signed(25655, LUT_AMPL_WIDTH),
		9382 => to_signed(25657, LUT_AMPL_WIDTH),
		9383 => to_signed(25659, LUT_AMPL_WIDTH),
		9384 => to_signed(25661, LUT_AMPL_WIDTH),
		9385 => to_signed(25663, LUT_AMPL_WIDTH),
		9386 => to_signed(25665, LUT_AMPL_WIDTH),
		9387 => to_signed(25667, LUT_AMPL_WIDTH),
		9388 => to_signed(25669, LUT_AMPL_WIDTH),
		9389 => to_signed(25671, LUT_AMPL_WIDTH),
		9390 => to_signed(25672, LUT_AMPL_WIDTH),
		9391 => to_signed(25674, LUT_AMPL_WIDTH),
		9392 => to_signed(25676, LUT_AMPL_WIDTH),
		9393 => to_signed(25678, LUT_AMPL_WIDTH),
		9394 => to_signed(25680, LUT_AMPL_WIDTH),
		9395 => to_signed(25682, LUT_AMPL_WIDTH),
		9396 => to_signed(25684, LUT_AMPL_WIDTH),
		9397 => to_signed(25686, LUT_AMPL_WIDTH),
		9398 => to_signed(25688, LUT_AMPL_WIDTH),
		9399 => to_signed(25690, LUT_AMPL_WIDTH),
		9400 => to_signed(25692, LUT_AMPL_WIDTH),
		9401 => to_signed(25694, LUT_AMPL_WIDTH),
		9402 => to_signed(25696, LUT_AMPL_WIDTH),
		9403 => to_signed(25698, LUT_AMPL_WIDTH),
		9404 => to_signed(25700, LUT_AMPL_WIDTH),
		9405 => to_signed(25702, LUT_AMPL_WIDTH),
		9406 => to_signed(25704, LUT_AMPL_WIDTH),
		9407 => to_signed(25706, LUT_AMPL_WIDTH),
		9408 => to_signed(25708, LUT_AMPL_WIDTH),
		9409 => to_signed(25710, LUT_AMPL_WIDTH),
		9410 => to_signed(25711, LUT_AMPL_WIDTH),
		9411 => to_signed(25713, LUT_AMPL_WIDTH),
		9412 => to_signed(25715, LUT_AMPL_WIDTH),
		9413 => to_signed(25717, LUT_AMPL_WIDTH),
		9414 => to_signed(25719, LUT_AMPL_WIDTH),
		9415 => to_signed(25721, LUT_AMPL_WIDTH),
		9416 => to_signed(25723, LUT_AMPL_WIDTH),
		9417 => to_signed(25725, LUT_AMPL_WIDTH),
		9418 => to_signed(25727, LUT_AMPL_WIDTH),
		9419 => to_signed(25729, LUT_AMPL_WIDTH),
		9420 => to_signed(25731, LUT_AMPL_WIDTH),
		9421 => to_signed(25733, LUT_AMPL_WIDTH),
		9422 => to_signed(25735, LUT_AMPL_WIDTH),
		9423 => to_signed(25737, LUT_AMPL_WIDTH),
		9424 => to_signed(25739, LUT_AMPL_WIDTH),
		9425 => to_signed(25741, LUT_AMPL_WIDTH),
		9426 => to_signed(25743, LUT_AMPL_WIDTH),
		9427 => to_signed(25745, LUT_AMPL_WIDTH),
		9428 => to_signed(25746, LUT_AMPL_WIDTH),
		9429 => to_signed(25748, LUT_AMPL_WIDTH),
		9430 => to_signed(25750, LUT_AMPL_WIDTH),
		9431 => to_signed(25752, LUT_AMPL_WIDTH),
		9432 => to_signed(25754, LUT_AMPL_WIDTH),
		9433 => to_signed(25756, LUT_AMPL_WIDTH),
		9434 => to_signed(25758, LUT_AMPL_WIDTH),
		9435 => to_signed(25760, LUT_AMPL_WIDTH),
		9436 => to_signed(25762, LUT_AMPL_WIDTH),
		9437 => to_signed(25764, LUT_AMPL_WIDTH),
		9438 => to_signed(25766, LUT_AMPL_WIDTH),
		9439 => to_signed(25768, LUT_AMPL_WIDTH),
		9440 => to_signed(25770, LUT_AMPL_WIDTH),
		9441 => to_signed(25772, LUT_AMPL_WIDTH),
		9442 => to_signed(25774, LUT_AMPL_WIDTH),
		9443 => to_signed(25776, LUT_AMPL_WIDTH),
		9444 => to_signed(25778, LUT_AMPL_WIDTH),
		9445 => to_signed(25779, LUT_AMPL_WIDTH),
		9446 => to_signed(25781, LUT_AMPL_WIDTH),
		9447 => to_signed(25783, LUT_AMPL_WIDTH),
		9448 => to_signed(25785, LUT_AMPL_WIDTH),
		9449 => to_signed(25787, LUT_AMPL_WIDTH),
		9450 => to_signed(25789, LUT_AMPL_WIDTH),
		9451 => to_signed(25791, LUT_AMPL_WIDTH),
		9452 => to_signed(25793, LUT_AMPL_WIDTH),
		9453 => to_signed(25795, LUT_AMPL_WIDTH),
		9454 => to_signed(25797, LUT_AMPL_WIDTH),
		9455 => to_signed(25799, LUT_AMPL_WIDTH),
		9456 => to_signed(25801, LUT_AMPL_WIDTH),
		9457 => to_signed(25803, LUT_AMPL_WIDTH),
		9458 => to_signed(25805, LUT_AMPL_WIDTH),
		9459 => to_signed(25807, LUT_AMPL_WIDTH),
		9460 => to_signed(25809, LUT_AMPL_WIDTH),
		9461 => to_signed(25810, LUT_AMPL_WIDTH),
		9462 => to_signed(25812, LUT_AMPL_WIDTH),
		9463 => to_signed(25814, LUT_AMPL_WIDTH),
		9464 => to_signed(25816, LUT_AMPL_WIDTH),
		9465 => to_signed(25818, LUT_AMPL_WIDTH),
		9466 => to_signed(25820, LUT_AMPL_WIDTH),
		9467 => to_signed(25822, LUT_AMPL_WIDTH),
		9468 => to_signed(25824, LUT_AMPL_WIDTH),
		9469 => to_signed(25826, LUT_AMPL_WIDTH),
		9470 => to_signed(25828, LUT_AMPL_WIDTH),
		9471 => to_signed(25830, LUT_AMPL_WIDTH),
		9472 => to_signed(25832, LUT_AMPL_WIDTH),
		9473 => to_signed(25834, LUT_AMPL_WIDTH),
		9474 => to_signed(25836, LUT_AMPL_WIDTH),
		9475 => to_signed(25838, LUT_AMPL_WIDTH),
		9476 => to_signed(25839, LUT_AMPL_WIDTH),
		9477 => to_signed(25841, LUT_AMPL_WIDTH),
		9478 => to_signed(25843, LUT_AMPL_WIDTH),
		9479 => to_signed(25845, LUT_AMPL_WIDTH),
		9480 => to_signed(25847, LUT_AMPL_WIDTH),
		9481 => to_signed(25849, LUT_AMPL_WIDTH),
		9482 => to_signed(25851, LUT_AMPL_WIDTH),
		9483 => to_signed(25853, LUT_AMPL_WIDTH),
		9484 => to_signed(25855, LUT_AMPL_WIDTH),
		9485 => to_signed(25857, LUT_AMPL_WIDTH),
		9486 => to_signed(25859, LUT_AMPL_WIDTH),
		9487 => to_signed(25861, LUT_AMPL_WIDTH),
		9488 => to_signed(25863, LUT_AMPL_WIDTH),
		9489 => to_signed(25865, LUT_AMPL_WIDTH),
		9490 => to_signed(25866, LUT_AMPL_WIDTH),
		9491 => to_signed(25868, LUT_AMPL_WIDTH),
		9492 => to_signed(25870, LUT_AMPL_WIDTH),
		9493 => to_signed(25872, LUT_AMPL_WIDTH),
		9494 => to_signed(25874, LUT_AMPL_WIDTH),
		9495 => to_signed(25876, LUT_AMPL_WIDTH),
		9496 => to_signed(25878, LUT_AMPL_WIDTH),
		9497 => to_signed(25880, LUT_AMPL_WIDTH),
		9498 => to_signed(25882, LUT_AMPL_WIDTH),
		9499 => to_signed(25884, LUT_AMPL_WIDTH),
		9500 => to_signed(25886, LUT_AMPL_WIDTH),
		9501 => to_signed(25888, LUT_AMPL_WIDTH),
		9502 => to_signed(25890, LUT_AMPL_WIDTH),
		9503 => to_signed(25892, LUT_AMPL_WIDTH),
		9504 => to_signed(25893, LUT_AMPL_WIDTH),
		9505 => to_signed(25895, LUT_AMPL_WIDTH),
		9506 => to_signed(25897, LUT_AMPL_WIDTH),
		9507 => to_signed(25899, LUT_AMPL_WIDTH),
		9508 => to_signed(25901, LUT_AMPL_WIDTH),
		9509 => to_signed(25903, LUT_AMPL_WIDTH),
		9510 => to_signed(25905, LUT_AMPL_WIDTH),
		9511 => to_signed(25907, LUT_AMPL_WIDTH),
		9512 => to_signed(25909, LUT_AMPL_WIDTH),
		9513 => to_signed(25911, LUT_AMPL_WIDTH),
		9514 => to_signed(25913, LUT_AMPL_WIDTH),
		9515 => to_signed(25915, LUT_AMPL_WIDTH),
		9516 => to_signed(25917, LUT_AMPL_WIDTH),
		9517 => to_signed(25918, LUT_AMPL_WIDTH),
		9518 => to_signed(25920, LUT_AMPL_WIDTH),
		9519 => to_signed(25922, LUT_AMPL_WIDTH),
		9520 => to_signed(25924, LUT_AMPL_WIDTH),
		9521 => to_signed(25926, LUT_AMPL_WIDTH),
		9522 => to_signed(25928, LUT_AMPL_WIDTH),
		9523 => to_signed(25930, LUT_AMPL_WIDTH),
		9524 => to_signed(25932, LUT_AMPL_WIDTH),
		9525 => to_signed(25934, LUT_AMPL_WIDTH),
		9526 => to_signed(25936, LUT_AMPL_WIDTH),
		9527 => to_signed(25938, LUT_AMPL_WIDTH),
		9528 => to_signed(25940, LUT_AMPL_WIDTH),
		9529 => to_signed(25942, LUT_AMPL_WIDTH),
		9530 => to_signed(25943, LUT_AMPL_WIDTH),
		9531 => to_signed(25945, LUT_AMPL_WIDTH),
		9532 => to_signed(25947, LUT_AMPL_WIDTH),
		9533 => to_signed(25949, LUT_AMPL_WIDTH),
		9534 => to_signed(25951, LUT_AMPL_WIDTH),
		9535 => to_signed(25953, LUT_AMPL_WIDTH),
		9536 => to_signed(25955, LUT_AMPL_WIDTH),
		9537 => to_signed(25957, LUT_AMPL_WIDTH),
		9538 => to_signed(25959, LUT_AMPL_WIDTH),
		9539 => to_signed(25961, LUT_AMPL_WIDTH),
		9540 => to_signed(25963, LUT_AMPL_WIDTH),
		9541 => to_signed(25965, LUT_AMPL_WIDTH),
		9542 => to_signed(25966, LUT_AMPL_WIDTH),
		9543 => to_signed(25968, LUT_AMPL_WIDTH),
		9544 => to_signed(25970, LUT_AMPL_WIDTH),
		9545 => to_signed(25972, LUT_AMPL_WIDTH),
		9546 => to_signed(25974, LUT_AMPL_WIDTH),
		9547 => to_signed(25976, LUT_AMPL_WIDTH),
		9548 => to_signed(25978, LUT_AMPL_WIDTH),
		9549 => to_signed(25980, LUT_AMPL_WIDTH),
		9550 => to_signed(25982, LUT_AMPL_WIDTH),
		9551 => to_signed(25984, LUT_AMPL_WIDTH),
		9552 => to_signed(25986, LUT_AMPL_WIDTH),
		9553 => to_signed(25988, LUT_AMPL_WIDTH),
		9554 => to_signed(25989, LUT_AMPL_WIDTH),
		9555 => to_signed(25991, LUT_AMPL_WIDTH),
		9556 => to_signed(25993, LUT_AMPL_WIDTH),
		9557 => to_signed(25995, LUT_AMPL_WIDTH),
		9558 => to_signed(25997, LUT_AMPL_WIDTH),
		9559 => to_signed(25999, LUT_AMPL_WIDTH),
		9560 => to_signed(26001, LUT_AMPL_WIDTH),
		9561 => to_signed(26003, LUT_AMPL_WIDTH),
		9562 => to_signed(26005, LUT_AMPL_WIDTH),
		9563 => to_signed(26007, LUT_AMPL_WIDTH),
		9564 => to_signed(26009, LUT_AMPL_WIDTH),
		9565 => to_signed(26010, LUT_AMPL_WIDTH),
		9566 => to_signed(26012, LUT_AMPL_WIDTH),
		9567 => to_signed(26014, LUT_AMPL_WIDTH),
		9568 => to_signed(26016, LUT_AMPL_WIDTH),
		9569 => to_signed(26018, LUT_AMPL_WIDTH),
		9570 => to_signed(26020, LUT_AMPL_WIDTH),
		9571 => to_signed(26022, LUT_AMPL_WIDTH),
		9572 => to_signed(26024, LUT_AMPL_WIDTH),
		9573 => to_signed(26026, LUT_AMPL_WIDTH),
		9574 => to_signed(26028, LUT_AMPL_WIDTH),
		9575 => to_signed(26030, LUT_AMPL_WIDTH),
		9576 => to_signed(26031, LUT_AMPL_WIDTH),
		9577 => to_signed(26033, LUT_AMPL_WIDTH),
		9578 => to_signed(26035, LUT_AMPL_WIDTH),
		9579 => to_signed(26037, LUT_AMPL_WIDTH),
		9580 => to_signed(26039, LUT_AMPL_WIDTH),
		9581 => to_signed(26041, LUT_AMPL_WIDTH),
		9582 => to_signed(26043, LUT_AMPL_WIDTH),
		9583 => to_signed(26045, LUT_AMPL_WIDTH),
		9584 => to_signed(26047, LUT_AMPL_WIDTH),
		9585 => to_signed(26049, LUT_AMPL_WIDTH),
		9586 => to_signed(26051, LUT_AMPL_WIDTH),
		9587 => to_signed(26052, LUT_AMPL_WIDTH),
		9588 => to_signed(26054, LUT_AMPL_WIDTH),
		9589 => to_signed(26056, LUT_AMPL_WIDTH),
		9590 => to_signed(26058, LUT_AMPL_WIDTH),
		9591 => to_signed(26060, LUT_AMPL_WIDTH),
		9592 => to_signed(26062, LUT_AMPL_WIDTH),
		9593 => to_signed(26064, LUT_AMPL_WIDTH),
		9594 => to_signed(26066, LUT_AMPL_WIDTH),
		9595 => to_signed(26068, LUT_AMPL_WIDTH),
		9596 => to_signed(26070, LUT_AMPL_WIDTH),
		9597 => to_signed(26071, LUT_AMPL_WIDTH),
		9598 => to_signed(26073, LUT_AMPL_WIDTH),
		9599 => to_signed(26075, LUT_AMPL_WIDTH),
		9600 => to_signed(26077, LUT_AMPL_WIDTH),
		9601 => to_signed(26079, LUT_AMPL_WIDTH),
		9602 => to_signed(26081, LUT_AMPL_WIDTH),
		9603 => to_signed(26083, LUT_AMPL_WIDTH),
		9604 => to_signed(26085, LUT_AMPL_WIDTH),
		9605 => to_signed(26087, LUT_AMPL_WIDTH),
		9606 => to_signed(26089, LUT_AMPL_WIDTH),
		9607 => to_signed(26090, LUT_AMPL_WIDTH),
		9608 => to_signed(26092, LUT_AMPL_WIDTH),
		9609 => to_signed(26094, LUT_AMPL_WIDTH),
		9610 => to_signed(26096, LUT_AMPL_WIDTH),
		9611 => to_signed(26098, LUT_AMPL_WIDTH),
		9612 => to_signed(26100, LUT_AMPL_WIDTH),
		9613 => to_signed(26102, LUT_AMPL_WIDTH),
		9614 => to_signed(26104, LUT_AMPL_WIDTH),
		9615 => to_signed(26106, LUT_AMPL_WIDTH),
		9616 => to_signed(26108, LUT_AMPL_WIDTH),
		9617 => to_signed(26109, LUT_AMPL_WIDTH),
		9618 => to_signed(26111, LUT_AMPL_WIDTH),
		9619 => to_signed(26113, LUT_AMPL_WIDTH),
		9620 => to_signed(26115, LUT_AMPL_WIDTH),
		9621 => to_signed(26117, LUT_AMPL_WIDTH),
		9622 => to_signed(26119, LUT_AMPL_WIDTH),
		9623 => to_signed(26121, LUT_AMPL_WIDTH),
		9624 => to_signed(26123, LUT_AMPL_WIDTH),
		9625 => to_signed(26125, LUT_AMPL_WIDTH),
		9626 => to_signed(26127, LUT_AMPL_WIDTH),
		9627 => to_signed(26128, LUT_AMPL_WIDTH),
		9628 => to_signed(26130, LUT_AMPL_WIDTH),
		9629 => to_signed(26132, LUT_AMPL_WIDTH),
		9630 => to_signed(26134, LUT_AMPL_WIDTH),
		9631 => to_signed(26136, LUT_AMPL_WIDTH),
		9632 => to_signed(26138, LUT_AMPL_WIDTH),
		9633 => to_signed(26140, LUT_AMPL_WIDTH),
		9634 => to_signed(26142, LUT_AMPL_WIDTH),
		9635 => to_signed(26144, LUT_AMPL_WIDTH),
		9636 => to_signed(26146, LUT_AMPL_WIDTH),
		9637 => to_signed(26147, LUT_AMPL_WIDTH),
		9638 => to_signed(26149, LUT_AMPL_WIDTH),
		9639 => to_signed(26151, LUT_AMPL_WIDTH),
		9640 => to_signed(26153, LUT_AMPL_WIDTH),
		9641 => to_signed(26155, LUT_AMPL_WIDTH),
		9642 => to_signed(26157, LUT_AMPL_WIDTH),
		9643 => to_signed(26159, LUT_AMPL_WIDTH),
		9644 => to_signed(26161, LUT_AMPL_WIDTH),
		9645 => to_signed(26163, LUT_AMPL_WIDTH),
		9646 => to_signed(26164, LUT_AMPL_WIDTH),
		9647 => to_signed(26166, LUT_AMPL_WIDTH),
		9648 => to_signed(26168, LUT_AMPL_WIDTH),
		9649 => to_signed(26170, LUT_AMPL_WIDTH),
		9650 => to_signed(26172, LUT_AMPL_WIDTH),
		9651 => to_signed(26174, LUT_AMPL_WIDTH),
		9652 => to_signed(26176, LUT_AMPL_WIDTH),
		9653 => to_signed(26178, LUT_AMPL_WIDTH),
		9654 => to_signed(26180, LUT_AMPL_WIDTH),
		9655 => to_signed(26181, LUT_AMPL_WIDTH),
		9656 => to_signed(26183, LUT_AMPL_WIDTH),
		9657 => to_signed(26185, LUT_AMPL_WIDTH),
		9658 => to_signed(26187, LUT_AMPL_WIDTH),
		9659 => to_signed(26189, LUT_AMPL_WIDTH),
		9660 => to_signed(26191, LUT_AMPL_WIDTH),
		9661 => to_signed(26193, LUT_AMPL_WIDTH),
		9662 => to_signed(26195, LUT_AMPL_WIDTH),
		9663 => to_signed(26197, LUT_AMPL_WIDTH),
		9664 => to_signed(26198, LUT_AMPL_WIDTH),
		9665 => to_signed(26200, LUT_AMPL_WIDTH),
		9666 => to_signed(26202, LUT_AMPL_WIDTH),
		9667 => to_signed(26204, LUT_AMPL_WIDTH),
		9668 => to_signed(26206, LUT_AMPL_WIDTH),
		9669 => to_signed(26208, LUT_AMPL_WIDTH),
		9670 => to_signed(26210, LUT_AMPL_WIDTH),
		9671 => to_signed(26212, LUT_AMPL_WIDTH),
		9672 => to_signed(26214, LUT_AMPL_WIDTH),
		9673 => to_signed(26215, LUT_AMPL_WIDTH),
		9674 => to_signed(26217, LUT_AMPL_WIDTH),
		9675 => to_signed(26219, LUT_AMPL_WIDTH),
		9676 => to_signed(26221, LUT_AMPL_WIDTH),
		9677 => to_signed(26223, LUT_AMPL_WIDTH),
		9678 => to_signed(26225, LUT_AMPL_WIDTH),
		9679 => to_signed(26227, LUT_AMPL_WIDTH),
		9680 => to_signed(26229, LUT_AMPL_WIDTH),
		9681 => to_signed(26230, LUT_AMPL_WIDTH),
		9682 => to_signed(26232, LUT_AMPL_WIDTH),
		9683 => to_signed(26234, LUT_AMPL_WIDTH),
		9684 => to_signed(26236, LUT_AMPL_WIDTH),
		9685 => to_signed(26238, LUT_AMPL_WIDTH),
		9686 => to_signed(26240, LUT_AMPL_WIDTH),
		9687 => to_signed(26242, LUT_AMPL_WIDTH),
		9688 => to_signed(26244, LUT_AMPL_WIDTH),
		9689 => to_signed(26246, LUT_AMPL_WIDTH),
		9690 => to_signed(26247, LUT_AMPL_WIDTH),
		9691 => to_signed(26249, LUT_AMPL_WIDTH),
		9692 => to_signed(26251, LUT_AMPL_WIDTH),
		9693 => to_signed(26253, LUT_AMPL_WIDTH),
		9694 => to_signed(26255, LUT_AMPL_WIDTH),
		9695 => to_signed(26257, LUT_AMPL_WIDTH),
		9696 => to_signed(26259, LUT_AMPL_WIDTH),
		9697 => to_signed(26261, LUT_AMPL_WIDTH),
		9698 => to_signed(26262, LUT_AMPL_WIDTH),
		9699 => to_signed(26264, LUT_AMPL_WIDTH),
		9700 => to_signed(26266, LUT_AMPL_WIDTH),
		9701 => to_signed(26268, LUT_AMPL_WIDTH),
		9702 => to_signed(26270, LUT_AMPL_WIDTH),
		9703 => to_signed(26272, LUT_AMPL_WIDTH),
		9704 => to_signed(26274, LUT_AMPL_WIDTH),
		9705 => to_signed(26276, LUT_AMPL_WIDTH),
		9706 => to_signed(26277, LUT_AMPL_WIDTH),
		9707 => to_signed(26279, LUT_AMPL_WIDTH),
		9708 => to_signed(26281, LUT_AMPL_WIDTH),
		9709 => to_signed(26283, LUT_AMPL_WIDTH),
		9710 => to_signed(26285, LUT_AMPL_WIDTH),
		9711 => to_signed(26287, LUT_AMPL_WIDTH),
		9712 => to_signed(26289, LUT_AMPL_WIDTH),
		9713 => to_signed(26291, LUT_AMPL_WIDTH),
		9714 => to_signed(26292, LUT_AMPL_WIDTH),
		9715 => to_signed(26294, LUT_AMPL_WIDTH),
		9716 => to_signed(26296, LUT_AMPL_WIDTH),
		9717 => to_signed(26298, LUT_AMPL_WIDTH),
		9718 => to_signed(26300, LUT_AMPL_WIDTH),
		9719 => to_signed(26302, LUT_AMPL_WIDTH),
		9720 => to_signed(26304, LUT_AMPL_WIDTH),
		9721 => to_signed(26306, LUT_AMPL_WIDTH),
		9722 => to_signed(26307, LUT_AMPL_WIDTH),
		9723 => to_signed(26309, LUT_AMPL_WIDTH),
		9724 => to_signed(26311, LUT_AMPL_WIDTH),
		9725 => to_signed(26313, LUT_AMPL_WIDTH),
		9726 => to_signed(26315, LUT_AMPL_WIDTH),
		9727 => to_signed(26317, LUT_AMPL_WIDTH),
		9728 => to_signed(26319, LUT_AMPL_WIDTH),
		9729 => to_signed(26321, LUT_AMPL_WIDTH),
		9730 => to_signed(26322, LUT_AMPL_WIDTH),
		9731 => to_signed(26324, LUT_AMPL_WIDTH),
		9732 => to_signed(26326, LUT_AMPL_WIDTH),
		9733 => to_signed(26328, LUT_AMPL_WIDTH),
		9734 => to_signed(26330, LUT_AMPL_WIDTH),
		9735 => to_signed(26332, LUT_AMPL_WIDTH),
		9736 => to_signed(26334, LUT_AMPL_WIDTH),
		9737 => to_signed(26336, LUT_AMPL_WIDTH),
		9738 => to_signed(26337, LUT_AMPL_WIDTH),
		9739 => to_signed(26339, LUT_AMPL_WIDTH),
		9740 => to_signed(26341, LUT_AMPL_WIDTH),
		9741 => to_signed(26343, LUT_AMPL_WIDTH),
		9742 => to_signed(26345, LUT_AMPL_WIDTH),
		9743 => to_signed(26347, LUT_AMPL_WIDTH),
		9744 => to_signed(26349, LUT_AMPL_WIDTH),
		9745 => to_signed(26350, LUT_AMPL_WIDTH),
		9746 => to_signed(26352, LUT_AMPL_WIDTH),
		9747 => to_signed(26354, LUT_AMPL_WIDTH),
		9748 => to_signed(26356, LUT_AMPL_WIDTH),
		9749 => to_signed(26358, LUT_AMPL_WIDTH),
		9750 => to_signed(26360, LUT_AMPL_WIDTH),
		9751 => to_signed(26362, LUT_AMPL_WIDTH),
		9752 => to_signed(26364, LUT_AMPL_WIDTH),
		9753 => to_signed(26365, LUT_AMPL_WIDTH),
		9754 => to_signed(26367, LUT_AMPL_WIDTH),
		9755 => to_signed(26369, LUT_AMPL_WIDTH),
		9756 => to_signed(26371, LUT_AMPL_WIDTH),
		9757 => to_signed(26373, LUT_AMPL_WIDTH),
		9758 => to_signed(26375, LUT_AMPL_WIDTH),
		9759 => to_signed(26377, LUT_AMPL_WIDTH),
		9760 => to_signed(26378, LUT_AMPL_WIDTH),
		9761 => to_signed(26380, LUT_AMPL_WIDTH),
		9762 => to_signed(26382, LUT_AMPL_WIDTH),
		9763 => to_signed(26384, LUT_AMPL_WIDTH),
		9764 => to_signed(26386, LUT_AMPL_WIDTH),
		9765 => to_signed(26388, LUT_AMPL_WIDTH),
		9766 => to_signed(26390, LUT_AMPL_WIDTH),
		9767 => to_signed(26392, LUT_AMPL_WIDTH),
		9768 => to_signed(26393, LUT_AMPL_WIDTH),
		9769 => to_signed(26395, LUT_AMPL_WIDTH),
		9770 => to_signed(26397, LUT_AMPL_WIDTH),
		9771 => to_signed(26399, LUT_AMPL_WIDTH),
		9772 => to_signed(26401, LUT_AMPL_WIDTH),
		9773 => to_signed(26403, LUT_AMPL_WIDTH),
		9774 => to_signed(26405, LUT_AMPL_WIDTH),
		9775 => to_signed(26406, LUT_AMPL_WIDTH),
		9776 => to_signed(26408, LUT_AMPL_WIDTH),
		9777 => to_signed(26410, LUT_AMPL_WIDTH),
		9778 => to_signed(26412, LUT_AMPL_WIDTH),
		9779 => to_signed(26414, LUT_AMPL_WIDTH),
		9780 => to_signed(26416, LUT_AMPL_WIDTH),
		9781 => to_signed(26418, LUT_AMPL_WIDTH),
		9782 => to_signed(26419, LUT_AMPL_WIDTH),
		9783 => to_signed(26421, LUT_AMPL_WIDTH),
		9784 => to_signed(26423, LUT_AMPL_WIDTH),
		9785 => to_signed(26425, LUT_AMPL_WIDTH),
		9786 => to_signed(26427, LUT_AMPL_WIDTH),
		9787 => to_signed(26429, LUT_AMPL_WIDTH),
		9788 => to_signed(26431, LUT_AMPL_WIDTH),
		9789 => to_signed(26432, LUT_AMPL_WIDTH),
		9790 => to_signed(26434, LUT_AMPL_WIDTH),
		9791 => to_signed(26436, LUT_AMPL_WIDTH),
		9792 => to_signed(26438, LUT_AMPL_WIDTH),
		9793 => to_signed(26440, LUT_AMPL_WIDTH),
		9794 => to_signed(26442, LUT_AMPL_WIDTH),
		9795 => to_signed(26444, LUT_AMPL_WIDTH),
		9796 => to_signed(26445, LUT_AMPL_WIDTH),
		9797 => to_signed(26447, LUT_AMPL_WIDTH),
		9798 => to_signed(26449, LUT_AMPL_WIDTH),
		9799 => to_signed(26451, LUT_AMPL_WIDTH),
		9800 => to_signed(26453, LUT_AMPL_WIDTH),
		9801 => to_signed(26455, LUT_AMPL_WIDTH),
		9802 => to_signed(26457, LUT_AMPL_WIDTH),
		9803 => to_signed(26458, LUT_AMPL_WIDTH),
		9804 => to_signed(26460, LUT_AMPL_WIDTH),
		9805 => to_signed(26462, LUT_AMPL_WIDTH),
		9806 => to_signed(26464, LUT_AMPL_WIDTH),
		9807 => to_signed(26466, LUT_AMPL_WIDTH),
		9808 => to_signed(26468, LUT_AMPL_WIDTH),
		9809 => to_signed(26469, LUT_AMPL_WIDTH),
		9810 => to_signed(26471, LUT_AMPL_WIDTH),
		9811 => to_signed(26473, LUT_AMPL_WIDTH),
		9812 => to_signed(26475, LUT_AMPL_WIDTH),
		9813 => to_signed(26477, LUT_AMPL_WIDTH),
		9814 => to_signed(26479, LUT_AMPL_WIDTH),
		9815 => to_signed(26481, LUT_AMPL_WIDTH),
		9816 => to_signed(26482, LUT_AMPL_WIDTH),
		9817 => to_signed(26484, LUT_AMPL_WIDTH),
		9818 => to_signed(26486, LUT_AMPL_WIDTH),
		9819 => to_signed(26488, LUT_AMPL_WIDTH),
		9820 => to_signed(26490, LUT_AMPL_WIDTH),
		9821 => to_signed(26492, LUT_AMPL_WIDTH),
		9822 => to_signed(26494, LUT_AMPL_WIDTH),
		9823 => to_signed(26495, LUT_AMPL_WIDTH),
		9824 => to_signed(26497, LUT_AMPL_WIDTH),
		9825 => to_signed(26499, LUT_AMPL_WIDTH),
		9826 => to_signed(26501, LUT_AMPL_WIDTH),
		9827 => to_signed(26503, LUT_AMPL_WIDTH),
		9828 => to_signed(26505, LUT_AMPL_WIDTH),
		9829 => to_signed(26506, LUT_AMPL_WIDTH),
		9830 => to_signed(26508, LUT_AMPL_WIDTH),
		9831 => to_signed(26510, LUT_AMPL_WIDTH),
		9832 => to_signed(26512, LUT_AMPL_WIDTH),
		9833 => to_signed(26514, LUT_AMPL_WIDTH),
		9834 => to_signed(26516, LUT_AMPL_WIDTH),
		9835 => to_signed(26518, LUT_AMPL_WIDTH),
		9836 => to_signed(26519, LUT_AMPL_WIDTH),
		9837 => to_signed(26521, LUT_AMPL_WIDTH),
		9838 => to_signed(26523, LUT_AMPL_WIDTH),
		9839 => to_signed(26525, LUT_AMPL_WIDTH),
		9840 => to_signed(26527, LUT_AMPL_WIDTH),
		9841 => to_signed(26529, LUT_AMPL_WIDTH),
		9842 => to_signed(26530, LUT_AMPL_WIDTH),
		9843 => to_signed(26532, LUT_AMPL_WIDTH),
		9844 => to_signed(26534, LUT_AMPL_WIDTH),
		9845 => to_signed(26536, LUT_AMPL_WIDTH),
		9846 => to_signed(26538, LUT_AMPL_WIDTH),
		9847 => to_signed(26540, LUT_AMPL_WIDTH),
		9848 => to_signed(26542, LUT_AMPL_WIDTH),
		9849 => to_signed(26543, LUT_AMPL_WIDTH),
		9850 => to_signed(26545, LUT_AMPL_WIDTH),
		9851 => to_signed(26547, LUT_AMPL_WIDTH),
		9852 => to_signed(26549, LUT_AMPL_WIDTH),
		9853 => to_signed(26551, LUT_AMPL_WIDTH),
		9854 => to_signed(26553, LUT_AMPL_WIDTH),
		9855 => to_signed(26554, LUT_AMPL_WIDTH),
		9856 => to_signed(26556, LUT_AMPL_WIDTH),
		9857 => to_signed(26558, LUT_AMPL_WIDTH),
		9858 => to_signed(26560, LUT_AMPL_WIDTH),
		9859 => to_signed(26562, LUT_AMPL_WIDTH),
		9860 => to_signed(26564, LUT_AMPL_WIDTH),
		9861 => to_signed(26565, LUT_AMPL_WIDTH),
		9862 => to_signed(26567, LUT_AMPL_WIDTH),
		9863 => to_signed(26569, LUT_AMPL_WIDTH),
		9864 => to_signed(26571, LUT_AMPL_WIDTH),
		9865 => to_signed(26573, LUT_AMPL_WIDTH),
		9866 => to_signed(26575, LUT_AMPL_WIDTH),
		9867 => to_signed(26576, LUT_AMPL_WIDTH),
		9868 => to_signed(26578, LUT_AMPL_WIDTH),
		9869 => to_signed(26580, LUT_AMPL_WIDTH),
		9870 => to_signed(26582, LUT_AMPL_WIDTH),
		9871 => to_signed(26584, LUT_AMPL_WIDTH),
		9872 => to_signed(26586, LUT_AMPL_WIDTH),
		9873 => to_signed(26588, LUT_AMPL_WIDTH),
		9874 => to_signed(26589, LUT_AMPL_WIDTH),
		9875 => to_signed(26591, LUT_AMPL_WIDTH),
		9876 => to_signed(26593, LUT_AMPL_WIDTH),
		9877 => to_signed(26595, LUT_AMPL_WIDTH),
		9878 => to_signed(26597, LUT_AMPL_WIDTH),
		9879 => to_signed(26599, LUT_AMPL_WIDTH),
		9880 => to_signed(26600, LUT_AMPL_WIDTH),
		9881 => to_signed(26602, LUT_AMPL_WIDTH),
		9882 => to_signed(26604, LUT_AMPL_WIDTH),
		9883 => to_signed(26606, LUT_AMPL_WIDTH),
		9884 => to_signed(26608, LUT_AMPL_WIDTH),
		9885 => to_signed(26610, LUT_AMPL_WIDTH),
		9886 => to_signed(26611, LUT_AMPL_WIDTH),
		9887 => to_signed(26613, LUT_AMPL_WIDTH),
		9888 => to_signed(26615, LUT_AMPL_WIDTH),
		9889 => to_signed(26617, LUT_AMPL_WIDTH),
		9890 => to_signed(26619, LUT_AMPL_WIDTH),
		9891 => to_signed(26621, LUT_AMPL_WIDTH),
		9892 => to_signed(26622, LUT_AMPL_WIDTH),
		9893 => to_signed(26624, LUT_AMPL_WIDTH),
		9894 => to_signed(26626, LUT_AMPL_WIDTH),
		9895 => to_signed(26628, LUT_AMPL_WIDTH),
		9896 => to_signed(26630, LUT_AMPL_WIDTH),
		9897 => to_signed(26631, LUT_AMPL_WIDTH),
		9898 => to_signed(26633, LUT_AMPL_WIDTH),
		9899 => to_signed(26635, LUT_AMPL_WIDTH),
		9900 => to_signed(26637, LUT_AMPL_WIDTH),
		9901 => to_signed(26639, LUT_AMPL_WIDTH),
		9902 => to_signed(26641, LUT_AMPL_WIDTH),
		9903 => to_signed(26642, LUT_AMPL_WIDTH),
		9904 => to_signed(26644, LUT_AMPL_WIDTH),
		9905 => to_signed(26646, LUT_AMPL_WIDTH),
		9906 => to_signed(26648, LUT_AMPL_WIDTH),
		9907 => to_signed(26650, LUT_AMPL_WIDTH),
		9908 => to_signed(26652, LUT_AMPL_WIDTH),
		9909 => to_signed(26653, LUT_AMPL_WIDTH),
		9910 => to_signed(26655, LUT_AMPL_WIDTH),
		9911 => to_signed(26657, LUT_AMPL_WIDTH),
		9912 => to_signed(26659, LUT_AMPL_WIDTH),
		9913 => to_signed(26661, LUT_AMPL_WIDTH),
		9914 => to_signed(26663, LUT_AMPL_WIDTH),
		9915 => to_signed(26664, LUT_AMPL_WIDTH),
		9916 => to_signed(26666, LUT_AMPL_WIDTH),
		9917 => to_signed(26668, LUT_AMPL_WIDTH),
		9918 => to_signed(26670, LUT_AMPL_WIDTH),
		9919 => to_signed(26672, LUT_AMPL_WIDTH),
		9920 => to_signed(26674, LUT_AMPL_WIDTH),
		9921 => to_signed(26675, LUT_AMPL_WIDTH),
		9922 => to_signed(26677, LUT_AMPL_WIDTH),
		9923 => to_signed(26679, LUT_AMPL_WIDTH),
		9924 => to_signed(26681, LUT_AMPL_WIDTH),
		9925 => to_signed(26683, LUT_AMPL_WIDTH),
		9926 => to_signed(26684, LUT_AMPL_WIDTH),
		9927 => to_signed(26686, LUT_AMPL_WIDTH),
		9928 => to_signed(26688, LUT_AMPL_WIDTH),
		9929 => to_signed(26690, LUT_AMPL_WIDTH),
		9930 => to_signed(26692, LUT_AMPL_WIDTH),
		9931 => to_signed(26694, LUT_AMPL_WIDTH),
		9932 => to_signed(26695, LUT_AMPL_WIDTH),
		9933 => to_signed(26697, LUT_AMPL_WIDTH),
		9934 => to_signed(26699, LUT_AMPL_WIDTH),
		9935 => to_signed(26701, LUT_AMPL_WIDTH),
		9936 => to_signed(26703, LUT_AMPL_WIDTH),
		9937 => to_signed(26705, LUT_AMPL_WIDTH),
		9938 => to_signed(26706, LUT_AMPL_WIDTH),
		9939 => to_signed(26708, LUT_AMPL_WIDTH),
		9940 => to_signed(26710, LUT_AMPL_WIDTH),
		9941 => to_signed(26712, LUT_AMPL_WIDTH),
		9942 => to_signed(26714, LUT_AMPL_WIDTH),
		9943 => to_signed(26715, LUT_AMPL_WIDTH),
		9944 => to_signed(26717, LUT_AMPL_WIDTH),
		9945 => to_signed(26719, LUT_AMPL_WIDTH),
		9946 => to_signed(26721, LUT_AMPL_WIDTH),
		9947 => to_signed(26723, LUT_AMPL_WIDTH),
		9948 => to_signed(26725, LUT_AMPL_WIDTH),
		9949 => to_signed(26726, LUT_AMPL_WIDTH),
		9950 => to_signed(26728, LUT_AMPL_WIDTH),
		9951 => to_signed(26730, LUT_AMPL_WIDTH),
		9952 => to_signed(26732, LUT_AMPL_WIDTH),
		9953 => to_signed(26734, LUT_AMPL_WIDTH),
		9954 => to_signed(26735, LUT_AMPL_WIDTH),
		9955 => to_signed(26737, LUT_AMPL_WIDTH),
		9956 => to_signed(26739, LUT_AMPL_WIDTH),
		9957 => to_signed(26741, LUT_AMPL_WIDTH),
		9958 => to_signed(26743, LUT_AMPL_WIDTH),
		9959 => to_signed(26745, LUT_AMPL_WIDTH),
		9960 => to_signed(26746, LUT_AMPL_WIDTH),
		9961 => to_signed(26748, LUT_AMPL_WIDTH),
		9962 => to_signed(26750, LUT_AMPL_WIDTH),
		9963 => to_signed(26752, LUT_AMPL_WIDTH),
		9964 => to_signed(26754, LUT_AMPL_WIDTH),
		9965 => to_signed(26755, LUT_AMPL_WIDTH),
		9966 => to_signed(26757, LUT_AMPL_WIDTH),
		9967 => to_signed(26759, LUT_AMPL_WIDTH),
		9968 => to_signed(26761, LUT_AMPL_WIDTH),
		9969 => to_signed(26763, LUT_AMPL_WIDTH),
		9970 => to_signed(26764, LUT_AMPL_WIDTH),
		9971 => to_signed(26766, LUT_AMPL_WIDTH),
		9972 => to_signed(26768, LUT_AMPL_WIDTH),
		9973 => to_signed(26770, LUT_AMPL_WIDTH),
		9974 => to_signed(26772, LUT_AMPL_WIDTH),
		9975 => to_signed(26774, LUT_AMPL_WIDTH),
		9976 => to_signed(26775, LUT_AMPL_WIDTH),
		9977 => to_signed(26777, LUT_AMPL_WIDTH),
		9978 => to_signed(26779, LUT_AMPL_WIDTH),
		9979 => to_signed(26781, LUT_AMPL_WIDTH),
		9980 => to_signed(26783, LUT_AMPL_WIDTH),
		9981 => to_signed(26784, LUT_AMPL_WIDTH),
		9982 => to_signed(26786, LUT_AMPL_WIDTH),
		9983 => to_signed(26788, LUT_AMPL_WIDTH),
		9984 => to_signed(26790, LUT_AMPL_WIDTH),
		9985 => to_signed(26792, LUT_AMPL_WIDTH),
		9986 => to_signed(26793, LUT_AMPL_WIDTH),
		9987 => to_signed(26795, LUT_AMPL_WIDTH),
		9988 => to_signed(26797, LUT_AMPL_WIDTH),
		9989 => to_signed(26799, LUT_AMPL_WIDTH),
		9990 => to_signed(26801, LUT_AMPL_WIDTH),
		9991 => to_signed(26802, LUT_AMPL_WIDTH),
		9992 => to_signed(26804, LUT_AMPL_WIDTH),
		9993 => to_signed(26806, LUT_AMPL_WIDTH),
		9994 => to_signed(26808, LUT_AMPL_WIDTH),
		9995 => to_signed(26810, LUT_AMPL_WIDTH),
		9996 => to_signed(26811, LUT_AMPL_WIDTH),
		9997 => to_signed(26813, LUT_AMPL_WIDTH),
		9998 => to_signed(26815, LUT_AMPL_WIDTH),
		9999 => to_signed(26817, LUT_AMPL_WIDTH),
		10000 => to_signed(26819, LUT_AMPL_WIDTH),
		10001 => to_signed(26821, LUT_AMPL_WIDTH),
		10002 => to_signed(26822, LUT_AMPL_WIDTH),
		10003 => to_signed(26824, LUT_AMPL_WIDTH),
		10004 => to_signed(26826, LUT_AMPL_WIDTH),
		10005 => to_signed(26828, LUT_AMPL_WIDTH),
		10006 => to_signed(26830, LUT_AMPL_WIDTH),
		10007 => to_signed(26831, LUT_AMPL_WIDTH),
		10008 => to_signed(26833, LUT_AMPL_WIDTH),
		10009 => to_signed(26835, LUT_AMPL_WIDTH),
		10010 => to_signed(26837, LUT_AMPL_WIDTH),
		10011 => to_signed(26839, LUT_AMPL_WIDTH),
		10012 => to_signed(26840, LUT_AMPL_WIDTH),
		10013 => to_signed(26842, LUT_AMPL_WIDTH),
		10014 => to_signed(26844, LUT_AMPL_WIDTH),
		10015 => to_signed(26846, LUT_AMPL_WIDTH),
		10016 => to_signed(26848, LUT_AMPL_WIDTH),
		10017 => to_signed(26849, LUT_AMPL_WIDTH),
		10018 => to_signed(26851, LUT_AMPL_WIDTH),
		10019 => to_signed(26853, LUT_AMPL_WIDTH),
		10020 => to_signed(26855, LUT_AMPL_WIDTH),
		10021 => to_signed(26857, LUT_AMPL_WIDTH),
		10022 => to_signed(26858, LUT_AMPL_WIDTH),
		10023 => to_signed(26860, LUT_AMPL_WIDTH),
		10024 => to_signed(26862, LUT_AMPL_WIDTH),
		10025 => to_signed(26864, LUT_AMPL_WIDTH),
		10026 => to_signed(26866, LUT_AMPL_WIDTH),
		10027 => to_signed(26867, LUT_AMPL_WIDTH),
		10028 => to_signed(26869, LUT_AMPL_WIDTH),
		10029 => to_signed(26871, LUT_AMPL_WIDTH),
		10030 => to_signed(26873, LUT_AMPL_WIDTH),
		10031 => to_signed(26875, LUT_AMPL_WIDTH),
		10032 => to_signed(26876, LUT_AMPL_WIDTH),
		10033 => to_signed(26878, LUT_AMPL_WIDTH),
		10034 => to_signed(26880, LUT_AMPL_WIDTH),
		10035 => to_signed(26882, LUT_AMPL_WIDTH),
		10036 => to_signed(26884, LUT_AMPL_WIDTH),
		10037 => to_signed(26885, LUT_AMPL_WIDTH),
		10038 => to_signed(26887, LUT_AMPL_WIDTH),
		10039 => to_signed(26889, LUT_AMPL_WIDTH),
		10040 => to_signed(26891, LUT_AMPL_WIDTH),
		10041 => to_signed(26893, LUT_AMPL_WIDTH),
		10042 => to_signed(26894, LUT_AMPL_WIDTH),
		10043 => to_signed(26896, LUT_AMPL_WIDTH),
		10044 => to_signed(26898, LUT_AMPL_WIDTH),
		10045 => to_signed(26900, LUT_AMPL_WIDTH),
		10046 => to_signed(26901, LUT_AMPL_WIDTH),
		10047 => to_signed(26903, LUT_AMPL_WIDTH),
		10048 => to_signed(26905, LUT_AMPL_WIDTH),
		10049 => to_signed(26907, LUT_AMPL_WIDTH),
		10050 => to_signed(26909, LUT_AMPL_WIDTH),
		10051 => to_signed(26910, LUT_AMPL_WIDTH),
		10052 => to_signed(26912, LUT_AMPL_WIDTH),
		10053 => to_signed(26914, LUT_AMPL_WIDTH),
		10054 => to_signed(26916, LUT_AMPL_WIDTH),
		10055 => to_signed(26918, LUT_AMPL_WIDTH),
		10056 => to_signed(26919, LUT_AMPL_WIDTH),
		10057 => to_signed(26921, LUT_AMPL_WIDTH),
		10058 => to_signed(26923, LUT_AMPL_WIDTH),
		10059 => to_signed(26925, LUT_AMPL_WIDTH),
		10060 => to_signed(26927, LUT_AMPL_WIDTH),
		10061 => to_signed(26928, LUT_AMPL_WIDTH),
		10062 => to_signed(26930, LUT_AMPL_WIDTH),
		10063 => to_signed(26932, LUT_AMPL_WIDTH),
		10064 => to_signed(26934, LUT_AMPL_WIDTH),
		10065 => to_signed(26936, LUT_AMPL_WIDTH),
		10066 => to_signed(26937, LUT_AMPL_WIDTH),
		10067 => to_signed(26939, LUT_AMPL_WIDTH),
		10068 => to_signed(26941, LUT_AMPL_WIDTH),
		10069 => to_signed(26943, LUT_AMPL_WIDTH),
		10070 => to_signed(26944, LUT_AMPL_WIDTH),
		10071 => to_signed(26946, LUT_AMPL_WIDTH),
		10072 => to_signed(26948, LUT_AMPL_WIDTH),
		10073 => to_signed(26950, LUT_AMPL_WIDTH),
		10074 => to_signed(26952, LUT_AMPL_WIDTH),
		10075 => to_signed(26953, LUT_AMPL_WIDTH),
		10076 => to_signed(26955, LUT_AMPL_WIDTH),
		10077 => to_signed(26957, LUT_AMPL_WIDTH),
		10078 => to_signed(26959, LUT_AMPL_WIDTH),
		10079 => to_signed(26961, LUT_AMPL_WIDTH),
		10080 => to_signed(26962, LUT_AMPL_WIDTH),
		10081 => to_signed(26964, LUT_AMPL_WIDTH),
		10082 => to_signed(26966, LUT_AMPL_WIDTH),
		10083 => to_signed(26968, LUT_AMPL_WIDTH),
		10084 => to_signed(26969, LUT_AMPL_WIDTH),
		10085 => to_signed(26971, LUT_AMPL_WIDTH),
		10086 => to_signed(26973, LUT_AMPL_WIDTH),
		10087 => to_signed(26975, LUT_AMPL_WIDTH),
		10088 => to_signed(26977, LUT_AMPL_WIDTH),
		10089 => to_signed(26978, LUT_AMPL_WIDTH),
		10090 => to_signed(26980, LUT_AMPL_WIDTH),
		10091 => to_signed(26982, LUT_AMPL_WIDTH),
		10092 => to_signed(26984, LUT_AMPL_WIDTH),
		10093 => to_signed(26986, LUT_AMPL_WIDTH),
		10094 => to_signed(26987, LUT_AMPL_WIDTH),
		10095 => to_signed(26989, LUT_AMPL_WIDTH),
		10096 => to_signed(26991, LUT_AMPL_WIDTH),
		10097 => to_signed(26993, LUT_AMPL_WIDTH),
		10098 => to_signed(26994, LUT_AMPL_WIDTH),
		10099 => to_signed(26996, LUT_AMPL_WIDTH),
		10100 => to_signed(26998, LUT_AMPL_WIDTH),
		10101 => to_signed(27000, LUT_AMPL_WIDTH),
		10102 => to_signed(27002, LUT_AMPL_WIDTH),
		10103 => to_signed(27003, LUT_AMPL_WIDTH),
		10104 => to_signed(27005, LUT_AMPL_WIDTH),
		10105 => to_signed(27007, LUT_AMPL_WIDTH),
		10106 => to_signed(27009, LUT_AMPL_WIDTH),
		10107 => to_signed(27010, LUT_AMPL_WIDTH),
		10108 => to_signed(27012, LUT_AMPL_WIDTH),
		10109 => to_signed(27014, LUT_AMPL_WIDTH),
		10110 => to_signed(27016, LUT_AMPL_WIDTH),
		10111 => to_signed(27018, LUT_AMPL_WIDTH),
		10112 => to_signed(27019, LUT_AMPL_WIDTH),
		10113 => to_signed(27021, LUT_AMPL_WIDTH),
		10114 => to_signed(27023, LUT_AMPL_WIDTH),
		10115 => to_signed(27025, LUT_AMPL_WIDTH),
		10116 => to_signed(27026, LUT_AMPL_WIDTH),
		10117 => to_signed(27028, LUT_AMPL_WIDTH),
		10118 => to_signed(27030, LUT_AMPL_WIDTH),
		10119 => to_signed(27032, LUT_AMPL_WIDTH),
		10120 => to_signed(27034, LUT_AMPL_WIDTH),
		10121 => to_signed(27035, LUT_AMPL_WIDTH),
		10122 => to_signed(27037, LUT_AMPL_WIDTH),
		10123 => to_signed(27039, LUT_AMPL_WIDTH),
		10124 => to_signed(27041, LUT_AMPL_WIDTH),
		10125 => to_signed(27042, LUT_AMPL_WIDTH),
		10126 => to_signed(27044, LUT_AMPL_WIDTH),
		10127 => to_signed(27046, LUT_AMPL_WIDTH),
		10128 => to_signed(27048, LUT_AMPL_WIDTH),
		10129 => to_signed(27049, LUT_AMPL_WIDTH),
		10130 => to_signed(27051, LUT_AMPL_WIDTH),
		10131 => to_signed(27053, LUT_AMPL_WIDTH),
		10132 => to_signed(27055, LUT_AMPL_WIDTH),
		10133 => to_signed(27057, LUT_AMPL_WIDTH),
		10134 => to_signed(27058, LUT_AMPL_WIDTH),
		10135 => to_signed(27060, LUT_AMPL_WIDTH),
		10136 => to_signed(27062, LUT_AMPL_WIDTH),
		10137 => to_signed(27064, LUT_AMPL_WIDTH),
		10138 => to_signed(27065, LUT_AMPL_WIDTH),
		10139 => to_signed(27067, LUT_AMPL_WIDTH),
		10140 => to_signed(27069, LUT_AMPL_WIDTH),
		10141 => to_signed(27071, LUT_AMPL_WIDTH),
		10142 => to_signed(27073, LUT_AMPL_WIDTH),
		10143 => to_signed(27074, LUT_AMPL_WIDTH),
		10144 => to_signed(27076, LUT_AMPL_WIDTH),
		10145 => to_signed(27078, LUT_AMPL_WIDTH),
		10146 => to_signed(27080, LUT_AMPL_WIDTH),
		10147 => to_signed(27081, LUT_AMPL_WIDTH),
		10148 => to_signed(27083, LUT_AMPL_WIDTH),
		10149 => to_signed(27085, LUT_AMPL_WIDTH),
		10150 => to_signed(27087, LUT_AMPL_WIDTH),
		10151 => to_signed(27088, LUT_AMPL_WIDTH),
		10152 => to_signed(27090, LUT_AMPL_WIDTH),
		10153 => to_signed(27092, LUT_AMPL_WIDTH),
		10154 => to_signed(27094, LUT_AMPL_WIDTH),
		10155 => to_signed(27096, LUT_AMPL_WIDTH),
		10156 => to_signed(27097, LUT_AMPL_WIDTH),
		10157 => to_signed(27099, LUT_AMPL_WIDTH),
		10158 => to_signed(27101, LUT_AMPL_WIDTH),
		10159 => to_signed(27103, LUT_AMPL_WIDTH),
		10160 => to_signed(27104, LUT_AMPL_WIDTH),
		10161 => to_signed(27106, LUT_AMPL_WIDTH),
		10162 => to_signed(27108, LUT_AMPL_WIDTH),
		10163 => to_signed(27110, LUT_AMPL_WIDTH),
		10164 => to_signed(27111, LUT_AMPL_WIDTH),
		10165 => to_signed(27113, LUT_AMPL_WIDTH),
		10166 => to_signed(27115, LUT_AMPL_WIDTH),
		10167 => to_signed(27117, LUT_AMPL_WIDTH),
		10168 => to_signed(27118, LUT_AMPL_WIDTH),
		10169 => to_signed(27120, LUT_AMPL_WIDTH),
		10170 => to_signed(27122, LUT_AMPL_WIDTH),
		10171 => to_signed(27124, LUT_AMPL_WIDTH),
		10172 => to_signed(27126, LUT_AMPL_WIDTH),
		10173 => to_signed(27127, LUT_AMPL_WIDTH),
		10174 => to_signed(27129, LUT_AMPL_WIDTH),
		10175 => to_signed(27131, LUT_AMPL_WIDTH),
		10176 => to_signed(27133, LUT_AMPL_WIDTH),
		10177 => to_signed(27134, LUT_AMPL_WIDTH),
		10178 => to_signed(27136, LUT_AMPL_WIDTH),
		10179 => to_signed(27138, LUT_AMPL_WIDTH),
		10180 => to_signed(27140, LUT_AMPL_WIDTH),
		10181 => to_signed(27141, LUT_AMPL_WIDTH),
		10182 => to_signed(27143, LUT_AMPL_WIDTH),
		10183 => to_signed(27145, LUT_AMPL_WIDTH),
		10184 => to_signed(27147, LUT_AMPL_WIDTH),
		10185 => to_signed(27148, LUT_AMPL_WIDTH),
		10186 => to_signed(27150, LUT_AMPL_WIDTH),
		10187 => to_signed(27152, LUT_AMPL_WIDTH),
		10188 => to_signed(27154, LUT_AMPL_WIDTH),
		10189 => to_signed(27155, LUT_AMPL_WIDTH),
		10190 => to_signed(27157, LUT_AMPL_WIDTH),
		10191 => to_signed(27159, LUT_AMPL_WIDTH),
		10192 => to_signed(27161, LUT_AMPL_WIDTH),
		10193 => to_signed(27162, LUT_AMPL_WIDTH),
		10194 => to_signed(27164, LUT_AMPL_WIDTH),
		10195 => to_signed(27166, LUT_AMPL_WIDTH),
		10196 => to_signed(27168, LUT_AMPL_WIDTH),
		10197 => to_signed(27169, LUT_AMPL_WIDTH),
		10198 => to_signed(27171, LUT_AMPL_WIDTH),
		10199 => to_signed(27173, LUT_AMPL_WIDTH),
		10200 => to_signed(27175, LUT_AMPL_WIDTH),
		10201 => to_signed(27177, LUT_AMPL_WIDTH),
		10202 => to_signed(27178, LUT_AMPL_WIDTH),
		10203 => to_signed(27180, LUT_AMPL_WIDTH),
		10204 => to_signed(27182, LUT_AMPL_WIDTH),
		10205 => to_signed(27184, LUT_AMPL_WIDTH),
		10206 => to_signed(27185, LUT_AMPL_WIDTH),
		10207 => to_signed(27187, LUT_AMPL_WIDTH),
		10208 => to_signed(27189, LUT_AMPL_WIDTH),
		10209 => to_signed(27191, LUT_AMPL_WIDTH),
		10210 => to_signed(27192, LUT_AMPL_WIDTH),
		10211 => to_signed(27194, LUT_AMPL_WIDTH),
		10212 => to_signed(27196, LUT_AMPL_WIDTH),
		10213 => to_signed(27198, LUT_AMPL_WIDTH),
		10214 => to_signed(27199, LUT_AMPL_WIDTH),
		10215 => to_signed(27201, LUT_AMPL_WIDTH),
		10216 => to_signed(27203, LUT_AMPL_WIDTH),
		10217 => to_signed(27205, LUT_AMPL_WIDTH),
		10218 => to_signed(27206, LUT_AMPL_WIDTH),
		10219 => to_signed(27208, LUT_AMPL_WIDTH),
		10220 => to_signed(27210, LUT_AMPL_WIDTH),
		10221 => to_signed(27212, LUT_AMPL_WIDTH),
		10222 => to_signed(27213, LUT_AMPL_WIDTH),
		10223 => to_signed(27215, LUT_AMPL_WIDTH),
		10224 => to_signed(27217, LUT_AMPL_WIDTH),
		10225 => to_signed(27219, LUT_AMPL_WIDTH),
		10226 => to_signed(27220, LUT_AMPL_WIDTH),
		10227 => to_signed(27222, LUT_AMPL_WIDTH),
		10228 => to_signed(27224, LUT_AMPL_WIDTH),
		10229 => to_signed(27226, LUT_AMPL_WIDTH),
		10230 => to_signed(27227, LUT_AMPL_WIDTH),
		10231 => to_signed(27229, LUT_AMPL_WIDTH),
		10232 => to_signed(27231, LUT_AMPL_WIDTH),
		10233 => to_signed(27233, LUT_AMPL_WIDTH),
		10234 => to_signed(27234, LUT_AMPL_WIDTH),
		10235 => to_signed(27236, LUT_AMPL_WIDTH),
		10236 => to_signed(27238, LUT_AMPL_WIDTH),
		10237 => to_signed(27240, LUT_AMPL_WIDTH),
		10238 => to_signed(27241, LUT_AMPL_WIDTH),
		10239 => to_signed(27243, LUT_AMPL_WIDTH),
		10240 => to_signed(27245, LUT_AMPL_WIDTH),
		10241 => to_signed(27247, LUT_AMPL_WIDTH),
		10242 => to_signed(27248, LUT_AMPL_WIDTH),
		10243 => to_signed(27250, LUT_AMPL_WIDTH),
		10244 => to_signed(27252, LUT_AMPL_WIDTH),
		10245 => to_signed(27253, LUT_AMPL_WIDTH),
		10246 => to_signed(27255, LUT_AMPL_WIDTH),
		10247 => to_signed(27257, LUT_AMPL_WIDTH),
		10248 => to_signed(27259, LUT_AMPL_WIDTH),
		10249 => to_signed(27260, LUT_AMPL_WIDTH),
		10250 => to_signed(27262, LUT_AMPL_WIDTH),
		10251 => to_signed(27264, LUT_AMPL_WIDTH),
		10252 => to_signed(27266, LUT_AMPL_WIDTH),
		10253 => to_signed(27267, LUT_AMPL_WIDTH),
		10254 => to_signed(27269, LUT_AMPL_WIDTH),
		10255 => to_signed(27271, LUT_AMPL_WIDTH),
		10256 => to_signed(27273, LUT_AMPL_WIDTH),
		10257 => to_signed(27274, LUT_AMPL_WIDTH),
		10258 => to_signed(27276, LUT_AMPL_WIDTH),
		10259 => to_signed(27278, LUT_AMPL_WIDTH),
		10260 => to_signed(27280, LUT_AMPL_WIDTH),
		10261 => to_signed(27281, LUT_AMPL_WIDTH),
		10262 => to_signed(27283, LUT_AMPL_WIDTH),
		10263 => to_signed(27285, LUT_AMPL_WIDTH),
		10264 => to_signed(27287, LUT_AMPL_WIDTH),
		10265 => to_signed(27288, LUT_AMPL_WIDTH),
		10266 => to_signed(27290, LUT_AMPL_WIDTH),
		10267 => to_signed(27292, LUT_AMPL_WIDTH),
		10268 => to_signed(27294, LUT_AMPL_WIDTH),
		10269 => to_signed(27295, LUT_AMPL_WIDTH),
		10270 => to_signed(27297, LUT_AMPL_WIDTH),
		10271 => to_signed(27299, LUT_AMPL_WIDTH),
		10272 => to_signed(27300, LUT_AMPL_WIDTH),
		10273 => to_signed(27302, LUT_AMPL_WIDTH),
		10274 => to_signed(27304, LUT_AMPL_WIDTH),
		10275 => to_signed(27306, LUT_AMPL_WIDTH),
		10276 => to_signed(27307, LUT_AMPL_WIDTH),
		10277 => to_signed(27309, LUT_AMPL_WIDTH),
		10278 => to_signed(27311, LUT_AMPL_WIDTH),
		10279 => to_signed(27313, LUT_AMPL_WIDTH),
		10280 => to_signed(27314, LUT_AMPL_WIDTH),
		10281 => to_signed(27316, LUT_AMPL_WIDTH),
		10282 => to_signed(27318, LUT_AMPL_WIDTH),
		10283 => to_signed(27320, LUT_AMPL_WIDTH),
		10284 => to_signed(27321, LUT_AMPL_WIDTH),
		10285 => to_signed(27323, LUT_AMPL_WIDTH),
		10286 => to_signed(27325, LUT_AMPL_WIDTH),
		10287 => to_signed(27327, LUT_AMPL_WIDTH),
		10288 => to_signed(27328, LUT_AMPL_WIDTH),
		10289 => to_signed(27330, LUT_AMPL_WIDTH),
		10290 => to_signed(27332, LUT_AMPL_WIDTH),
		10291 => to_signed(27333, LUT_AMPL_WIDTH),
		10292 => to_signed(27335, LUT_AMPL_WIDTH),
		10293 => to_signed(27337, LUT_AMPL_WIDTH),
		10294 => to_signed(27339, LUT_AMPL_WIDTH),
		10295 => to_signed(27340, LUT_AMPL_WIDTH),
		10296 => to_signed(27342, LUT_AMPL_WIDTH),
		10297 => to_signed(27344, LUT_AMPL_WIDTH),
		10298 => to_signed(27346, LUT_AMPL_WIDTH),
		10299 => to_signed(27347, LUT_AMPL_WIDTH),
		10300 => to_signed(27349, LUT_AMPL_WIDTH),
		10301 => to_signed(27351, LUT_AMPL_WIDTH),
		10302 => to_signed(27352, LUT_AMPL_WIDTH),
		10303 => to_signed(27354, LUT_AMPL_WIDTH),
		10304 => to_signed(27356, LUT_AMPL_WIDTH),
		10305 => to_signed(27358, LUT_AMPL_WIDTH),
		10306 => to_signed(27359, LUT_AMPL_WIDTH),
		10307 => to_signed(27361, LUT_AMPL_WIDTH),
		10308 => to_signed(27363, LUT_AMPL_WIDTH),
		10309 => to_signed(27365, LUT_AMPL_WIDTH),
		10310 => to_signed(27366, LUT_AMPL_WIDTH),
		10311 => to_signed(27368, LUT_AMPL_WIDTH),
		10312 => to_signed(27370, LUT_AMPL_WIDTH),
		10313 => to_signed(27372, LUT_AMPL_WIDTH),
		10314 => to_signed(27373, LUT_AMPL_WIDTH),
		10315 => to_signed(27375, LUT_AMPL_WIDTH),
		10316 => to_signed(27377, LUT_AMPL_WIDTH),
		10317 => to_signed(27378, LUT_AMPL_WIDTH),
		10318 => to_signed(27380, LUT_AMPL_WIDTH),
		10319 => to_signed(27382, LUT_AMPL_WIDTH),
		10320 => to_signed(27384, LUT_AMPL_WIDTH),
		10321 => to_signed(27385, LUT_AMPL_WIDTH),
		10322 => to_signed(27387, LUT_AMPL_WIDTH),
		10323 => to_signed(27389, LUT_AMPL_WIDTH),
		10324 => to_signed(27390, LUT_AMPL_WIDTH),
		10325 => to_signed(27392, LUT_AMPL_WIDTH),
		10326 => to_signed(27394, LUT_AMPL_WIDTH),
		10327 => to_signed(27396, LUT_AMPL_WIDTH),
		10328 => to_signed(27397, LUT_AMPL_WIDTH),
		10329 => to_signed(27399, LUT_AMPL_WIDTH),
		10330 => to_signed(27401, LUT_AMPL_WIDTH),
		10331 => to_signed(27403, LUT_AMPL_WIDTH),
		10332 => to_signed(27404, LUT_AMPL_WIDTH),
		10333 => to_signed(27406, LUT_AMPL_WIDTH),
		10334 => to_signed(27408, LUT_AMPL_WIDTH),
		10335 => to_signed(27409, LUT_AMPL_WIDTH),
		10336 => to_signed(27411, LUT_AMPL_WIDTH),
		10337 => to_signed(27413, LUT_AMPL_WIDTH),
		10338 => to_signed(27415, LUT_AMPL_WIDTH),
		10339 => to_signed(27416, LUT_AMPL_WIDTH),
		10340 => to_signed(27418, LUT_AMPL_WIDTH),
		10341 => to_signed(27420, LUT_AMPL_WIDTH),
		10342 => to_signed(27421, LUT_AMPL_WIDTH),
		10343 => to_signed(27423, LUT_AMPL_WIDTH),
		10344 => to_signed(27425, LUT_AMPL_WIDTH),
		10345 => to_signed(27427, LUT_AMPL_WIDTH),
		10346 => to_signed(27428, LUT_AMPL_WIDTH),
		10347 => to_signed(27430, LUT_AMPL_WIDTH),
		10348 => to_signed(27432, LUT_AMPL_WIDTH),
		10349 => to_signed(27434, LUT_AMPL_WIDTH),
		10350 => to_signed(27435, LUT_AMPL_WIDTH),
		10351 => to_signed(27437, LUT_AMPL_WIDTH),
		10352 => to_signed(27439, LUT_AMPL_WIDTH),
		10353 => to_signed(27440, LUT_AMPL_WIDTH),
		10354 => to_signed(27442, LUT_AMPL_WIDTH),
		10355 => to_signed(27444, LUT_AMPL_WIDTH),
		10356 => to_signed(27446, LUT_AMPL_WIDTH),
		10357 => to_signed(27447, LUT_AMPL_WIDTH),
		10358 => to_signed(27449, LUT_AMPL_WIDTH),
		10359 => to_signed(27451, LUT_AMPL_WIDTH),
		10360 => to_signed(27452, LUT_AMPL_WIDTH),
		10361 => to_signed(27454, LUT_AMPL_WIDTH),
		10362 => to_signed(27456, LUT_AMPL_WIDTH),
		10363 => to_signed(27458, LUT_AMPL_WIDTH),
		10364 => to_signed(27459, LUT_AMPL_WIDTH),
		10365 => to_signed(27461, LUT_AMPL_WIDTH),
		10366 => to_signed(27463, LUT_AMPL_WIDTH),
		10367 => to_signed(27464, LUT_AMPL_WIDTH),
		10368 => to_signed(27466, LUT_AMPL_WIDTH),
		10369 => to_signed(27468, LUT_AMPL_WIDTH),
		10370 => to_signed(27470, LUT_AMPL_WIDTH),
		10371 => to_signed(27471, LUT_AMPL_WIDTH),
		10372 => to_signed(27473, LUT_AMPL_WIDTH),
		10373 => to_signed(27475, LUT_AMPL_WIDTH),
		10374 => to_signed(27476, LUT_AMPL_WIDTH),
		10375 => to_signed(27478, LUT_AMPL_WIDTH),
		10376 => to_signed(27480, LUT_AMPL_WIDTH),
		10377 => to_signed(27482, LUT_AMPL_WIDTH),
		10378 => to_signed(27483, LUT_AMPL_WIDTH),
		10379 => to_signed(27485, LUT_AMPL_WIDTH),
		10380 => to_signed(27487, LUT_AMPL_WIDTH),
		10381 => to_signed(27488, LUT_AMPL_WIDTH),
		10382 => to_signed(27490, LUT_AMPL_WIDTH),
		10383 => to_signed(27492, LUT_AMPL_WIDTH),
		10384 => to_signed(27493, LUT_AMPL_WIDTH),
		10385 => to_signed(27495, LUT_AMPL_WIDTH),
		10386 => to_signed(27497, LUT_AMPL_WIDTH),
		10387 => to_signed(27499, LUT_AMPL_WIDTH),
		10388 => to_signed(27500, LUT_AMPL_WIDTH),
		10389 => to_signed(27502, LUT_AMPL_WIDTH),
		10390 => to_signed(27504, LUT_AMPL_WIDTH),
		10391 => to_signed(27505, LUT_AMPL_WIDTH),
		10392 => to_signed(27507, LUT_AMPL_WIDTH),
		10393 => to_signed(27509, LUT_AMPL_WIDTH),
		10394 => to_signed(27511, LUT_AMPL_WIDTH),
		10395 => to_signed(27512, LUT_AMPL_WIDTH),
		10396 => to_signed(27514, LUT_AMPL_WIDTH),
		10397 => to_signed(27516, LUT_AMPL_WIDTH),
		10398 => to_signed(27517, LUT_AMPL_WIDTH),
		10399 => to_signed(27519, LUT_AMPL_WIDTH),
		10400 => to_signed(27521, LUT_AMPL_WIDTH),
		10401 => to_signed(27523, LUT_AMPL_WIDTH),
		10402 => to_signed(27524, LUT_AMPL_WIDTH),
		10403 => to_signed(27526, LUT_AMPL_WIDTH),
		10404 => to_signed(27528, LUT_AMPL_WIDTH),
		10405 => to_signed(27529, LUT_AMPL_WIDTH),
		10406 => to_signed(27531, LUT_AMPL_WIDTH),
		10407 => to_signed(27533, LUT_AMPL_WIDTH),
		10408 => to_signed(27534, LUT_AMPL_WIDTH),
		10409 => to_signed(27536, LUT_AMPL_WIDTH),
		10410 => to_signed(27538, LUT_AMPL_WIDTH),
		10411 => to_signed(27540, LUT_AMPL_WIDTH),
		10412 => to_signed(27541, LUT_AMPL_WIDTH),
		10413 => to_signed(27543, LUT_AMPL_WIDTH),
		10414 => to_signed(27545, LUT_AMPL_WIDTH),
		10415 => to_signed(27546, LUT_AMPL_WIDTH),
		10416 => to_signed(27548, LUT_AMPL_WIDTH),
		10417 => to_signed(27550, LUT_AMPL_WIDTH),
		10418 => to_signed(27551, LUT_AMPL_WIDTH),
		10419 => to_signed(27553, LUT_AMPL_WIDTH),
		10420 => to_signed(27555, LUT_AMPL_WIDTH),
		10421 => to_signed(27557, LUT_AMPL_WIDTH),
		10422 => to_signed(27558, LUT_AMPL_WIDTH),
		10423 => to_signed(27560, LUT_AMPL_WIDTH),
		10424 => to_signed(27562, LUT_AMPL_WIDTH),
		10425 => to_signed(27563, LUT_AMPL_WIDTH),
		10426 => to_signed(27565, LUT_AMPL_WIDTH),
		10427 => to_signed(27567, LUT_AMPL_WIDTH),
		10428 => to_signed(27568, LUT_AMPL_WIDTH),
		10429 => to_signed(27570, LUT_AMPL_WIDTH),
		10430 => to_signed(27572, LUT_AMPL_WIDTH),
		10431 => to_signed(27574, LUT_AMPL_WIDTH),
		10432 => to_signed(27575, LUT_AMPL_WIDTH),
		10433 => to_signed(27577, LUT_AMPL_WIDTH),
		10434 => to_signed(27579, LUT_AMPL_WIDTH),
		10435 => to_signed(27580, LUT_AMPL_WIDTH),
		10436 => to_signed(27582, LUT_AMPL_WIDTH),
		10437 => to_signed(27584, LUT_AMPL_WIDTH),
		10438 => to_signed(27585, LUT_AMPL_WIDTH),
		10439 => to_signed(27587, LUT_AMPL_WIDTH),
		10440 => to_signed(27589, LUT_AMPL_WIDTH),
		10441 => to_signed(27590, LUT_AMPL_WIDTH),
		10442 => to_signed(27592, LUT_AMPL_WIDTH),
		10443 => to_signed(27594, LUT_AMPL_WIDTH),
		10444 => to_signed(27596, LUT_AMPL_WIDTH),
		10445 => to_signed(27597, LUT_AMPL_WIDTH),
		10446 => to_signed(27599, LUT_AMPL_WIDTH),
		10447 => to_signed(27601, LUT_AMPL_WIDTH),
		10448 => to_signed(27602, LUT_AMPL_WIDTH),
		10449 => to_signed(27604, LUT_AMPL_WIDTH),
		10450 => to_signed(27606, LUT_AMPL_WIDTH),
		10451 => to_signed(27607, LUT_AMPL_WIDTH),
		10452 => to_signed(27609, LUT_AMPL_WIDTH),
		10453 => to_signed(27611, LUT_AMPL_WIDTH),
		10454 => to_signed(27613, LUT_AMPL_WIDTH),
		10455 => to_signed(27614, LUT_AMPL_WIDTH),
		10456 => to_signed(27616, LUT_AMPL_WIDTH),
		10457 => to_signed(27618, LUT_AMPL_WIDTH),
		10458 => to_signed(27619, LUT_AMPL_WIDTH),
		10459 => to_signed(27621, LUT_AMPL_WIDTH),
		10460 => to_signed(27623, LUT_AMPL_WIDTH),
		10461 => to_signed(27624, LUT_AMPL_WIDTH),
		10462 => to_signed(27626, LUT_AMPL_WIDTH),
		10463 => to_signed(27628, LUT_AMPL_WIDTH),
		10464 => to_signed(27629, LUT_AMPL_WIDTH),
		10465 => to_signed(27631, LUT_AMPL_WIDTH),
		10466 => to_signed(27633, LUT_AMPL_WIDTH),
		10467 => to_signed(27634, LUT_AMPL_WIDTH),
		10468 => to_signed(27636, LUT_AMPL_WIDTH),
		10469 => to_signed(27638, LUT_AMPL_WIDTH),
		10470 => to_signed(27640, LUT_AMPL_WIDTH),
		10471 => to_signed(27641, LUT_AMPL_WIDTH),
		10472 => to_signed(27643, LUT_AMPL_WIDTH),
		10473 => to_signed(27645, LUT_AMPL_WIDTH),
		10474 => to_signed(27646, LUT_AMPL_WIDTH),
		10475 => to_signed(27648, LUT_AMPL_WIDTH),
		10476 => to_signed(27650, LUT_AMPL_WIDTH),
		10477 => to_signed(27651, LUT_AMPL_WIDTH),
		10478 => to_signed(27653, LUT_AMPL_WIDTH),
		10479 => to_signed(27655, LUT_AMPL_WIDTH),
		10480 => to_signed(27656, LUT_AMPL_WIDTH),
		10481 => to_signed(27658, LUT_AMPL_WIDTH),
		10482 => to_signed(27660, LUT_AMPL_WIDTH),
		10483 => to_signed(27661, LUT_AMPL_WIDTH),
		10484 => to_signed(27663, LUT_AMPL_WIDTH),
		10485 => to_signed(27665, LUT_AMPL_WIDTH),
		10486 => to_signed(27666, LUT_AMPL_WIDTH),
		10487 => to_signed(27668, LUT_AMPL_WIDTH),
		10488 => to_signed(27670, LUT_AMPL_WIDTH),
		10489 => to_signed(27672, LUT_AMPL_WIDTH),
		10490 => to_signed(27673, LUT_AMPL_WIDTH),
		10491 => to_signed(27675, LUT_AMPL_WIDTH),
		10492 => to_signed(27677, LUT_AMPL_WIDTH),
		10493 => to_signed(27678, LUT_AMPL_WIDTH),
		10494 => to_signed(27680, LUT_AMPL_WIDTH),
		10495 => to_signed(27682, LUT_AMPL_WIDTH),
		10496 => to_signed(27683, LUT_AMPL_WIDTH),
		10497 => to_signed(27685, LUT_AMPL_WIDTH),
		10498 => to_signed(27687, LUT_AMPL_WIDTH),
		10499 => to_signed(27688, LUT_AMPL_WIDTH),
		10500 => to_signed(27690, LUT_AMPL_WIDTH),
		10501 => to_signed(27692, LUT_AMPL_WIDTH),
		10502 => to_signed(27693, LUT_AMPL_WIDTH),
		10503 => to_signed(27695, LUT_AMPL_WIDTH),
		10504 => to_signed(27697, LUT_AMPL_WIDTH),
		10505 => to_signed(27698, LUT_AMPL_WIDTH),
		10506 => to_signed(27700, LUT_AMPL_WIDTH),
		10507 => to_signed(27702, LUT_AMPL_WIDTH),
		10508 => to_signed(27703, LUT_AMPL_WIDTH),
		10509 => to_signed(27705, LUT_AMPL_WIDTH),
		10510 => to_signed(27707, LUT_AMPL_WIDTH),
		10511 => to_signed(27708, LUT_AMPL_WIDTH),
		10512 => to_signed(27710, LUT_AMPL_WIDTH),
		10513 => to_signed(27712, LUT_AMPL_WIDTH),
		10514 => to_signed(27714, LUT_AMPL_WIDTH),
		10515 => to_signed(27715, LUT_AMPL_WIDTH),
		10516 => to_signed(27717, LUT_AMPL_WIDTH),
		10517 => to_signed(27719, LUT_AMPL_WIDTH),
		10518 => to_signed(27720, LUT_AMPL_WIDTH),
		10519 => to_signed(27722, LUT_AMPL_WIDTH),
		10520 => to_signed(27724, LUT_AMPL_WIDTH),
		10521 => to_signed(27725, LUT_AMPL_WIDTH),
		10522 => to_signed(27727, LUT_AMPL_WIDTH),
		10523 => to_signed(27729, LUT_AMPL_WIDTH),
		10524 => to_signed(27730, LUT_AMPL_WIDTH),
		10525 => to_signed(27732, LUT_AMPL_WIDTH),
		10526 => to_signed(27734, LUT_AMPL_WIDTH),
		10527 => to_signed(27735, LUT_AMPL_WIDTH),
		10528 => to_signed(27737, LUT_AMPL_WIDTH),
		10529 => to_signed(27739, LUT_AMPL_WIDTH),
		10530 => to_signed(27740, LUT_AMPL_WIDTH),
		10531 => to_signed(27742, LUT_AMPL_WIDTH),
		10532 => to_signed(27744, LUT_AMPL_WIDTH),
		10533 => to_signed(27745, LUT_AMPL_WIDTH),
		10534 => to_signed(27747, LUT_AMPL_WIDTH),
		10535 => to_signed(27749, LUT_AMPL_WIDTH),
		10536 => to_signed(27750, LUT_AMPL_WIDTH),
		10537 => to_signed(27752, LUT_AMPL_WIDTH),
		10538 => to_signed(27754, LUT_AMPL_WIDTH),
		10539 => to_signed(27755, LUT_AMPL_WIDTH),
		10540 => to_signed(27757, LUT_AMPL_WIDTH),
		10541 => to_signed(27759, LUT_AMPL_WIDTH),
		10542 => to_signed(27760, LUT_AMPL_WIDTH),
		10543 => to_signed(27762, LUT_AMPL_WIDTH),
		10544 => to_signed(27764, LUT_AMPL_WIDTH),
		10545 => to_signed(27765, LUT_AMPL_WIDTH),
		10546 => to_signed(27767, LUT_AMPL_WIDTH),
		10547 => to_signed(27769, LUT_AMPL_WIDTH),
		10548 => to_signed(27770, LUT_AMPL_WIDTH),
		10549 => to_signed(27772, LUT_AMPL_WIDTH),
		10550 => to_signed(27774, LUT_AMPL_WIDTH),
		10551 => to_signed(27775, LUT_AMPL_WIDTH),
		10552 => to_signed(27777, LUT_AMPL_WIDTH),
		10553 => to_signed(27779, LUT_AMPL_WIDTH),
		10554 => to_signed(27780, LUT_AMPL_WIDTH),
		10555 => to_signed(27782, LUT_AMPL_WIDTH),
		10556 => to_signed(27784, LUT_AMPL_WIDTH),
		10557 => to_signed(27785, LUT_AMPL_WIDTH),
		10558 => to_signed(27787, LUT_AMPL_WIDTH),
		10559 => to_signed(27789, LUT_AMPL_WIDTH),
		10560 => to_signed(27790, LUT_AMPL_WIDTH),
		10561 => to_signed(27792, LUT_AMPL_WIDTH),
		10562 => to_signed(27794, LUT_AMPL_WIDTH),
		10563 => to_signed(27795, LUT_AMPL_WIDTH),
		10564 => to_signed(27797, LUT_AMPL_WIDTH),
		10565 => to_signed(27799, LUT_AMPL_WIDTH),
		10566 => to_signed(27800, LUT_AMPL_WIDTH),
		10567 => to_signed(27802, LUT_AMPL_WIDTH),
		10568 => to_signed(27804, LUT_AMPL_WIDTH),
		10569 => to_signed(27805, LUT_AMPL_WIDTH),
		10570 => to_signed(27807, LUT_AMPL_WIDTH),
		10571 => to_signed(27809, LUT_AMPL_WIDTH),
		10572 => to_signed(27810, LUT_AMPL_WIDTH),
		10573 => to_signed(27812, LUT_AMPL_WIDTH),
		10574 => to_signed(27814, LUT_AMPL_WIDTH),
		10575 => to_signed(27815, LUT_AMPL_WIDTH),
		10576 => to_signed(27817, LUT_AMPL_WIDTH),
		10577 => to_signed(27819, LUT_AMPL_WIDTH),
		10578 => to_signed(27820, LUT_AMPL_WIDTH),
		10579 => to_signed(27822, LUT_AMPL_WIDTH),
		10580 => to_signed(27824, LUT_AMPL_WIDTH),
		10581 => to_signed(27825, LUT_AMPL_WIDTH),
		10582 => to_signed(27827, LUT_AMPL_WIDTH),
		10583 => to_signed(27829, LUT_AMPL_WIDTH),
		10584 => to_signed(27830, LUT_AMPL_WIDTH),
		10585 => to_signed(27832, LUT_AMPL_WIDTH),
		10586 => to_signed(27834, LUT_AMPL_WIDTH),
		10587 => to_signed(27835, LUT_AMPL_WIDTH),
		10588 => to_signed(27837, LUT_AMPL_WIDTH),
		10589 => to_signed(27839, LUT_AMPL_WIDTH),
		10590 => to_signed(27840, LUT_AMPL_WIDTH),
		10591 => to_signed(27842, LUT_AMPL_WIDTH),
		10592 => to_signed(27843, LUT_AMPL_WIDTH),
		10593 => to_signed(27845, LUT_AMPL_WIDTH),
		10594 => to_signed(27847, LUT_AMPL_WIDTH),
		10595 => to_signed(27848, LUT_AMPL_WIDTH),
		10596 => to_signed(27850, LUT_AMPL_WIDTH),
		10597 => to_signed(27852, LUT_AMPL_WIDTH),
		10598 => to_signed(27853, LUT_AMPL_WIDTH),
		10599 => to_signed(27855, LUT_AMPL_WIDTH),
		10600 => to_signed(27857, LUT_AMPL_WIDTH),
		10601 => to_signed(27858, LUT_AMPL_WIDTH),
		10602 => to_signed(27860, LUT_AMPL_WIDTH),
		10603 => to_signed(27862, LUT_AMPL_WIDTH),
		10604 => to_signed(27863, LUT_AMPL_WIDTH),
		10605 => to_signed(27865, LUT_AMPL_WIDTH),
		10606 => to_signed(27867, LUT_AMPL_WIDTH),
		10607 => to_signed(27868, LUT_AMPL_WIDTH),
		10608 => to_signed(27870, LUT_AMPL_WIDTH),
		10609 => to_signed(27872, LUT_AMPL_WIDTH),
		10610 => to_signed(27873, LUT_AMPL_WIDTH),
		10611 => to_signed(27875, LUT_AMPL_WIDTH),
		10612 => to_signed(27877, LUT_AMPL_WIDTH),
		10613 => to_signed(27878, LUT_AMPL_WIDTH),
		10614 => to_signed(27880, LUT_AMPL_WIDTH),
		10615 => to_signed(27882, LUT_AMPL_WIDTH),
		10616 => to_signed(27883, LUT_AMPL_WIDTH),
		10617 => to_signed(27885, LUT_AMPL_WIDTH),
		10618 => to_signed(27886, LUT_AMPL_WIDTH),
		10619 => to_signed(27888, LUT_AMPL_WIDTH),
		10620 => to_signed(27890, LUT_AMPL_WIDTH),
		10621 => to_signed(27891, LUT_AMPL_WIDTH),
		10622 => to_signed(27893, LUT_AMPL_WIDTH),
		10623 => to_signed(27895, LUT_AMPL_WIDTH),
		10624 => to_signed(27896, LUT_AMPL_WIDTH),
		10625 => to_signed(27898, LUT_AMPL_WIDTH),
		10626 => to_signed(27900, LUT_AMPL_WIDTH),
		10627 => to_signed(27901, LUT_AMPL_WIDTH),
		10628 => to_signed(27903, LUT_AMPL_WIDTH),
		10629 => to_signed(27905, LUT_AMPL_WIDTH),
		10630 => to_signed(27906, LUT_AMPL_WIDTH),
		10631 => to_signed(27908, LUT_AMPL_WIDTH),
		10632 => to_signed(27910, LUT_AMPL_WIDTH),
		10633 => to_signed(27911, LUT_AMPL_WIDTH),
		10634 => to_signed(27913, LUT_AMPL_WIDTH),
		10635 => to_signed(27914, LUT_AMPL_WIDTH),
		10636 => to_signed(27916, LUT_AMPL_WIDTH),
		10637 => to_signed(27918, LUT_AMPL_WIDTH),
		10638 => to_signed(27919, LUT_AMPL_WIDTH),
		10639 => to_signed(27921, LUT_AMPL_WIDTH),
		10640 => to_signed(27923, LUT_AMPL_WIDTH),
		10641 => to_signed(27924, LUT_AMPL_WIDTH),
		10642 => to_signed(27926, LUT_AMPL_WIDTH),
		10643 => to_signed(27928, LUT_AMPL_WIDTH),
		10644 => to_signed(27929, LUT_AMPL_WIDTH),
		10645 => to_signed(27931, LUT_AMPL_WIDTH),
		10646 => to_signed(27933, LUT_AMPL_WIDTH),
		10647 => to_signed(27934, LUT_AMPL_WIDTH),
		10648 => to_signed(27936, LUT_AMPL_WIDTH),
		10649 => to_signed(27937, LUT_AMPL_WIDTH),
		10650 => to_signed(27939, LUT_AMPL_WIDTH),
		10651 => to_signed(27941, LUT_AMPL_WIDTH),
		10652 => to_signed(27942, LUT_AMPL_WIDTH),
		10653 => to_signed(27944, LUT_AMPL_WIDTH),
		10654 => to_signed(27946, LUT_AMPL_WIDTH),
		10655 => to_signed(27947, LUT_AMPL_WIDTH),
		10656 => to_signed(27949, LUT_AMPL_WIDTH),
		10657 => to_signed(27951, LUT_AMPL_WIDTH),
		10658 => to_signed(27952, LUT_AMPL_WIDTH),
		10659 => to_signed(27954, LUT_AMPL_WIDTH),
		10660 => to_signed(27956, LUT_AMPL_WIDTH),
		10661 => to_signed(27957, LUT_AMPL_WIDTH),
		10662 => to_signed(27959, LUT_AMPL_WIDTH),
		10663 => to_signed(27960, LUT_AMPL_WIDTH),
		10664 => to_signed(27962, LUT_AMPL_WIDTH),
		10665 => to_signed(27964, LUT_AMPL_WIDTH),
		10666 => to_signed(27965, LUT_AMPL_WIDTH),
		10667 => to_signed(27967, LUT_AMPL_WIDTH),
		10668 => to_signed(27969, LUT_AMPL_WIDTH),
		10669 => to_signed(27970, LUT_AMPL_WIDTH),
		10670 => to_signed(27972, LUT_AMPL_WIDTH),
		10671 => to_signed(27974, LUT_AMPL_WIDTH),
		10672 => to_signed(27975, LUT_AMPL_WIDTH),
		10673 => to_signed(27977, LUT_AMPL_WIDTH),
		10674 => to_signed(27978, LUT_AMPL_WIDTH),
		10675 => to_signed(27980, LUT_AMPL_WIDTH),
		10676 => to_signed(27982, LUT_AMPL_WIDTH),
		10677 => to_signed(27983, LUT_AMPL_WIDTH),
		10678 => to_signed(27985, LUT_AMPL_WIDTH),
		10679 => to_signed(27987, LUT_AMPL_WIDTH),
		10680 => to_signed(27988, LUT_AMPL_WIDTH),
		10681 => to_signed(27990, LUT_AMPL_WIDTH),
		10682 => to_signed(27992, LUT_AMPL_WIDTH),
		10683 => to_signed(27993, LUT_AMPL_WIDTH),
		10684 => to_signed(27995, LUT_AMPL_WIDTH),
		10685 => to_signed(27996, LUT_AMPL_WIDTH),
		10686 => to_signed(27998, LUT_AMPL_WIDTH),
		10687 => to_signed(28000, LUT_AMPL_WIDTH),
		10688 => to_signed(28001, LUT_AMPL_WIDTH),
		10689 => to_signed(28003, LUT_AMPL_WIDTH),
		10690 => to_signed(28005, LUT_AMPL_WIDTH),
		10691 => to_signed(28006, LUT_AMPL_WIDTH),
		10692 => to_signed(28008, LUT_AMPL_WIDTH),
		10693 => to_signed(28009, LUT_AMPL_WIDTH),
		10694 => to_signed(28011, LUT_AMPL_WIDTH),
		10695 => to_signed(28013, LUT_AMPL_WIDTH),
		10696 => to_signed(28014, LUT_AMPL_WIDTH),
		10697 => to_signed(28016, LUT_AMPL_WIDTH),
		10698 => to_signed(28018, LUT_AMPL_WIDTH),
		10699 => to_signed(28019, LUT_AMPL_WIDTH),
		10700 => to_signed(28021, LUT_AMPL_WIDTH),
		10701 => to_signed(28022, LUT_AMPL_WIDTH),
		10702 => to_signed(28024, LUT_AMPL_WIDTH),
		10703 => to_signed(28026, LUT_AMPL_WIDTH),
		10704 => to_signed(28027, LUT_AMPL_WIDTH),
		10705 => to_signed(28029, LUT_AMPL_WIDTH),
		10706 => to_signed(28031, LUT_AMPL_WIDTH),
		10707 => to_signed(28032, LUT_AMPL_WIDTH),
		10708 => to_signed(28034, LUT_AMPL_WIDTH),
		10709 => to_signed(28036, LUT_AMPL_WIDTH),
		10710 => to_signed(28037, LUT_AMPL_WIDTH),
		10711 => to_signed(28039, LUT_AMPL_WIDTH),
		10712 => to_signed(28040, LUT_AMPL_WIDTH),
		10713 => to_signed(28042, LUT_AMPL_WIDTH),
		10714 => to_signed(28044, LUT_AMPL_WIDTH),
		10715 => to_signed(28045, LUT_AMPL_WIDTH),
		10716 => to_signed(28047, LUT_AMPL_WIDTH),
		10717 => to_signed(28049, LUT_AMPL_WIDTH),
		10718 => to_signed(28050, LUT_AMPL_WIDTH),
		10719 => to_signed(28052, LUT_AMPL_WIDTH),
		10720 => to_signed(28053, LUT_AMPL_WIDTH),
		10721 => to_signed(28055, LUT_AMPL_WIDTH),
		10722 => to_signed(28057, LUT_AMPL_WIDTH),
		10723 => to_signed(28058, LUT_AMPL_WIDTH),
		10724 => to_signed(28060, LUT_AMPL_WIDTH),
		10725 => to_signed(28061, LUT_AMPL_WIDTH),
		10726 => to_signed(28063, LUT_AMPL_WIDTH),
		10727 => to_signed(28065, LUT_AMPL_WIDTH),
		10728 => to_signed(28066, LUT_AMPL_WIDTH),
		10729 => to_signed(28068, LUT_AMPL_WIDTH),
		10730 => to_signed(28070, LUT_AMPL_WIDTH),
		10731 => to_signed(28071, LUT_AMPL_WIDTH),
		10732 => to_signed(28073, LUT_AMPL_WIDTH),
		10733 => to_signed(28074, LUT_AMPL_WIDTH),
		10734 => to_signed(28076, LUT_AMPL_WIDTH),
		10735 => to_signed(28078, LUT_AMPL_WIDTH),
		10736 => to_signed(28079, LUT_AMPL_WIDTH),
		10737 => to_signed(28081, LUT_AMPL_WIDTH),
		10738 => to_signed(28083, LUT_AMPL_WIDTH),
		10739 => to_signed(28084, LUT_AMPL_WIDTH),
		10740 => to_signed(28086, LUT_AMPL_WIDTH),
		10741 => to_signed(28087, LUT_AMPL_WIDTH),
		10742 => to_signed(28089, LUT_AMPL_WIDTH),
		10743 => to_signed(28091, LUT_AMPL_WIDTH),
		10744 => to_signed(28092, LUT_AMPL_WIDTH),
		10745 => to_signed(28094, LUT_AMPL_WIDTH),
		10746 => to_signed(28095, LUT_AMPL_WIDTH),
		10747 => to_signed(28097, LUT_AMPL_WIDTH),
		10748 => to_signed(28099, LUT_AMPL_WIDTH),
		10749 => to_signed(28100, LUT_AMPL_WIDTH),
		10750 => to_signed(28102, LUT_AMPL_WIDTH),
		10751 => to_signed(28104, LUT_AMPL_WIDTH),
		10752 => to_signed(28105, LUT_AMPL_WIDTH),
		10753 => to_signed(28107, LUT_AMPL_WIDTH),
		10754 => to_signed(28108, LUT_AMPL_WIDTH),
		10755 => to_signed(28110, LUT_AMPL_WIDTH),
		10756 => to_signed(28112, LUT_AMPL_WIDTH),
		10757 => to_signed(28113, LUT_AMPL_WIDTH),
		10758 => to_signed(28115, LUT_AMPL_WIDTH),
		10759 => to_signed(28116, LUT_AMPL_WIDTH),
		10760 => to_signed(28118, LUT_AMPL_WIDTH),
		10761 => to_signed(28120, LUT_AMPL_WIDTH),
		10762 => to_signed(28121, LUT_AMPL_WIDTH),
		10763 => to_signed(28123, LUT_AMPL_WIDTH),
		10764 => to_signed(28125, LUT_AMPL_WIDTH),
		10765 => to_signed(28126, LUT_AMPL_WIDTH),
		10766 => to_signed(28128, LUT_AMPL_WIDTH),
		10767 => to_signed(28129, LUT_AMPL_WIDTH),
		10768 => to_signed(28131, LUT_AMPL_WIDTH),
		10769 => to_signed(28133, LUT_AMPL_WIDTH),
		10770 => to_signed(28134, LUT_AMPL_WIDTH),
		10771 => to_signed(28136, LUT_AMPL_WIDTH),
		10772 => to_signed(28137, LUT_AMPL_WIDTH),
		10773 => to_signed(28139, LUT_AMPL_WIDTH),
		10774 => to_signed(28141, LUT_AMPL_WIDTH),
		10775 => to_signed(28142, LUT_AMPL_WIDTH),
		10776 => to_signed(28144, LUT_AMPL_WIDTH),
		10777 => to_signed(28145, LUT_AMPL_WIDTH),
		10778 => to_signed(28147, LUT_AMPL_WIDTH),
		10779 => to_signed(28149, LUT_AMPL_WIDTH),
		10780 => to_signed(28150, LUT_AMPL_WIDTH),
		10781 => to_signed(28152, LUT_AMPL_WIDTH),
		10782 => to_signed(28154, LUT_AMPL_WIDTH),
		10783 => to_signed(28155, LUT_AMPL_WIDTH),
		10784 => to_signed(28157, LUT_AMPL_WIDTH),
		10785 => to_signed(28158, LUT_AMPL_WIDTH),
		10786 => to_signed(28160, LUT_AMPL_WIDTH),
		10787 => to_signed(28162, LUT_AMPL_WIDTH),
		10788 => to_signed(28163, LUT_AMPL_WIDTH),
		10789 => to_signed(28165, LUT_AMPL_WIDTH),
		10790 => to_signed(28166, LUT_AMPL_WIDTH),
		10791 => to_signed(28168, LUT_AMPL_WIDTH),
		10792 => to_signed(28170, LUT_AMPL_WIDTH),
		10793 => to_signed(28171, LUT_AMPL_WIDTH),
		10794 => to_signed(28173, LUT_AMPL_WIDTH),
		10795 => to_signed(28174, LUT_AMPL_WIDTH),
		10796 => to_signed(28176, LUT_AMPL_WIDTH),
		10797 => to_signed(28178, LUT_AMPL_WIDTH),
		10798 => to_signed(28179, LUT_AMPL_WIDTH),
		10799 => to_signed(28181, LUT_AMPL_WIDTH),
		10800 => to_signed(28182, LUT_AMPL_WIDTH),
		10801 => to_signed(28184, LUT_AMPL_WIDTH),
		10802 => to_signed(28186, LUT_AMPL_WIDTH),
		10803 => to_signed(28187, LUT_AMPL_WIDTH),
		10804 => to_signed(28189, LUT_AMPL_WIDTH),
		10805 => to_signed(28190, LUT_AMPL_WIDTH),
		10806 => to_signed(28192, LUT_AMPL_WIDTH),
		10807 => to_signed(28194, LUT_AMPL_WIDTH),
		10808 => to_signed(28195, LUT_AMPL_WIDTH),
		10809 => to_signed(28197, LUT_AMPL_WIDTH),
		10810 => to_signed(28198, LUT_AMPL_WIDTH),
		10811 => to_signed(28200, LUT_AMPL_WIDTH),
		10812 => to_signed(28202, LUT_AMPL_WIDTH),
		10813 => to_signed(28203, LUT_AMPL_WIDTH),
		10814 => to_signed(28205, LUT_AMPL_WIDTH),
		10815 => to_signed(28206, LUT_AMPL_WIDTH),
		10816 => to_signed(28208, LUT_AMPL_WIDTH),
		10817 => to_signed(28210, LUT_AMPL_WIDTH),
		10818 => to_signed(28211, LUT_AMPL_WIDTH),
		10819 => to_signed(28213, LUT_AMPL_WIDTH),
		10820 => to_signed(28214, LUT_AMPL_WIDTH),
		10821 => to_signed(28216, LUT_AMPL_WIDTH),
		10822 => to_signed(28218, LUT_AMPL_WIDTH),
		10823 => to_signed(28219, LUT_AMPL_WIDTH),
		10824 => to_signed(28221, LUT_AMPL_WIDTH),
		10825 => to_signed(28222, LUT_AMPL_WIDTH),
		10826 => to_signed(28224, LUT_AMPL_WIDTH),
		10827 => to_signed(28226, LUT_AMPL_WIDTH),
		10828 => to_signed(28227, LUT_AMPL_WIDTH),
		10829 => to_signed(28229, LUT_AMPL_WIDTH),
		10830 => to_signed(28230, LUT_AMPL_WIDTH),
		10831 => to_signed(28232, LUT_AMPL_WIDTH),
		10832 => to_signed(28234, LUT_AMPL_WIDTH),
		10833 => to_signed(28235, LUT_AMPL_WIDTH),
		10834 => to_signed(28237, LUT_AMPL_WIDTH),
		10835 => to_signed(28238, LUT_AMPL_WIDTH),
		10836 => to_signed(28240, LUT_AMPL_WIDTH),
		10837 => to_signed(28242, LUT_AMPL_WIDTH),
		10838 => to_signed(28243, LUT_AMPL_WIDTH),
		10839 => to_signed(28245, LUT_AMPL_WIDTH),
		10840 => to_signed(28246, LUT_AMPL_WIDTH),
		10841 => to_signed(28248, LUT_AMPL_WIDTH),
		10842 => to_signed(28249, LUT_AMPL_WIDTH),
		10843 => to_signed(28251, LUT_AMPL_WIDTH),
		10844 => to_signed(28253, LUT_AMPL_WIDTH),
		10845 => to_signed(28254, LUT_AMPL_WIDTH),
		10846 => to_signed(28256, LUT_AMPL_WIDTH),
		10847 => to_signed(28257, LUT_AMPL_WIDTH),
		10848 => to_signed(28259, LUT_AMPL_WIDTH),
		10849 => to_signed(28261, LUT_AMPL_WIDTH),
		10850 => to_signed(28262, LUT_AMPL_WIDTH),
		10851 => to_signed(28264, LUT_AMPL_WIDTH),
		10852 => to_signed(28265, LUT_AMPL_WIDTH),
		10853 => to_signed(28267, LUT_AMPL_WIDTH),
		10854 => to_signed(28269, LUT_AMPL_WIDTH),
		10855 => to_signed(28270, LUT_AMPL_WIDTH),
		10856 => to_signed(28272, LUT_AMPL_WIDTH),
		10857 => to_signed(28273, LUT_AMPL_WIDTH),
		10858 => to_signed(28275, LUT_AMPL_WIDTH),
		10859 => to_signed(28277, LUT_AMPL_WIDTH),
		10860 => to_signed(28278, LUT_AMPL_WIDTH),
		10861 => to_signed(28280, LUT_AMPL_WIDTH),
		10862 => to_signed(28281, LUT_AMPL_WIDTH),
		10863 => to_signed(28283, LUT_AMPL_WIDTH),
		10864 => to_signed(28284, LUT_AMPL_WIDTH),
		10865 => to_signed(28286, LUT_AMPL_WIDTH),
		10866 => to_signed(28288, LUT_AMPL_WIDTH),
		10867 => to_signed(28289, LUT_AMPL_WIDTH),
		10868 => to_signed(28291, LUT_AMPL_WIDTH),
		10869 => to_signed(28292, LUT_AMPL_WIDTH),
		10870 => to_signed(28294, LUT_AMPL_WIDTH),
		10871 => to_signed(28296, LUT_AMPL_WIDTH),
		10872 => to_signed(28297, LUT_AMPL_WIDTH),
		10873 => to_signed(28299, LUT_AMPL_WIDTH),
		10874 => to_signed(28300, LUT_AMPL_WIDTH),
		10875 => to_signed(28302, LUT_AMPL_WIDTH),
		10876 => to_signed(28303, LUT_AMPL_WIDTH),
		10877 => to_signed(28305, LUT_AMPL_WIDTH),
		10878 => to_signed(28307, LUT_AMPL_WIDTH),
		10879 => to_signed(28308, LUT_AMPL_WIDTH),
		10880 => to_signed(28310, LUT_AMPL_WIDTH),
		10881 => to_signed(28311, LUT_AMPL_WIDTH),
		10882 => to_signed(28313, LUT_AMPL_WIDTH),
		10883 => to_signed(28315, LUT_AMPL_WIDTH),
		10884 => to_signed(28316, LUT_AMPL_WIDTH),
		10885 => to_signed(28318, LUT_AMPL_WIDTH),
		10886 => to_signed(28319, LUT_AMPL_WIDTH),
		10887 => to_signed(28321, LUT_AMPL_WIDTH),
		10888 => to_signed(28322, LUT_AMPL_WIDTH),
		10889 => to_signed(28324, LUT_AMPL_WIDTH),
		10890 => to_signed(28326, LUT_AMPL_WIDTH),
		10891 => to_signed(28327, LUT_AMPL_WIDTH),
		10892 => to_signed(28329, LUT_AMPL_WIDTH),
		10893 => to_signed(28330, LUT_AMPL_WIDTH),
		10894 => to_signed(28332, LUT_AMPL_WIDTH),
		10895 => to_signed(28333, LUT_AMPL_WIDTH),
		10896 => to_signed(28335, LUT_AMPL_WIDTH),
		10897 => to_signed(28337, LUT_AMPL_WIDTH),
		10898 => to_signed(28338, LUT_AMPL_WIDTH),
		10899 => to_signed(28340, LUT_AMPL_WIDTH),
		10900 => to_signed(28341, LUT_AMPL_WIDTH),
		10901 => to_signed(28343, LUT_AMPL_WIDTH),
		10902 => to_signed(28345, LUT_AMPL_WIDTH),
		10903 => to_signed(28346, LUT_AMPL_WIDTH),
		10904 => to_signed(28348, LUT_AMPL_WIDTH),
		10905 => to_signed(28349, LUT_AMPL_WIDTH),
		10906 => to_signed(28351, LUT_AMPL_WIDTH),
		10907 => to_signed(28352, LUT_AMPL_WIDTH),
		10908 => to_signed(28354, LUT_AMPL_WIDTH),
		10909 => to_signed(28356, LUT_AMPL_WIDTH),
		10910 => to_signed(28357, LUT_AMPL_WIDTH),
		10911 => to_signed(28359, LUT_AMPL_WIDTH),
		10912 => to_signed(28360, LUT_AMPL_WIDTH),
		10913 => to_signed(28362, LUT_AMPL_WIDTH),
		10914 => to_signed(28363, LUT_AMPL_WIDTH),
		10915 => to_signed(28365, LUT_AMPL_WIDTH),
		10916 => to_signed(28367, LUT_AMPL_WIDTH),
		10917 => to_signed(28368, LUT_AMPL_WIDTH),
		10918 => to_signed(28370, LUT_AMPL_WIDTH),
		10919 => to_signed(28371, LUT_AMPL_WIDTH),
		10920 => to_signed(28373, LUT_AMPL_WIDTH),
		10921 => to_signed(28374, LUT_AMPL_WIDTH),
		10922 => to_signed(28376, LUT_AMPL_WIDTH),
		10923 => to_signed(28378, LUT_AMPL_WIDTH),
		10924 => to_signed(28379, LUT_AMPL_WIDTH),
		10925 => to_signed(28381, LUT_AMPL_WIDTH),
		10926 => to_signed(28382, LUT_AMPL_WIDTH),
		10927 => to_signed(28384, LUT_AMPL_WIDTH),
		10928 => to_signed(28385, LUT_AMPL_WIDTH),
		10929 => to_signed(28387, LUT_AMPL_WIDTH),
		10930 => to_signed(28389, LUT_AMPL_WIDTH),
		10931 => to_signed(28390, LUT_AMPL_WIDTH),
		10932 => to_signed(28392, LUT_AMPL_WIDTH),
		10933 => to_signed(28393, LUT_AMPL_WIDTH),
		10934 => to_signed(28395, LUT_AMPL_WIDTH),
		10935 => to_signed(28396, LUT_AMPL_WIDTH),
		10936 => to_signed(28398, LUT_AMPL_WIDTH),
		10937 => to_signed(28400, LUT_AMPL_WIDTH),
		10938 => to_signed(28401, LUT_AMPL_WIDTH),
		10939 => to_signed(28403, LUT_AMPL_WIDTH),
		10940 => to_signed(28404, LUT_AMPL_WIDTH),
		10941 => to_signed(28406, LUT_AMPL_WIDTH),
		10942 => to_signed(28407, LUT_AMPL_WIDTH),
		10943 => to_signed(28409, LUT_AMPL_WIDTH),
		10944 => to_signed(28411, LUT_AMPL_WIDTH),
		10945 => to_signed(28412, LUT_AMPL_WIDTH),
		10946 => to_signed(28414, LUT_AMPL_WIDTH),
		10947 => to_signed(28415, LUT_AMPL_WIDTH),
		10948 => to_signed(28417, LUT_AMPL_WIDTH),
		10949 => to_signed(28418, LUT_AMPL_WIDTH),
		10950 => to_signed(28420, LUT_AMPL_WIDTH),
		10951 => to_signed(28421, LUT_AMPL_WIDTH),
		10952 => to_signed(28423, LUT_AMPL_WIDTH),
		10953 => to_signed(28425, LUT_AMPL_WIDTH),
		10954 => to_signed(28426, LUT_AMPL_WIDTH),
		10955 => to_signed(28428, LUT_AMPL_WIDTH),
		10956 => to_signed(28429, LUT_AMPL_WIDTH),
		10957 => to_signed(28431, LUT_AMPL_WIDTH),
		10958 => to_signed(28432, LUT_AMPL_WIDTH),
		10959 => to_signed(28434, LUT_AMPL_WIDTH),
		10960 => to_signed(28436, LUT_AMPL_WIDTH),
		10961 => to_signed(28437, LUT_AMPL_WIDTH),
		10962 => to_signed(28439, LUT_AMPL_WIDTH),
		10963 => to_signed(28440, LUT_AMPL_WIDTH),
		10964 => to_signed(28442, LUT_AMPL_WIDTH),
		10965 => to_signed(28443, LUT_AMPL_WIDTH),
		10966 => to_signed(28445, LUT_AMPL_WIDTH),
		10967 => to_signed(28446, LUT_AMPL_WIDTH),
		10968 => to_signed(28448, LUT_AMPL_WIDTH),
		10969 => to_signed(28450, LUT_AMPL_WIDTH),
		10970 => to_signed(28451, LUT_AMPL_WIDTH),
		10971 => to_signed(28453, LUT_AMPL_WIDTH),
		10972 => to_signed(28454, LUT_AMPL_WIDTH),
		10973 => to_signed(28456, LUT_AMPL_WIDTH),
		10974 => to_signed(28457, LUT_AMPL_WIDTH),
		10975 => to_signed(28459, LUT_AMPL_WIDTH),
		10976 => to_signed(28460, LUT_AMPL_WIDTH),
		10977 => to_signed(28462, LUT_AMPL_WIDTH),
		10978 => to_signed(28464, LUT_AMPL_WIDTH),
		10979 => to_signed(28465, LUT_AMPL_WIDTH),
		10980 => to_signed(28467, LUT_AMPL_WIDTH),
		10981 => to_signed(28468, LUT_AMPL_WIDTH),
		10982 => to_signed(28470, LUT_AMPL_WIDTH),
		10983 => to_signed(28471, LUT_AMPL_WIDTH),
		10984 => to_signed(28473, LUT_AMPL_WIDTH),
		10985 => to_signed(28474, LUT_AMPL_WIDTH),
		10986 => to_signed(28476, LUT_AMPL_WIDTH),
		10987 => to_signed(28478, LUT_AMPL_WIDTH),
		10988 => to_signed(28479, LUT_AMPL_WIDTH),
		10989 => to_signed(28481, LUT_AMPL_WIDTH),
		10990 => to_signed(28482, LUT_AMPL_WIDTH),
		10991 => to_signed(28484, LUT_AMPL_WIDTH),
		10992 => to_signed(28485, LUT_AMPL_WIDTH),
		10993 => to_signed(28487, LUT_AMPL_WIDTH),
		10994 => to_signed(28488, LUT_AMPL_WIDTH),
		10995 => to_signed(28490, LUT_AMPL_WIDTH),
		10996 => to_signed(28492, LUT_AMPL_WIDTH),
		10997 => to_signed(28493, LUT_AMPL_WIDTH),
		10998 => to_signed(28495, LUT_AMPL_WIDTH),
		10999 => to_signed(28496, LUT_AMPL_WIDTH),
		11000 => to_signed(28498, LUT_AMPL_WIDTH),
		11001 => to_signed(28499, LUT_AMPL_WIDTH),
		11002 => to_signed(28501, LUT_AMPL_WIDTH),
		11003 => to_signed(28502, LUT_AMPL_WIDTH),
		11004 => to_signed(28504, LUT_AMPL_WIDTH),
		11005 => to_signed(28505, LUT_AMPL_WIDTH),
		11006 => to_signed(28507, LUT_AMPL_WIDTH),
		11007 => to_signed(28509, LUT_AMPL_WIDTH),
		11008 => to_signed(28510, LUT_AMPL_WIDTH),
		11009 => to_signed(28512, LUT_AMPL_WIDTH),
		11010 => to_signed(28513, LUT_AMPL_WIDTH),
		11011 => to_signed(28515, LUT_AMPL_WIDTH),
		11012 => to_signed(28516, LUT_AMPL_WIDTH),
		11013 => to_signed(28518, LUT_AMPL_WIDTH),
		11014 => to_signed(28519, LUT_AMPL_WIDTH),
		11015 => to_signed(28521, LUT_AMPL_WIDTH),
		11016 => to_signed(28523, LUT_AMPL_WIDTH),
		11017 => to_signed(28524, LUT_AMPL_WIDTH),
		11018 => to_signed(28526, LUT_AMPL_WIDTH),
		11019 => to_signed(28527, LUT_AMPL_WIDTH),
		11020 => to_signed(28529, LUT_AMPL_WIDTH),
		11021 => to_signed(28530, LUT_AMPL_WIDTH),
		11022 => to_signed(28532, LUT_AMPL_WIDTH),
		11023 => to_signed(28533, LUT_AMPL_WIDTH),
		11024 => to_signed(28535, LUT_AMPL_WIDTH),
		11025 => to_signed(28536, LUT_AMPL_WIDTH),
		11026 => to_signed(28538, LUT_AMPL_WIDTH),
		11027 => to_signed(28540, LUT_AMPL_WIDTH),
		11028 => to_signed(28541, LUT_AMPL_WIDTH),
		11029 => to_signed(28543, LUT_AMPL_WIDTH),
		11030 => to_signed(28544, LUT_AMPL_WIDTH),
		11031 => to_signed(28546, LUT_AMPL_WIDTH),
		11032 => to_signed(28547, LUT_AMPL_WIDTH),
		11033 => to_signed(28549, LUT_AMPL_WIDTH),
		11034 => to_signed(28550, LUT_AMPL_WIDTH),
		11035 => to_signed(28552, LUT_AMPL_WIDTH),
		11036 => to_signed(28553, LUT_AMPL_WIDTH),
		11037 => to_signed(28555, LUT_AMPL_WIDTH),
		11038 => to_signed(28556, LUT_AMPL_WIDTH),
		11039 => to_signed(28558, LUT_AMPL_WIDTH),
		11040 => to_signed(28560, LUT_AMPL_WIDTH),
		11041 => to_signed(28561, LUT_AMPL_WIDTH),
		11042 => to_signed(28563, LUT_AMPL_WIDTH),
		11043 => to_signed(28564, LUT_AMPL_WIDTH),
		11044 => to_signed(28566, LUT_AMPL_WIDTH),
		11045 => to_signed(28567, LUT_AMPL_WIDTH),
		11046 => to_signed(28569, LUT_AMPL_WIDTH),
		11047 => to_signed(28570, LUT_AMPL_WIDTH),
		11048 => to_signed(28572, LUT_AMPL_WIDTH),
		11049 => to_signed(28573, LUT_AMPL_WIDTH),
		11050 => to_signed(28575, LUT_AMPL_WIDTH),
		11051 => to_signed(28576, LUT_AMPL_WIDTH),
		11052 => to_signed(28578, LUT_AMPL_WIDTH),
		11053 => to_signed(28580, LUT_AMPL_WIDTH),
		11054 => to_signed(28581, LUT_AMPL_WIDTH),
		11055 => to_signed(28583, LUT_AMPL_WIDTH),
		11056 => to_signed(28584, LUT_AMPL_WIDTH),
		11057 => to_signed(28586, LUT_AMPL_WIDTH),
		11058 => to_signed(28587, LUT_AMPL_WIDTH),
		11059 => to_signed(28589, LUT_AMPL_WIDTH),
		11060 => to_signed(28590, LUT_AMPL_WIDTH),
		11061 => to_signed(28592, LUT_AMPL_WIDTH),
		11062 => to_signed(28593, LUT_AMPL_WIDTH),
		11063 => to_signed(28595, LUT_AMPL_WIDTH),
		11064 => to_signed(28596, LUT_AMPL_WIDTH),
		11065 => to_signed(28598, LUT_AMPL_WIDTH),
		11066 => to_signed(28600, LUT_AMPL_WIDTH),
		11067 => to_signed(28601, LUT_AMPL_WIDTH),
		11068 => to_signed(28603, LUT_AMPL_WIDTH),
		11069 => to_signed(28604, LUT_AMPL_WIDTH),
		11070 => to_signed(28606, LUT_AMPL_WIDTH),
		11071 => to_signed(28607, LUT_AMPL_WIDTH),
		11072 => to_signed(28609, LUT_AMPL_WIDTH),
		11073 => to_signed(28610, LUT_AMPL_WIDTH),
		11074 => to_signed(28612, LUT_AMPL_WIDTH),
		11075 => to_signed(28613, LUT_AMPL_WIDTH),
		11076 => to_signed(28615, LUT_AMPL_WIDTH),
		11077 => to_signed(28616, LUT_AMPL_WIDTH),
		11078 => to_signed(28618, LUT_AMPL_WIDTH),
		11079 => to_signed(28619, LUT_AMPL_WIDTH),
		11080 => to_signed(28621, LUT_AMPL_WIDTH),
		11081 => to_signed(28622, LUT_AMPL_WIDTH),
		11082 => to_signed(28624, LUT_AMPL_WIDTH),
		11083 => to_signed(28626, LUT_AMPL_WIDTH),
		11084 => to_signed(28627, LUT_AMPL_WIDTH),
		11085 => to_signed(28629, LUT_AMPL_WIDTH),
		11086 => to_signed(28630, LUT_AMPL_WIDTH),
		11087 => to_signed(28632, LUT_AMPL_WIDTH),
		11088 => to_signed(28633, LUT_AMPL_WIDTH),
		11089 => to_signed(28635, LUT_AMPL_WIDTH),
		11090 => to_signed(28636, LUT_AMPL_WIDTH),
		11091 => to_signed(28638, LUT_AMPL_WIDTH),
		11092 => to_signed(28639, LUT_AMPL_WIDTH),
		11093 => to_signed(28641, LUT_AMPL_WIDTH),
		11094 => to_signed(28642, LUT_AMPL_WIDTH),
		11095 => to_signed(28644, LUT_AMPL_WIDTH),
		11096 => to_signed(28645, LUT_AMPL_WIDTH),
		11097 => to_signed(28647, LUT_AMPL_WIDTH),
		11098 => to_signed(28648, LUT_AMPL_WIDTH),
		11099 => to_signed(28650, LUT_AMPL_WIDTH),
		11100 => to_signed(28651, LUT_AMPL_WIDTH),
		11101 => to_signed(28653, LUT_AMPL_WIDTH),
		11102 => to_signed(28655, LUT_AMPL_WIDTH),
		11103 => to_signed(28656, LUT_AMPL_WIDTH),
		11104 => to_signed(28658, LUT_AMPL_WIDTH),
		11105 => to_signed(28659, LUT_AMPL_WIDTH),
		11106 => to_signed(28661, LUT_AMPL_WIDTH),
		11107 => to_signed(28662, LUT_AMPL_WIDTH),
		11108 => to_signed(28664, LUT_AMPL_WIDTH),
		11109 => to_signed(28665, LUT_AMPL_WIDTH),
		11110 => to_signed(28667, LUT_AMPL_WIDTH),
		11111 => to_signed(28668, LUT_AMPL_WIDTH),
		11112 => to_signed(28670, LUT_AMPL_WIDTH),
		11113 => to_signed(28671, LUT_AMPL_WIDTH),
		11114 => to_signed(28673, LUT_AMPL_WIDTH),
		11115 => to_signed(28674, LUT_AMPL_WIDTH),
		11116 => to_signed(28676, LUT_AMPL_WIDTH),
		11117 => to_signed(28677, LUT_AMPL_WIDTH),
		11118 => to_signed(28679, LUT_AMPL_WIDTH),
		11119 => to_signed(28680, LUT_AMPL_WIDTH),
		11120 => to_signed(28682, LUT_AMPL_WIDTH),
		11121 => to_signed(28683, LUT_AMPL_WIDTH),
		11122 => to_signed(28685, LUT_AMPL_WIDTH),
		11123 => to_signed(28686, LUT_AMPL_WIDTH),
		11124 => to_signed(28688, LUT_AMPL_WIDTH),
		11125 => to_signed(28690, LUT_AMPL_WIDTH),
		11126 => to_signed(28691, LUT_AMPL_WIDTH),
		11127 => to_signed(28693, LUT_AMPL_WIDTH),
		11128 => to_signed(28694, LUT_AMPL_WIDTH),
		11129 => to_signed(28696, LUT_AMPL_WIDTH),
		11130 => to_signed(28697, LUT_AMPL_WIDTH),
		11131 => to_signed(28699, LUT_AMPL_WIDTH),
		11132 => to_signed(28700, LUT_AMPL_WIDTH),
		11133 => to_signed(28702, LUT_AMPL_WIDTH),
		11134 => to_signed(28703, LUT_AMPL_WIDTH),
		11135 => to_signed(28705, LUT_AMPL_WIDTH),
		11136 => to_signed(28706, LUT_AMPL_WIDTH),
		11137 => to_signed(28708, LUT_AMPL_WIDTH),
		11138 => to_signed(28709, LUT_AMPL_WIDTH),
		11139 => to_signed(28711, LUT_AMPL_WIDTH),
		11140 => to_signed(28712, LUT_AMPL_WIDTH),
		11141 => to_signed(28714, LUT_AMPL_WIDTH),
		11142 => to_signed(28715, LUT_AMPL_WIDTH),
		11143 => to_signed(28717, LUT_AMPL_WIDTH),
		11144 => to_signed(28718, LUT_AMPL_WIDTH),
		11145 => to_signed(28720, LUT_AMPL_WIDTH),
		11146 => to_signed(28721, LUT_AMPL_WIDTH),
		11147 => to_signed(28723, LUT_AMPL_WIDTH),
		11148 => to_signed(28724, LUT_AMPL_WIDTH),
		11149 => to_signed(28726, LUT_AMPL_WIDTH),
		11150 => to_signed(28727, LUT_AMPL_WIDTH),
		11151 => to_signed(28729, LUT_AMPL_WIDTH),
		11152 => to_signed(28730, LUT_AMPL_WIDTH),
		11153 => to_signed(28732, LUT_AMPL_WIDTH),
		11154 => to_signed(28733, LUT_AMPL_WIDTH),
		11155 => to_signed(28735, LUT_AMPL_WIDTH),
		11156 => to_signed(28736, LUT_AMPL_WIDTH),
		11157 => to_signed(28738, LUT_AMPL_WIDTH),
		11158 => to_signed(28739, LUT_AMPL_WIDTH),
		11159 => to_signed(28741, LUT_AMPL_WIDTH),
		11160 => to_signed(28742, LUT_AMPL_WIDTH),
		11161 => to_signed(28744, LUT_AMPL_WIDTH),
		11162 => to_signed(28745, LUT_AMPL_WIDTH),
		11163 => to_signed(28747, LUT_AMPL_WIDTH),
		11164 => to_signed(28748, LUT_AMPL_WIDTH),
		11165 => to_signed(28750, LUT_AMPL_WIDTH),
		11166 => to_signed(28752, LUT_AMPL_WIDTH),
		11167 => to_signed(28753, LUT_AMPL_WIDTH),
		11168 => to_signed(28755, LUT_AMPL_WIDTH),
		11169 => to_signed(28756, LUT_AMPL_WIDTH),
		11170 => to_signed(28758, LUT_AMPL_WIDTH),
		11171 => to_signed(28759, LUT_AMPL_WIDTH),
		11172 => to_signed(28761, LUT_AMPL_WIDTH),
		11173 => to_signed(28762, LUT_AMPL_WIDTH),
		11174 => to_signed(28764, LUT_AMPL_WIDTH),
		11175 => to_signed(28765, LUT_AMPL_WIDTH),
		11176 => to_signed(28767, LUT_AMPL_WIDTH),
		11177 => to_signed(28768, LUT_AMPL_WIDTH),
		11178 => to_signed(28770, LUT_AMPL_WIDTH),
		11179 => to_signed(28771, LUT_AMPL_WIDTH),
		11180 => to_signed(28773, LUT_AMPL_WIDTH),
		11181 => to_signed(28774, LUT_AMPL_WIDTH),
		11182 => to_signed(28776, LUT_AMPL_WIDTH),
		11183 => to_signed(28777, LUT_AMPL_WIDTH),
		11184 => to_signed(28779, LUT_AMPL_WIDTH),
		11185 => to_signed(28780, LUT_AMPL_WIDTH),
		11186 => to_signed(28782, LUT_AMPL_WIDTH),
		11187 => to_signed(28783, LUT_AMPL_WIDTH),
		11188 => to_signed(28785, LUT_AMPL_WIDTH),
		11189 => to_signed(28786, LUT_AMPL_WIDTH),
		11190 => to_signed(28788, LUT_AMPL_WIDTH),
		11191 => to_signed(28789, LUT_AMPL_WIDTH),
		11192 => to_signed(28791, LUT_AMPL_WIDTH),
		11193 => to_signed(28792, LUT_AMPL_WIDTH),
		11194 => to_signed(28794, LUT_AMPL_WIDTH),
		11195 => to_signed(28795, LUT_AMPL_WIDTH),
		11196 => to_signed(28797, LUT_AMPL_WIDTH),
		11197 => to_signed(28798, LUT_AMPL_WIDTH),
		11198 => to_signed(28800, LUT_AMPL_WIDTH),
		11199 => to_signed(28801, LUT_AMPL_WIDTH),
		11200 => to_signed(28803, LUT_AMPL_WIDTH),
		11201 => to_signed(28804, LUT_AMPL_WIDTH),
		11202 => to_signed(28806, LUT_AMPL_WIDTH),
		11203 => to_signed(28807, LUT_AMPL_WIDTH),
		11204 => to_signed(28809, LUT_AMPL_WIDTH),
		11205 => to_signed(28810, LUT_AMPL_WIDTH),
		11206 => to_signed(28812, LUT_AMPL_WIDTH),
		11207 => to_signed(28813, LUT_AMPL_WIDTH),
		11208 => to_signed(28815, LUT_AMPL_WIDTH),
		11209 => to_signed(28816, LUT_AMPL_WIDTH),
		11210 => to_signed(28818, LUT_AMPL_WIDTH),
		11211 => to_signed(28819, LUT_AMPL_WIDTH),
		11212 => to_signed(28821, LUT_AMPL_WIDTH),
		11213 => to_signed(28822, LUT_AMPL_WIDTH),
		11214 => to_signed(28824, LUT_AMPL_WIDTH),
		11215 => to_signed(28825, LUT_AMPL_WIDTH),
		11216 => to_signed(28827, LUT_AMPL_WIDTH),
		11217 => to_signed(28828, LUT_AMPL_WIDTH),
		11218 => to_signed(28830, LUT_AMPL_WIDTH),
		11219 => to_signed(28831, LUT_AMPL_WIDTH),
		11220 => to_signed(28832, LUT_AMPL_WIDTH),
		11221 => to_signed(28834, LUT_AMPL_WIDTH),
		11222 => to_signed(28835, LUT_AMPL_WIDTH),
		11223 => to_signed(28837, LUT_AMPL_WIDTH),
		11224 => to_signed(28838, LUT_AMPL_WIDTH),
		11225 => to_signed(28840, LUT_AMPL_WIDTH),
		11226 => to_signed(28841, LUT_AMPL_WIDTH),
		11227 => to_signed(28843, LUT_AMPL_WIDTH),
		11228 => to_signed(28844, LUT_AMPL_WIDTH),
		11229 => to_signed(28846, LUT_AMPL_WIDTH),
		11230 => to_signed(28847, LUT_AMPL_WIDTH),
		11231 => to_signed(28849, LUT_AMPL_WIDTH),
		11232 => to_signed(28850, LUT_AMPL_WIDTH),
		11233 => to_signed(28852, LUT_AMPL_WIDTH),
		11234 => to_signed(28853, LUT_AMPL_WIDTH),
		11235 => to_signed(28855, LUT_AMPL_WIDTH),
		11236 => to_signed(28856, LUT_AMPL_WIDTH),
		11237 => to_signed(28858, LUT_AMPL_WIDTH),
		11238 => to_signed(28859, LUT_AMPL_WIDTH),
		11239 => to_signed(28861, LUT_AMPL_WIDTH),
		11240 => to_signed(28862, LUT_AMPL_WIDTH),
		11241 => to_signed(28864, LUT_AMPL_WIDTH),
		11242 => to_signed(28865, LUT_AMPL_WIDTH),
		11243 => to_signed(28867, LUT_AMPL_WIDTH),
		11244 => to_signed(28868, LUT_AMPL_WIDTH),
		11245 => to_signed(28870, LUT_AMPL_WIDTH),
		11246 => to_signed(28871, LUT_AMPL_WIDTH),
		11247 => to_signed(28873, LUT_AMPL_WIDTH),
		11248 => to_signed(28874, LUT_AMPL_WIDTH),
		11249 => to_signed(28876, LUT_AMPL_WIDTH),
		11250 => to_signed(28877, LUT_AMPL_WIDTH),
		11251 => to_signed(28879, LUT_AMPL_WIDTH),
		11252 => to_signed(28880, LUT_AMPL_WIDTH),
		11253 => to_signed(28882, LUT_AMPL_WIDTH),
		11254 => to_signed(28883, LUT_AMPL_WIDTH),
		11255 => to_signed(28885, LUT_AMPL_WIDTH),
		11256 => to_signed(28886, LUT_AMPL_WIDTH),
		11257 => to_signed(28888, LUT_AMPL_WIDTH),
		11258 => to_signed(28889, LUT_AMPL_WIDTH),
		11259 => to_signed(28891, LUT_AMPL_WIDTH),
		11260 => to_signed(28892, LUT_AMPL_WIDTH),
		11261 => to_signed(28893, LUT_AMPL_WIDTH),
		11262 => to_signed(28895, LUT_AMPL_WIDTH),
		11263 => to_signed(28896, LUT_AMPL_WIDTH),
		11264 => to_signed(28898, LUT_AMPL_WIDTH),
		11265 => to_signed(28899, LUT_AMPL_WIDTH),
		11266 => to_signed(28901, LUT_AMPL_WIDTH),
		11267 => to_signed(28902, LUT_AMPL_WIDTH),
		11268 => to_signed(28904, LUT_AMPL_WIDTH),
		11269 => to_signed(28905, LUT_AMPL_WIDTH),
		11270 => to_signed(28907, LUT_AMPL_WIDTH),
		11271 => to_signed(28908, LUT_AMPL_WIDTH),
		11272 => to_signed(28910, LUT_AMPL_WIDTH),
		11273 => to_signed(28911, LUT_AMPL_WIDTH),
		11274 => to_signed(28913, LUT_AMPL_WIDTH),
		11275 => to_signed(28914, LUT_AMPL_WIDTH),
		11276 => to_signed(28916, LUT_AMPL_WIDTH),
		11277 => to_signed(28917, LUT_AMPL_WIDTH),
		11278 => to_signed(28919, LUT_AMPL_WIDTH),
		11279 => to_signed(28920, LUT_AMPL_WIDTH),
		11280 => to_signed(28922, LUT_AMPL_WIDTH),
		11281 => to_signed(28923, LUT_AMPL_WIDTH),
		11282 => to_signed(28925, LUT_AMPL_WIDTH),
		11283 => to_signed(28926, LUT_AMPL_WIDTH),
		11284 => to_signed(28927, LUT_AMPL_WIDTH),
		11285 => to_signed(28929, LUT_AMPL_WIDTH),
		11286 => to_signed(28930, LUT_AMPL_WIDTH),
		11287 => to_signed(28932, LUT_AMPL_WIDTH),
		11288 => to_signed(28933, LUT_AMPL_WIDTH),
		11289 => to_signed(28935, LUT_AMPL_WIDTH),
		11290 => to_signed(28936, LUT_AMPL_WIDTH),
		11291 => to_signed(28938, LUT_AMPL_WIDTH),
		11292 => to_signed(28939, LUT_AMPL_WIDTH),
		11293 => to_signed(28941, LUT_AMPL_WIDTH),
		11294 => to_signed(28942, LUT_AMPL_WIDTH),
		11295 => to_signed(28944, LUT_AMPL_WIDTH),
		11296 => to_signed(28945, LUT_AMPL_WIDTH),
		11297 => to_signed(28947, LUT_AMPL_WIDTH),
		11298 => to_signed(28948, LUT_AMPL_WIDTH),
		11299 => to_signed(28950, LUT_AMPL_WIDTH),
		11300 => to_signed(28951, LUT_AMPL_WIDTH),
		11301 => to_signed(28953, LUT_AMPL_WIDTH),
		11302 => to_signed(28954, LUT_AMPL_WIDTH),
		11303 => to_signed(28955, LUT_AMPL_WIDTH),
		11304 => to_signed(28957, LUT_AMPL_WIDTH),
		11305 => to_signed(28958, LUT_AMPL_WIDTH),
		11306 => to_signed(28960, LUT_AMPL_WIDTH),
		11307 => to_signed(28961, LUT_AMPL_WIDTH),
		11308 => to_signed(28963, LUT_AMPL_WIDTH),
		11309 => to_signed(28964, LUT_AMPL_WIDTH),
		11310 => to_signed(28966, LUT_AMPL_WIDTH),
		11311 => to_signed(28967, LUT_AMPL_WIDTH),
		11312 => to_signed(28969, LUT_AMPL_WIDTH),
		11313 => to_signed(28970, LUT_AMPL_WIDTH),
		11314 => to_signed(28972, LUT_AMPL_WIDTH),
		11315 => to_signed(28973, LUT_AMPL_WIDTH),
		11316 => to_signed(28975, LUT_AMPL_WIDTH),
		11317 => to_signed(28976, LUT_AMPL_WIDTH),
		11318 => to_signed(28977, LUT_AMPL_WIDTH),
		11319 => to_signed(28979, LUT_AMPL_WIDTH),
		11320 => to_signed(28980, LUT_AMPL_WIDTH),
		11321 => to_signed(28982, LUT_AMPL_WIDTH),
		11322 => to_signed(28983, LUT_AMPL_WIDTH),
		11323 => to_signed(28985, LUT_AMPL_WIDTH),
		11324 => to_signed(28986, LUT_AMPL_WIDTH),
		11325 => to_signed(28988, LUT_AMPL_WIDTH),
		11326 => to_signed(28989, LUT_AMPL_WIDTH),
		11327 => to_signed(28991, LUT_AMPL_WIDTH),
		11328 => to_signed(28992, LUT_AMPL_WIDTH),
		11329 => to_signed(28994, LUT_AMPL_WIDTH),
		11330 => to_signed(28995, LUT_AMPL_WIDTH),
		11331 => to_signed(28997, LUT_AMPL_WIDTH),
		11332 => to_signed(28998, LUT_AMPL_WIDTH),
		11333 => to_signed(28999, LUT_AMPL_WIDTH),
		11334 => to_signed(29001, LUT_AMPL_WIDTH),
		11335 => to_signed(29002, LUT_AMPL_WIDTH),
		11336 => to_signed(29004, LUT_AMPL_WIDTH),
		11337 => to_signed(29005, LUT_AMPL_WIDTH),
		11338 => to_signed(29007, LUT_AMPL_WIDTH),
		11339 => to_signed(29008, LUT_AMPL_WIDTH),
		11340 => to_signed(29010, LUT_AMPL_WIDTH),
		11341 => to_signed(29011, LUT_AMPL_WIDTH),
		11342 => to_signed(29013, LUT_AMPL_WIDTH),
		11343 => to_signed(29014, LUT_AMPL_WIDTH),
		11344 => to_signed(29016, LUT_AMPL_WIDTH),
		11345 => to_signed(29017, LUT_AMPL_WIDTH),
		11346 => to_signed(29018, LUT_AMPL_WIDTH),
		11347 => to_signed(29020, LUT_AMPL_WIDTH),
		11348 => to_signed(29021, LUT_AMPL_WIDTH),
		11349 => to_signed(29023, LUT_AMPL_WIDTH),
		11350 => to_signed(29024, LUT_AMPL_WIDTH),
		11351 => to_signed(29026, LUT_AMPL_WIDTH),
		11352 => to_signed(29027, LUT_AMPL_WIDTH),
		11353 => to_signed(29029, LUT_AMPL_WIDTH),
		11354 => to_signed(29030, LUT_AMPL_WIDTH),
		11355 => to_signed(29032, LUT_AMPL_WIDTH),
		11356 => to_signed(29033, LUT_AMPL_WIDTH),
		11357 => to_signed(29034, LUT_AMPL_WIDTH),
		11358 => to_signed(29036, LUT_AMPL_WIDTH),
		11359 => to_signed(29037, LUT_AMPL_WIDTH),
		11360 => to_signed(29039, LUT_AMPL_WIDTH),
		11361 => to_signed(29040, LUT_AMPL_WIDTH),
		11362 => to_signed(29042, LUT_AMPL_WIDTH),
		11363 => to_signed(29043, LUT_AMPL_WIDTH),
		11364 => to_signed(29045, LUT_AMPL_WIDTH),
		11365 => to_signed(29046, LUT_AMPL_WIDTH),
		11366 => to_signed(29048, LUT_AMPL_WIDTH),
		11367 => to_signed(29049, LUT_AMPL_WIDTH),
		11368 => to_signed(29050, LUT_AMPL_WIDTH),
		11369 => to_signed(29052, LUT_AMPL_WIDTH),
		11370 => to_signed(29053, LUT_AMPL_WIDTH),
		11371 => to_signed(29055, LUT_AMPL_WIDTH),
		11372 => to_signed(29056, LUT_AMPL_WIDTH),
		11373 => to_signed(29058, LUT_AMPL_WIDTH),
		11374 => to_signed(29059, LUT_AMPL_WIDTH),
		11375 => to_signed(29061, LUT_AMPL_WIDTH),
		11376 => to_signed(29062, LUT_AMPL_WIDTH),
		11377 => to_signed(29064, LUT_AMPL_WIDTH),
		11378 => to_signed(29065, LUT_AMPL_WIDTH),
		11379 => to_signed(29066, LUT_AMPL_WIDTH),
		11380 => to_signed(29068, LUT_AMPL_WIDTH),
		11381 => to_signed(29069, LUT_AMPL_WIDTH),
		11382 => to_signed(29071, LUT_AMPL_WIDTH),
		11383 => to_signed(29072, LUT_AMPL_WIDTH),
		11384 => to_signed(29074, LUT_AMPL_WIDTH),
		11385 => to_signed(29075, LUT_AMPL_WIDTH),
		11386 => to_signed(29077, LUT_AMPL_WIDTH),
		11387 => to_signed(29078, LUT_AMPL_WIDTH),
		11388 => to_signed(29079, LUT_AMPL_WIDTH),
		11389 => to_signed(29081, LUT_AMPL_WIDTH),
		11390 => to_signed(29082, LUT_AMPL_WIDTH),
		11391 => to_signed(29084, LUT_AMPL_WIDTH),
		11392 => to_signed(29085, LUT_AMPL_WIDTH),
		11393 => to_signed(29087, LUT_AMPL_WIDTH),
		11394 => to_signed(29088, LUT_AMPL_WIDTH),
		11395 => to_signed(29090, LUT_AMPL_WIDTH),
		11396 => to_signed(29091, LUT_AMPL_WIDTH),
		11397 => to_signed(29093, LUT_AMPL_WIDTH),
		11398 => to_signed(29094, LUT_AMPL_WIDTH),
		11399 => to_signed(29095, LUT_AMPL_WIDTH),
		11400 => to_signed(29097, LUT_AMPL_WIDTH),
		11401 => to_signed(29098, LUT_AMPL_WIDTH),
		11402 => to_signed(29100, LUT_AMPL_WIDTH),
		11403 => to_signed(29101, LUT_AMPL_WIDTH),
		11404 => to_signed(29103, LUT_AMPL_WIDTH),
		11405 => to_signed(29104, LUT_AMPL_WIDTH),
		11406 => to_signed(29106, LUT_AMPL_WIDTH),
		11407 => to_signed(29107, LUT_AMPL_WIDTH),
		11408 => to_signed(29108, LUT_AMPL_WIDTH),
		11409 => to_signed(29110, LUT_AMPL_WIDTH),
		11410 => to_signed(29111, LUT_AMPL_WIDTH),
		11411 => to_signed(29113, LUT_AMPL_WIDTH),
		11412 => to_signed(29114, LUT_AMPL_WIDTH),
		11413 => to_signed(29116, LUT_AMPL_WIDTH),
		11414 => to_signed(29117, LUT_AMPL_WIDTH),
		11415 => to_signed(29118, LUT_AMPL_WIDTH),
		11416 => to_signed(29120, LUT_AMPL_WIDTH),
		11417 => to_signed(29121, LUT_AMPL_WIDTH),
		11418 => to_signed(29123, LUT_AMPL_WIDTH),
		11419 => to_signed(29124, LUT_AMPL_WIDTH),
		11420 => to_signed(29126, LUT_AMPL_WIDTH),
		11421 => to_signed(29127, LUT_AMPL_WIDTH),
		11422 => to_signed(29129, LUT_AMPL_WIDTH),
		11423 => to_signed(29130, LUT_AMPL_WIDTH),
		11424 => to_signed(29131, LUT_AMPL_WIDTH),
		11425 => to_signed(29133, LUT_AMPL_WIDTH),
		11426 => to_signed(29134, LUT_AMPL_WIDTH),
		11427 => to_signed(29136, LUT_AMPL_WIDTH),
		11428 => to_signed(29137, LUT_AMPL_WIDTH),
		11429 => to_signed(29139, LUT_AMPL_WIDTH),
		11430 => to_signed(29140, LUT_AMPL_WIDTH),
		11431 => to_signed(29142, LUT_AMPL_WIDTH),
		11432 => to_signed(29143, LUT_AMPL_WIDTH),
		11433 => to_signed(29144, LUT_AMPL_WIDTH),
		11434 => to_signed(29146, LUT_AMPL_WIDTH),
		11435 => to_signed(29147, LUT_AMPL_WIDTH),
		11436 => to_signed(29149, LUT_AMPL_WIDTH),
		11437 => to_signed(29150, LUT_AMPL_WIDTH),
		11438 => to_signed(29152, LUT_AMPL_WIDTH),
		11439 => to_signed(29153, LUT_AMPL_WIDTH),
		11440 => to_signed(29154, LUT_AMPL_WIDTH),
		11441 => to_signed(29156, LUT_AMPL_WIDTH),
		11442 => to_signed(29157, LUT_AMPL_WIDTH),
		11443 => to_signed(29159, LUT_AMPL_WIDTH),
		11444 => to_signed(29160, LUT_AMPL_WIDTH),
		11445 => to_signed(29162, LUT_AMPL_WIDTH),
		11446 => to_signed(29163, LUT_AMPL_WIDTH),
		11447 => to_signed(29164, LUT_AMPL_WIDTH),
		11448 => to_signed(29166, LUT_AMPL_WIDTH),
		11449 => to_signed(29167, LUT_AMPL_WIDTH),
		11450 => to_signed(29169, LUT_AMPL_WIDTH),
		11451 => to_signed(29170, LUT_AMPL_WIDTH),
		11452 => to_signed(29172, LUT_AMPL_WIDTH),
		11453 => to_signed(29173, LUT_AMPL_WIDTH),
		11454 => to_signed(29174, LUT_AMPL_WIDTH),
		11455 => to_signed(29176, LUT_AMPL_WIDTH),
		11456 => to_signed(29177, LUT_AMPL_WIDTH),
		11457 => to_signed(29179, LUT_AMPL_WIDTH),
		11458 => to_signed(29180, LUT_AMPL_WIDTH),
		11459 => to_signed(29182, LUT_AMPL_WIDTH),
		11460 => to_signed(29183, LUT_AMPL_WIDTH),
		11461 => to_signed(29184, LUT_AMPL_WIDTH),
		11462 => to_signed(29186, LUT_AMPL_WIDTH),
		11463 => to_signed(29187, LUT_AMPL_WIDTH),
		11464 => to_signed(29189, LUT_AMPL_WIDTH),
		11465 => to_signed(29190, LUT_AMPL_WIDTH),
		11466 => to_signed(29192, LUT_AMPL_WIDTH),
		11467 => to_signed(29193, LUT_AMPL_WIDTH),
		11468 => to_signed(29194, LUT_AMPL_WIDTH),
		11469 => to_signed(29196, LUT_AMPL_WIDTH),
		11470 => to_signed(29197, LUT_AMPL_WIDTH),
		11471 => to_signed(29199, LUT_AMPL_WIDTH),
		11472 => to_signed(29200, LUT_AMPL_WIDTH),
		11473 => to_signed(29202, LUT_AMPL_WIDTH),
		11474 => to_signed(29203, LUT_AMPL_WIDTH),
		11475 => to_signed(29204, LUT_AMPL_WIDTH),
		11476 => to_signed(29206, LUT_AMPL_WIDTH),
		11477 => to_signed(29207, LUT_AMPL_WIDTH),
		11478 => to_signed(29209, LUT_AMPL_WIDTH),
		11479 => to_signed(29210, LUT_AMPL_WIDTH),
		11480 => to_signed(29212, LUT_AMPL_WIDTH),
		11481 => to_signed(29213, LUT_AMPL_WIDTH),
		11482 => to_signed(29214, LUT_AMPL_WIDTH),
		11483 => to_signed(29216, LUT_AMPL_WIDTH),
		11484 => to_signed(29217, LUT_AMPL_WIDTH),
		11485 => to_signed(29219, LUT_AMPL_WIDTH),
		11486 => to_signed(29220, LUT_AMPL_WIDTH),
		11487 => to_signed(29222, LUT_AMPL_WIDTH),
		11488 => to_signed(29223, LUT_AMPL_WIDTH),
		11489 => to_signed(29224, LUT_AMPL_WIDTH),
		11490 => to_signed(29226, LUT_AMPL_WIDTH),
		11491 => to_signed(29227, LUT_AMPL_WIDTH),
		11492 => to_signed(29229, LUT_AMPL_WIDTH),
		11493 => to_signed(29230, LUT_AMPL_WIDTH),
		11494 => to_signed(29231, LUT_AMPL_WIDTH),
		11495 => to_signed(29233, LUT_AMPL_WIDTH),
		11496 => to_signed(29234, LUT_AMPL_WIDTH),
		11497 => to_signed(29236, LUT_AMPL_WIDTH),
		11498 => to_signed(29237, LUT_AMPL_WIDTH),
		11499 => to_signed(29239, LUT_AMPL_WIDTH),
		11500 => to_signed(29240, LUT_AMPL_WIDTH),
		11501 => to_signed(29241, LUT_AMPL_WIDTH),
		11502 => to_signed(29243, LUT_AMPL_WIDTH),
		11503 => to_signed(29244, LUT_AMPL_WIDTH),
		11504 => to_signed(29246, LUT_AMPL_WIDTH),
		11505 => to_signed(29247, LUT_AMPL_WIDTH),
		11506 => to_signed(29248, LUT_AMPL_WIDTH),
		11507 => to_signed(29250, LUT_AMPL_WIDTH),
		11508 => to_signed(29251, LUT_AMPL_WIDTH),
		11509 => to_signed(29253, LUT_AMPL_WIDTH),
		11510 => to_signed(29254, LUT_AMPL_WIDTH),
		11511 => to_signed(29256, LUT_AMPL_WIDTH),
		11512 => to_signed(29257, LUT_AMPL_WIDTH),
		11513 => to_signed(29258, LUT_AMPL_WIDTH),
		11514 => to_signed(29260, LUT_AMPL_WIDTH),
		11515 => to_signed(29261, LUT_AMPL_WIDTH),
		11516 => to_signed(29263, LUT_AMPL_WIDTH),
		11517 => to_signed(29264, LUT_AMPL_WIDTH),
		11518 => to_signed(29265, LUT_AMPL_WIDTH),
		11519 => to_signed(29267, LUT_AMPL_WIDTH),
		11520 => to_signed(29268, LUT_AMPL_WIDTH),
		11521 => to_signed(29270, LUT_AMPL_WIDTH),
		11522 => to_signed(29271, LUT_AMPL_WIDTH),
		11523 => to_signed(29273, LUT_AMPL_WIDTH),
		11524 => to_signed(29274, LUT_AMPL_WIDTH),
		11525 => to_signed(29275, LUT_AMPL_WIDTH),
		11526 => to_signed(29277, LUT_AMPL_WIDTH),
		11527 => to_signed(29278, LUT_AMPL_WIDTH),
		11528 => to_signed(29280, LUT_AMPL_WIDTH),
		11529 => to_signed(29281, LUT_AMPL_WIDTH),
		11530 => to_signed(29282, LUT_AMPL_WIDTH),
		11531 => to_signed(29284, LUT_AMPL_WIDTH),
		11532 => to_signed(29285, LUT_AMPL_WIDTH),
		11533 => to_signed(29287, LUT_AMPL_WIDTH),
		11534 => to_signed(29288, LUT_AMPL_WIDTH),
		11535 => to_signed(29289, LUT_AMPL_WIDTH),
		11536 => to_signed(29291, LUT_AMPL_WIDTH),
		11537 => to_signed(29292, LUT_AMPL_WIDTH),
		11538 => to_signed(29294, LUT_AMPL_WIDTH),
		11539 => to_signed(29295, LUT_AMPL_WIDTH),
		11540 => to_signed(29296, LUT_AMPL_WIDTH),
		11541 => to_signed(29298, LUT_AMPL_WIDTH),
		11542 => to_signed(29299, LUT_AMPL_WIDTH),
		11543 => to_signed(29301, LUT_AMPL_WIDTH),
		11544 => to_signed(29302, LUT_AMPL_WIDTH),
		11545 => to_signed(29304, LUT_AMPL_WIDTH),
		11546 => to_signed(29305, LUT_AMPL_WIDTH),
		11547 => to_signed(29306, LUT_AMPL_WIDTH),
		11548 => to_signed(29308, LUT_AMPL_WIDTH),
		11549 => to_signed(29309, LUT_AMPL_WIDTH),
		11550 => to_signed(29311, LUT_AMPL_WIDTH),
		11551 => to_signed(29312, LUT_AMPL_WIDTH),
		11552 => to_signed(29313, LUT_AMPL_WIDTH),
		11553 => to_signed(29315, LUT_AMPL_WIDTH),
		11554 => to_signed(29316, LUT_AMPL_WIDTH),
		11555 => to_signed(29318, LUT_AMPL_WIDTH),
		11556 => to_signed(29319, LUT_AMPL_WIDTH),
		11557 => to_signed(29320, LUT_AMPL_WIDTH),
		11558 => to_signed(29322, LUT_AMPL_WIDTH),
		11559 => to_signed(29323, LUT_AMPL_WIDTH),
		11560 => to_signed(29325, LUT_AMPL_WIDTH),
		11561 => to_signed(29326, LUT_AMPL_WIDTH),
		11562 => to_signed(29327, LUT_AMPL_WIDTH),
		11563 => to_signed(29329, LUT_AMPL_WIDTH),
		11564 => to_signed(29330, LUT_AMPL_WIDTH),
		11565 => to_signed(29332, LUT_AMPL_WIDTH),
		11566 => to_signed(29333, LUT_AMPL_WIDTH),
		11567 => to_signed(29334, LUT_AMPL_WIDTH),
		11568 => to_signed(29336, LUT_AMPL_WIDTH),
		11569 => to_signed(29337, LUT_AMPL_WIDTH),
		11570 => to_signed(29339, LUT_AMPL_WIDTH),
		11571 => to_signed(29340, LUT_AMPL_WIDTH),
		11572 => to_signed(29341, LUT_AMPL_WIDTH),
		11573 => to_signed(29343, LUT_AMPL_WIDTH),
		11574 => to_signed(29344, LUT_AMPL_WIDTH),
		11575 => to_signed(29346, LUT_AMPL_WIDTH),
		11576 => to_signed(29347, LUT_AMPL_WIDTH),
		11577 => to_signed(29348, LUT_AMPL_WIDTH),
		11578 => to_signed(29350, LUT_AMPL_WIDTH),
		11579 => to_signed(29351, LUT_AMPL_WIDTH),
		11580 => to_signed(29353, LUT_AMPL_WIDTH),
		11581 => to_signed(29354, LUT_AMPL_WIDTH),
		11582 => to_signed(29355, LUT_AMPL_WIDTH),
		11583 => to_signed(29357, LUT_AMPL_WIDTH),
		11584 => to_signed(29358, LUT_AMPL_WIDTH),
		11585 => to_signed(29360, LUT_AMPL_WIDTH),
		11586 => to_signed(29361, LUT_AMPL_WIDTH),
		11587 => to_signed(29362, LUT_AMPL_WIDTH),
		11588 => to_signed(29364, LUT_AMPL_WIDTH),
		11589 => to_signed(29365, LUT_AMPL_WIDTH),
		11590 => to_signed(29366, LUT_AMPL_WIDTH),
		11591 => to_signed(29368, LUT_AMPL_WIDTH),
		11592 => to_signed(29369, LUT_AMPL_WIDTH),
		11593 => to_signed(29371, LUT_AMPL_WIDTH),
		11594 => to_signed(29372, LUT_AMPL_WIDTH),
		11595 => to_signed(29373, LUT_AMPL_WIDTH),
		11596 => to_signed(29375, LUT_AMPL_WIDTH),
		11597 => to_signed(29376, LUT_AMPL_WIDTH),
		11598 => to_signed(29378, LUT_AMPL_WIDTH),
		11599 => to_signed(29379, LUT_AMPL_WIDTH),
		11600 => to_signed(29380, LUT_AMPL_WIDTH),
		11601 => to_signed(29382, LUT_AMPL_WIDTH),
		11602 => to_signed(29383, LUT_AMPL_WIDTH),
		11603 => to_signed(29385, LUT_AMPL_WIDTH),
		11604 => to_signed(29386, LUT_AMPL_WIDTH),
		11605 => to_signed(29387, LUT_AMPL_WIDTH),
		11606 => to_signed(29389, LUT_AMPL_WIDTH),
		11607 => to_signed(29390, LUT_AMPL_WIDTH),
		11608 => to_signed(29392, LUT_AMPL_WIDTH),
		11609 => to_signed(29393, LUT_AMPL_WIDTH),
		11610 => to_signed(29394, LUT_AMPL_WIDTH),
		11611 => to_signed(29396, LUT_AMPL_WIDTH),
		11612 => to_signed(29397, LUT_AMPL_WIDTH),
		11613 => to_signed(29398, LUT_AMPL_WIDTH),
		11614 => to_signed(29400, LUT_AMPL_WIDTH),
		11615 => to_signed(29401, LUT_AMPL_WIDTH),
		11616 => to_signed(29403, LUT_AMPL_WIDTH),
		11617 => to_signed(29404, LUT_AMPL_WIDTH),
		11618 => to_signed(29405, LUT_AMPL_WIDTH),
		11619 => to_signed(29407, LUT_AMPL_WIDTH),
		11620 => to_signed(29408, LUT_AMPL_WIDTH),
		11621 => to_signed(29410, LUT_AMPL_WIDTH),
		11622 => to_signed(29411, LUT_AMPL_WIDTH),
		11623 => to_signed(29412, LUT_AMPL_WIDTH),
		11624 => to_signed(29414, LUT_AMPL_WIDTH),
		11625 => to_signed(29415, LUT_AMPL_WIDTH),
		11626 => to_signed(29416, LUT_AMPL_WIDTH),
		11627 => to_signed(29418, LUT_AMPL_WIDTH),
		11628 => to_signed(29419, LUT_AMPL_WIDTH),
		11629 => to_signed(29421, LUT_AMPL_WIDTH),
		11630 => to_signed(29422, LUT_AMPL_WIDTH),
		11631 => to_signed(29423, LUT_AMPL_WIDTH),
		11632 => to_signed(29425, LUT_AMPL_WIDTH),
		11633 => to_signed(29426, LUT_AMPL_WIDTH),
		11634 => to_signed(29428, LUT_AMPL_WIDTH),
		11635 => to_signed(29429, LUT_AMPL_WIDTH),
		11636 => to_signed(29430, LUT_AMPL_WIDTH),
		11637 => to_signed(29432, LUT_AMPL_WIDTH),
		11638 => to_signed(29433, LUT_AMPL_WIDTH),
		11639 => to_signed(29434, LUT_AMPL_WIDTH),
		11640 => to_signed(29436, LUT_AMPL_WIDTH),
		11641 => to_signed(29437, LUT_AMPL_WIDTH),
		11642 => to_signed(29439, LUT_AMPL_WIDTH),
		11643 => to_signed(29440, LUT_AMPL_WIDTH),
		11644 => to_signed(29441, LUT_AMPL_WIDTH),
		11645 => to_signed(29443, LUT_AMPL_WIDTH),
		11646 => to_signed(29444, LUT_AMPL_WIDTH),
		11647 => to_signed(29445, LUT_AMPL_WIDTH),
		11648 => to_signed(29447, LUT_AMPL_WIDTH),
		11649 => to_signed(29448, LUT_AMPL_WIDTH),
		11650 => to_signed(29450, LUT_AMPL_WIDTH),
		11651 => to_signed(29451, LUT_AMPL_WIDTH),
		11652 => to_signed(29452, LUT_AMPL_WIDTH),
		11653 => to_signed(29454, LUT_AMPL_WIDTH),
		11654 => to_signed(29455, LUT_AMPL_WIDTH),
		11655 => to_signed(29457, LUT_AMPL_WIDTH),
		11656 => to_signed(29458, LUT_AMPL_WIDTH),
		11657 => to_signed(29459, LUT_AMPL_WIDTH),
		11658 => to_signed(29461, LUT_AMPL_WIDTH),
		11659 => to_signed(29462, LUT_AMPL_WIDTH),
		11660 => to_signed(29463, LUT_AMPL_WIDTH),
		11661 => to_signed(29465, LUT_AMPL_WIDTH),
		11662 => to_signed(29466, LUT_AMPL_WIDTH),
		11663 => to_signed(29468, LUT_AMPL_WIDTH),
		11664 => to_signed(29469, LUT_AMPL_WIDTH),
		11665 => to_signed(29470, LUT_AMPL_WIDTH),
		11666 => to_signed(29472, LUT_AMPL_WIDTH),
		11667 => to_signed(29473, LUT_AMPL_WIDTH),
		11668 => to_signed(29474, LUT_AMPL_WIDTH),
		11669 => to_signed(29476, LUT_AMPL_WIDTH),
		11670 => to_signed(29477, LUT_AMPL_WIDTH),
		11671 => to_signed(29478, LUT_AMPL_WIDTH),
		11672 => to_signed(29480, LUT_AMPL_WIDTH),
		11673 => to_signed(29481, LUT_AMPL_WIDTH),
		11674 => to_signed(29483, LUT_AMPL_WIDTH),
		11675 => to_signed(29484, LUT_AMPL_WIDTH),
		11676 => to_signed(29485, LUT_AMPL_WIDTH),
		11677 => to_signed(29487, LUT_AMPL_WIDTH),
		11678 => to_signed(29488, LUT_AMPL_WIDTH),
		11679 => to_signed(29489, LUT_AMPL_WIDTH),
		11680 => to_signed(29491, LUT_AMPL_WIDTH),
		11681 => to_signed(29492, LUT_AMPL_WIDTH),
		11682 => to_signed(29494, LUT_AMPL_WIDTH),
		11683 => to_signed(29495, LUT_AMPL_WIDTH),
		11684 => to_signed(29496, LUT_AMPL_WIDTH),
		11685 => to_signed(29498, LUT_AMPL_WIDTH),
		11686 => to_signed(29499, LUT_AMPL_WIDTH),
		11687 => to_signed(29500, LUT_AMPL_WIDTH),
		11688 => to_signed(29502, LUT_AMPL_WIDTH),
		11689 => to_signed(29503, LUT_AMPL_WIDTH),
		11690 => to_signed(29504, LUT_AMPL_WIDTH),
		11691 => to_signed(29506, LUT_AMPL_WIDTH),
		11692 => to_signed(29507, LUT_AMPL_WIDTH),
		11693 => to_signed(29509, LUT_AMPL_WIDTH),
		11694 => to_signed(29510, LUT_AMPL_WIDTH),
		11695 => to_signed(29511, LUT_AMPL_WIDTH),
		11696 => to_signed(29513, LUT_AMPL_WIDTH),
		11697 => to_signed(29514, LUT_AMPL_WIDTH),
		11698 => to_signed(29515, LUT_AMPL_WIDTH),
		11699 => to_signed(29517, LUT_AMPL_WIDTH),
		11700 => to_signed(29518, LUT_AMPL_WIDTH),
		11701 => to_signed(29520, LUT_AMPL_WIDTH),
		11702 => to_signed(29521, LUT_AMPL_WIDTH),
		11703 => to_signed(29522, LUT_AMPL_WIDTH),
		11704 => to_signed(29524, LUT_AMPL_WIDTH),
		11705 => to_signed(29525, LUT_AMPL_WIDTH),
		11706 => to_signed(29526, LUT_AMPL_WIDTH),
		11707 => to_signed(29528, LUT_AMPL_WIDTH),
		11708 => to_signed(29529, LUT_AMPL_WIDTH),
		11709 => to_signed(29530, LUT_AMPL_WIDTH),
		11710 => to_signed(29532, LUT_AMPL_WIDTH),
		11711 => to_signed(29533, LUT_AMPL_WIDTH),
		11712 => to_signed(29534, LUT_AMPL_WIDTH),
		11713 => to_signed(29536, LUT_AMPL_WIDTH),
		11714 => to_signed(29537, LUT_AMPL_WIDTH),
		11715 => to_signed(29539, LUT_AMPL_WIDTH),
		11716 => to_signed(29540, LUT_AMPL_WIDTH),
		11717 => to_signed(29541, LUT_AMPL_WIDTH),
		11718 => to_signed(29543, LUT_AMPL_WIDTH),
		11719 => to_signed(29544, LUT_AMPL_WIDTH),
		11720 => to_signed(29545, LUT_AMPL_WIDTH),
		11721 => to_signed(29547, LUT_AMPL_WIDTH),
		11722 => to_signed(29548, LUT_AMPL_WIDTH),
		11723 => to_signed(29549, LUT_AMPL_WIDTH),
		11724 => to_signed(29551, LUT_AMPL_WIDTH),
		11725 => to_signed(29552, LUT_AMPL_WIDTH),
		11726 => to_signed(29554, LUT_AMPL_WIDTH),
		11727 => to_signed(29555, LUT_AMPL_WIDTH),
		11728 => to_signed(29556, LUT_AMPL_WIDTH),
		11729 => to_signed(29558, LUT_AMPL_WIDTH),
		11730 => to_signed(29559, LUT_AMPL_WIDTH),
		11731 => to_signed(29560, LUT_AMPL_WIDTH),
		11732 => to_signed(29562, LUT_AMPL_WIDTH),
		11733 => to_signed(29563, LUT_AMPL_WIDTH),
		11734 => to_signed(29564, LUT_AMPL_WIDTH),
		11735 => to_signed(29566, LUT_AMPL_WIDTH),
		11736 => to_signed(29567, LUT_AMPL_WIDTH),
		11737 => to_signed(29568, LUT_AMPL_WIDTH),
		11738 => to_signed(29570, LUT_AMPL_WIDTH),
		11739 => to_signed(29571, LUT_AMPL_WIDTH),
		11740 => to_signed(29572, LUT_AMPL_WIDTH),
		11741 => to_signed(29574, LUT_AMPL_WIDTH),
		11742 => to_signed(29575, LUT_AMPL_WIDTH),
		11743 => to_signed(29577, LUT_AMPL_WIDTH),
		11744 => to_signed(29578, LUT_AMPL_WIDTH),
		11745 => to_signed(29579, LUT_AMPL_WIDTH),
		11746 => to_signed(29581, LUT_AMPL_WIDTH),
		11747 => to_signed(29582, LUT_AMPL_WIDTH),
		11748 => to_signed(29583, LUT_AMPL_WIDTH),
		11749 => to_signed(29585, LUT_AMPL_WIDTH),
		11750 => to_signed(29586, LUT_AMPL_WIDTH),
		11751 => to_signed(29587, LUT_AMPL_WIDTH),
		11752 => to_signed(29589, LUT_AMPL_WIDTH),
		11753 => to_signed(29590, LUT_AMPL_WIDTH),
		11754 => to_signed(29591, LUT_AMPL_WIDTH),
		11755 => to_signed(29593, LUT_AMPL_WIDTH),
		11756 => to_signed(29594, LUT_AMPL_WIDTH),
		11757 => to_signed(29595, LUT_AMPL_WIDTH),
		11758 => to_signed(29597, LUT_AMPL_WIDTH),
		11759 => to_signed(29598, LUT_AMPL_WIDTH),
		11760 => to_signed(29599, LUT_AMPL_WIDTH),
		11761 => to_signed(29601, LUT_AMPL_WIDTH),
		11762 => to_signed(29602, LUT_AMPL_WIDTH),
		11763 => to_signed(29604, LUT_AMPL_WIDTH),
		11764 => to_signed(29605, LUT_AMPL_WIDTH),
		11765 => to_signed(29606, LUT_AMPL_WIDTH),
		11766 => to_signed(29608, LUT_AMPL_WIDTH),
		11767 => to_signed(29609, LUT_AMPL_WIDTH),
		11768 => to_signed(29610, LUT_AMPL_WIDTH),
		11769 => to_signed(29612, LUT_AMPL_WIDTH),
		11770 => to_signed(29613, LUT_AMPL_WIDTH),
		11771 => to_signed(29614, LUT_AMPL_WIDTH),
		11772 => to_signed(29616, LUT_AMPL_WIDTH),
		11773 => to_signed(29617, LUT_AMPL_WIDTH),
		11774 => to_signed(29618, LUT_AMPL_WIDTH),
		11775 => to_signed(29620, LUT_AMPL_WIDTH),
		11776 => to_signed(29621, LUT_AMPL_WIDTH),
		11777 => to_signed(29622, LUT_AMPL_WIDTH),
		11778 => to_signed(29624, LUT_AMPL_WIDTH),
		11779 => to_signed(29625, LUT_AMPL_WIDTH),
		11780 => to_signed(29626, LUT_AMPL_WIDTH),
		11781 => to_signed(29628, LUT_AMPL_WIDTH),
		11782 => to_signed(29629, LUT_AMPL_WIDTH),
		11783 => to_signed(29630, LUT_AMPL_WIDTH),
		11784 => to_signed(29632, LUT_AMPL_WIDTH),
		11785 => to_signed(29633, LUT_AMPL_WIDTH),
		11786 => to_signed(29634, LUT_AMPL_WIDTH),
		11787 => to_signed(29636, LUT_AMPL_WIDTH),
		11788 => to_signed(29637, LUT_AMPL_WIDTH),
		11789 => to_signed(29638, LUT_AMPL_WIDTH),
		11790 => to_signed(29640, LUT_AMPL_WIDTH),
		11791 => to_signed(29641, LUT_AMPL_WIDTH),
		11792 => to_signed(29642, LUT_AMPL_WIDTH),
		11793 => to_signed(29644, LUT_AMPL_WIDTH),
		11794 => to_signed(29645, LUT_AMPL_WIDTH),
		11795 => to_signed(29646, LUT_AMPL_WIDTH),
		11796 => to_signed(29648, LUT_AMPL_WIDTH),
		11797 => to_signed(29649, LUT_AMPL_WIDTH),
		11798 => to_signed(29651, LUT_AMPL_WIDTH),
		11799 => to_signed(29652, LUT_AMPL_WIDTH),
		11800 => to_signed(29653, LUT_AMPL_WIDTH),
		11801 => to_signed(29655, LUT_AMPL_WIDTH),
		11802 => to_signed(29656, LUT_AMPL_WIDTH),
		11803 => to_signed(29657, LUT_AMPL_WIDTH),
		11804 => to_signed(29659, LUT_AMPL_WIDTH),
		11805 => to_signed(29660, LUT_AMPL_WIDTH),
		11806 => to_signed(29661, LUT_AMPL_WIDTH),
		11807 => to_signed(29663, LUT_AMPL_WIDTH),
		11808 => to_signed(29664, LUT_AMPL_WIDTH),
		11809 => to_signed(29665, LUT_AMPL_WIDTH),
		11810 => to_signed(29667, LUT_AMPL_WIDTH),
		11811 => to_signed(29668, LUT_AMPL_WIDTH),
		11812 => to_signed(29669, LUT_AMPL_WIDTH),
		11813 => to_signed(29671, LUT_AMPL_WIDTH),
		11814 => to_signed(29672, LUT_AMPL_WIDTH),
		11815 => to_signed(29673, LUT_AMPL_WIDTH),
		11816 => to_signed(29675, LUT_AMPL_WIDTH),
		11817 => to_signed(29676, LUT_AMPL_WIDTH),
		11818 => to_signed(29677, LUT_AMPL_WIDTH),
		11819 => to_signed(29679, LUT_AMPL_WIDTH),
		11820 => to_signed(29680, LUT_AMPL_WIDTH),
		11821 => to_signed(29681, LUT_AMPL_WIDTH),
		11822 => to_signed(29683, LUT_AMPL_WIDTH),
		11823 => to_signed(29684, LUT_AMPL_WIDTH),
		11824 => to_signed(29685, LUT_AMPL_WIDTH),
		11825 => to_signed(29687, LUT_AMPL_WIDTH),
		11826 => to_signed(29688, LUT_AMPL_WIDTH),
		11827 => to_signed(29689, LUT_AMPL_WIDTH),
		11828 => to_signed(29690, LUT_AMPL_WIDTH),
		11829 => to_signed(29692, LUT_AMPL_WIDTH),
		11830 => to_signed(29693, LUT_AMPL_WIDTH),
		11831 => to_signed(29694, LUT_AMPL_WIDTH),
		11832 => to_signed(29696, LUT_AMPL_WIDTH),
		11833 => to_signed(29697, LUT_AMPL_WIDTH),
		11834 => to_signed(29698, LUT_AMPL_WIDTH),
		11835 => to_signed(29700, LUT_AMPL_WIDTH),
		11836 => to_signed(29701, LUT_AMPL_WIDTH),
		11837 => to_signed(29702, LUT_AMPL_WIDTH),
		11838 => to_signed(29704, LUT_AMPL_WIDTH),
		11839 => to_signed(29705, LUT_AMPL_WIDTH),
		11840 => to_signed(29706, LUT_AMPL_WIDTH),
		11841 => to_signed(29708, LUT_AMPL_WIDTH),
		11842 => to_signed(29709, LUT_AMPL_WIDTH),
		11843 => to_signed(29710, LUT_AMPL_WIDTH),
		11844 => to_signed(29712, LUT_AMPL_WIDTH),
		11845 => to_signed(29713, LUT_AMPL_WIDTH),
		11846 => to_signed(29714, LUT_AMPL_WIDTH),
		11847 => to_signed(29716, LUT_AMPL_WIDTH),
		11848 => to_signed(29717, LUT_AMPL_WIDTH),
		11849 => to_signed(29718, LUT_AMPL_WIDTH),
		11850 => to_signed(29720, LUT_AMPL_WIDTH),
		11851 => to_signed(29721, LUT_AMPL_WIDTH),
		11852 => to_signed(29722, LUT_AMPL_WIDTH),
		11853 => to_signed(29724, LUT_AMPL_WIDTH),
		11854 => to_signed(29725, LUT_AMPL_WIDTH),
		11855 => to_signed(29726, LUT_AMPL_WIDTH),
		11856 => to_signed(29728, LUT_AMPL_WIDTH),
		11857 => to_signed(29729, LUT_AMPL_WIDTH),
		11858 => to_signed(29730, LUT_AMPL_WIDTH),
		11859 => to_signed(29732, LUT_AMPL_WIDTH),
		11860 => to_signed(29733, LUT_AMPL_WIDTH),
		11861 => to_signed(29734, LUT_AMPL_WIDTH),
		11862 => to_signed(29736, LUT_AMPL_WIDTH),
		11863 => to_signed(29737, LUT_AMPL_WIDTH),
		11864 => to_signed(29738, LUT_AMPL_WIDTH),
		11865 => to_signed(29739, LUT_AMPL_WIDTH),
		11866 => to_signed(29741, LUT_AMPL_WIDTH),
		11867 => to_signed(29742, LUT_AMPL_WIDTH),
		11868 => to_signed(29743, LUT_AMPL_WIDTH),
		11869 => to_signed(29745, LUT_AMPL_WIDTH),
		11870 => to_signed(29746, LUT_AMPL_WIDTH),
		11871 => to_signed(29747, LUT_AMPL_WIDTH),
		11872 => to_signed(29749, LUT_AMPL_WIDTH),
		11873 => to_signed(29750, LUT_AMPL_WIDTH),
		11874 => to_signed(29751, LUT_AMPL_WIDTH),
		11875 => to_signed(29753, LUT_AMPL_WIDTH),
		11876 => to_signed(29754, LUT_AMPL_WIDTH),
		11877 => to_signed(29755, LUT_AMPL_WIDTH),
		11878 => to_signed(29757, LUT_AMPL_WIDTH),
		11879 => to_signed(29758, LUT_AMPL_WIDTH),
		11880 => to_signed(29759, LUT_AMPL_WIDTH),
		11881 => to_signed(29761, LUT_AMPL_WIDTH),
		11882 => to_signed(29762, LUT_AMPL_WIDTH),
		11883 => to_signed(29763, LUT_AMPL_WIDTH),
		11884 => to_signed(29764, LUT_AMPL_WIDTH),
		11885 => to_signed(29766, LUT_AMPL_WIDTH),
		11886 => to_signed(29767, LUT_AMPL_WIDTH),
		11887 => to_signed(29768, LUT_AMPL_WIDTH),
		11888 => to_signed(29770, LUT_AMPL_WIDTH),
		11889 => to_signed(29771, LUT_AMPL_WIDTH),
		11890 => to_signed(29772, LUT_AMPL_WIDTH),
		11891 => to_signed(29774, LUT_AMPL_WIDTH),
		11892 => to_signed(29775, LUT_AMPL_WIDTH),
		11893 => to_signed(29776, LUT_AMPL_WIDTH),
		11894 => to_signed(29778, LUT_AMPL_WIDTH),
		11895 => to_signed(29779, LUT_AMPL_WIDTH),
		11896 => to_signed(29780, LUT_AMPL_WIDTH),
		11897 => to_signed(29782, LUT_AMPL_WIDTH),
		11898 => to_signed(29783, LUT_AMPL_WIDTH),
		11899 => to_signed(29784, LUT_AMPL_WIDTH),
		11900 => to_signed(29785, LUT_AMPL_WIDTH),
		11901 => to_signed(29787, LUT_AMPL_WIDTH),
		11902 => to_signed(29788, LUT_AMPL_WIDTH),
		11903 => to_signed(29789, LUT_AMPL_WIDTH),
		11904 => to_signed(29791, LUT_AMPL_WIDTH),
		11905 => to_signed(29792, LUT_AMPL_WIDTH),
		11906 => to_signed(29793, LUT_AMPL_WIDTH),
		11907 => to_signed(29795, LUT_AMPL_WIDTH),
		11908 => to_signed(29796, LUT_AMPL_WIDTH),
		11909 => to_signed(29797, LUT_AMPL_WIDTH),
		11910 => to_signed(29799, LUT_AMPL_WIDTH),
		11911 => to_signed(29800, LUT_AMPL_WIDTH),
		11912 => to_signed(29801, LUT_AMPL_WIDTH),
		11913 => to_signed(29802, LUT_AMPL_WIDTH),
		11914 => to_signed(29804, LUT_AMPL_WIDTH),
		11915 => to_signed(29805, LUT_AMPL_WIDTH),
		11916 => to_signed(29806, LUT_AMPL_WIDTH),
		11917 => to_signed(29808, LUT_AMPL_WIDTH),
		11918 => to_signed(29809, LUT_AMPL_WIDTH),
		11919 => to_signed(29810, LUT_AMPL_WIDTH),
		11920 => to_signed(29812, LUT_AMPL_WIDTH),
		11921 => to_signed(29813, LUT_AMPL_WIDTH),
		11922 => to_signed(29814, LUT_AMPL_WIDTH),
		11923 => to_signed(29816, LUT_AMPL_WIDTH),
		11924 => to_signed(29817, LUT_AMPL_WIDTH),
		11925 => to_signed(29818, LUT_AMPL_WIDTH),
		11926 => to_signed(29819, LUT_AMPL_WIDTH),
		11927 => to_signed(29821, LUT_AMPL_WIDTH),
		11928 => to_signed(29822, LUT_AMPL_WIDTH),
		11929 => to_signed(29823, LUT_AMPL_WIDTH),
		11930 => to_signed(29825, LUT_AMPL_WIDTH),
		11931 => to_signed(29826, LUT_AMPL_WIDTH),
		11932 => to_signed(29827, LUT_AMPL_WIDTH),
		11933 => to_signed(29829, LUT_AMPL_WIDTH),
		11934 => to_signed(29830, LUT_AMPL_WIDTH),
		11935 => to_signed(29831, LUT_AMPL_WIDTH),
		11936 => to_signed(29832, LUT_AMPL_WIDTH),
		11937 => to_signed(29834, LUT_AMPL_WIDTH),
		11938 => to_signed(29835, LUT_AMPL_WIDTH),
		11939 => to_signed(29836, LUT_AMPL_WIDTH),
		11940 => to_signed(29838, LUT_AMPL_WIDTH),
		11941 => to_signed(29839, LUT_AMPL_WIDTH),
		11942 => to_signed(29840, LUT_AMPL_WIDTH),
		11943 => to_signed(29842, LUT_AMPL_WIDTH),
		11944 => to_signed(29843, LUT_AMPL_WIDTH),
		11945 => to_signed(29844, LUT_AMPL_WIDTH),
		11946 => to_signed(29845, LUT_AMPL_WIDTH),
		11947 => to_signed(29847, LUT_AMPL_WIDTH),
		11948 => to_signed(29848, LUT_AMPL_WIDTH),
		11949 => to_signed(29849, LUT_AMPL_WIDTH),
		11950 => to_signed(29851, LUT_AMPL_WIDTH),
		11951 => to_signed(29852, LUT_AMPL_WIDTH),
		11952 => to_signed(29853, LUT_AMPL_WIDTH),
		11953 => to_signed(29854, LUT_AMPL_WIDTH),
		11954 => to_signed(29856, LUT_AMPL_WIDTH),
		11955 => to_signed(29857, LUT_AMPL_WIDTH),
		11956 => to_signed(29858, LUT_AMPL_WIDTH),
		11957 => to_signed(29860, LUT_AMPL_WIDTH),
		11958 => to_signed(29861, LUT_AMPL_WIDTH),
		11959 => to_signed(29862, LUT_AMPL_WIDTH),
		11960 => to_signed(29864, LUT_AMPL_WIDTH),
		11961 => to_signed(29865, LUT_AMPL_WIDTH),
		11962 => to_signed(29866, LUT_AMPL_WIDTH),
		11963 => to_signed(29867, LUT_AMPL_WIDTH),
		11964 => to_signed(29869, LUT_AMPL_WIDTH),
		11965 => to_signed(29870, LUT_AMPL_WIDTH),
		11966 => to_signed(29871, LUT_AMPL_WIDTH),
		11967 => to_signed(29873, LUT_AMPL_WIDTH),
		11968 => to_signed(29874, LUT_AMPL_WIDTH),
		11969 => to_signed(29875, LUT_AMPL_WIDTH),
		11970 => to_signed(29876, LUT_AMPL_WIDTH),
		11971 => to_signed(29878, LUT_AMPL_WIDTH),
		11972 => to_signed(29879, LUT_AMPL_WIDTH),
		11973 => to_signed(29880, LUT_AMPL_WIDTH),
		11974 => to_signed(29882, LUT_AMPL_WIDTH),
		11975 => to_signed(29883, LUT_AMPL_WIDTH),
		11976 => to_signed(29884, LUT_AMPL_WIDTH),
		11977 => to_signed(29885, LUT_AMPL_WIDTH),
		11978 => to_signed(29887, LUT_AMPL_WIDTH),
		11979 => to_signed(29888, LUT_AMPL_WIDTH),
		11980 => to_signed(29889, LUT_AMPL_WIDTH),
		11981 => to_signed(29891, LUT_AMPL_WIDTH),
		11982 => to_signed(29892, LUT_AMPL_WIDTH),
		11983 => to_signed(29893, LUT_AMPL_WIDTH),
		11984 => to_signed(29894, LUT_AMPL_WIDTH),
		11985 => to_signed(29896, LUT_AMPL_WIDTH),
		11986 => to_signed(29897, LUT_AMPL_WIDTH),
		11987 => to_signed(29898, LUT_AMPL_WIDTH),
		11988 => to_signed(29900, LUT_AMPL_WIDTH),
		11989 => to_signed(29901, LUT_AMPL_WIDTH),
		11990 => to_signed(29902, LUT_AMPL_WIDTH),
		11991 => to_signed(29903, LUT_AMPL_WIDTH),
		11992 => to_signed(29905, LUT_AMPL_WIDTH),
		11993 => to_signed(29906, LUT_AMPL_WIDTH),
		11994 => to_signed(29907, LUT_AMPL_WIDTH),
		11995 => to_signed(29909, LUT_AMPL_WIDTH),
		11996 => to_signed(29910, LUT_AMPL_WIDTH),
		11997 => to_signed(29911, LUT_AMPL_WIDTH),
		11998 => to_signed(29912, LUT_AMPL_WIDTH),
		11999 => to_signed(29914, LUT_AMPL_WIDTH),
		12000 => to_signed(29915, LUT_AMPL_WIDTH),
		12001 => to_signed(29916, LUT_AMPL_WIDTH),
		12002 => to_signed(29918, LUT_AMPL_WIDTH),
		12003 => to_signed(29919, LUT_AMPL_WIDTH),
		12004 => to_signed(29920, LUT_AMPL_WIDTH),
		12005 => to_signed(29921, LUT_AMPL_WIDTH),
		12006 => to_signed(29923, LUT_AMPL_WIDTH),
		12007 => to_signed(29924, LUT_AMPL_WIDTH),
		12008 => to_signed(29925, LUT_AMPL_WIDTH),
		12009 => to_signed(29927, LUT_AMPL_WIDTH),
		12010 => to_signed(29928, LUT_AMPL_WIDTH),
		12011 => to_signed(29929, LUT_AMPL_WIDTH),
		12012 => to_signed(29930, LUT_AMPL_WIDTH),
		12013 => to_signed(29932, LUT_AMPL_WIDTH),
		12014 => to_signed(29933, LUT_AMPL_WIDTH),
		12015 => to_signed(29934, LUT_AMPL_WIDTH),
		12016 => to_signed(29936, LUT_AMPL_WIDTH),
		12017 => to_signed(29937, LUT_AMPL_WIDTH),
		12018 => to_signed(29938, LUT_AMPL_WIDTH),
		12019 => to_signed(29939, LUT_AMPL_WIDTH),
		12020 => to_signed(29941, LUT_AMPL_WIDTH),
		12021 => to_signed(29942, LUT_AMPL_WIDTH),
		12022 => to_signed(29943, LUT_AMPL_WIDTH),
		12023 => to_signed(29944, LUT_AMPL_WIDTH),
		12024 => to_signed(29946, LUT_AMPL_WIDTH),
		12025 => to_signed(29947, LUT_AMPL_WIDTH),
		12026 => to_signed(29948, LUT_AMPL_WIDTH),
		12027 => to_signed(29950, LUT_AMPL_WIDTH),
		12028 => to_signed(29951, LUT_AMPL_WIDTH),
		12029 => to_signed(29952, LUT_AMPL_WIDTH),
		12030 => to_signed(29953, LUT_AMPL_WIDTH),
		12031 => to_signed(29955, LUT_AMPL_WIDTH),
		12032 => to_signed(29956, LUT_AMPL_WIDTH),
		12033 => to_signed(29957, LUT_AMPL_WIDTH),
		12034 => to_signed(29958, LUT_AMPL_WIDTH),
		12035 => to_signed(29960, LUT_AMPL_WIDTH),
		12036 => to_signed(29961, LUT_AMPL_WIDTH),
		12037 => to_signed(29962, LUT_AMPL_WIDTH),
		12038 => to_signed(29964, LUT_AMPL_WIDTH),
		12039 => to_signed(29965, LUT_AMPL_WIDTH),
		12040 => to_signed(29966, LUT_AMPL_WIDTH),
		12041 => to_signed(29967, LUT_AMPL_WIDTH),
		12042 => to_signed(29969, LUT_AMPL_WIDTH),
		12043 => to_signed(29970, LUT_AMPL_WIDTH),
		12044 => to_signed(29971, LUT_AMPL_WIDTH),
		12045 => to_signed(29972, LUT_AMPL_WIDTH),
		12046 => to_signed(29974, LUT_AMPL_WIDTH),
		12047 => to_signed(29975, LUT_AMPL_WIDTH),
		12048 => to_signed(29976, LUT_AMPL_WIDTH),
		12049 => to_signed(29978, LUT_AMPL_WIDTH),
		12050 => to_signed(29979, LUT_AMPL_WIDTH),
		12051 => to_signed(29980, LUT_AMPL_WIDTH),
		12052 => to_signed(29981, LUT_AMPL_WIDTH),
		12053 => to_signed(29983, LUT_AMPL_WIDTH),
		12054 => to_signed(29984, LUT_AMPL_WIDTH),
		12055 => to_signed(29985, LUT_AMPL_WIDTH),
		12056 => to_signed(29986, LUT_AMPL_WIDTH),
		12057 => to_signed(29988, LUT_AMPL_WIDTH),
		12058 => to_signed(29989, LUT_AMPL_WIDTH),
		12059 => to_signed(29990, LUT_AMPL_WIDTH),
		12060 => to_signed(29991, LUT_AMPL_WIDTH),
		12061 => to_signed(29993, LUT_AMPL_WIDTH),
		12062 => to_signed(29994, LUT_AMPL_WIDTH),
		12063 => to_signed(29995, LUT_AMPL_WIDTH),
		12064 => to_signed(29997, LUT_AMPL_WIDTH),
		12065 => to_signed(29998, LUT_AMPL_WIDTH),
		12066 => to_signed(29999, LUT_AMPL_WIDTH),
		12067 => to_signed(30000, LUT_AMPL_WIDTH),
		12068 => to_signed(30002, LUT_AMPL_WIDTH),
		12069 => to_signed(30003, LUT_AMPL_WIDTH),
		12070 => to_signed(30004, LUT_AMPL_WIDTH),
		12071 => to_signed(30005, LUT_AMPL_WIDTH),
		12072 => to_signed(30007, LUT_AMPL_WIDTH),
		12073 => to_signed(30008, LUT_AMPL_WIDTH),
		12074 => to_signed(30009, LUT_AMPL_WIDTH),
		12075 => to_signed(30010, LUT_AMPL_WIDTH),
		12076 => to_signed(30012, LUT_AMPL_WIDTH),
		12077 => to_signed(30013, LUT_AMPL_WIDTH),
		12078 => to_signed(30014, LUT_AMPL_WIDTH),
		12079 => to_signed(30015, LUT_AMPL_WIDTH),
		12080 => to_signed(30017, LUT_AMPL_WIDTH),
		12081 => to_signed(30018, LUT_AMPL_WIDTH),
		12082 => to_signed(30019, LUT_AMPL_WIDTH),
		12083 => to_signed(30020, LUT_AMPL_WIDTH),
		12084 => to_signed(30022, LUT_AMPL_WIDTH),
		12085 => to_signed(30023, LUT_AMPL_WIDTH),
		12086 => to_signed(30024, LUT_AMPL_WIDTH),
		12087 => to_signed(30026, LUT_AMPL_WIDTH),
		12088 => to_signed(30027, LUT_AMPL_WIDTH),
		12089 => to_signed(30028, LUT_AMPL_WIDTH),
		12090 => to_signed(30029, LUT_AMPL_WIDTH),
		12091 => to_signed(30031, LUT_AMPL_WIDTH),
		12092 => to_signed(30032, LUT_AMPL_WIDTH),
		12093 => to_signed(30033, LUT_AMPL_WIDTH),
		12094 => to_signed(30034, LUT_AMPL_WIDTH),
		12095 => to_signed(30036, LUT_AMPL_WIDTH),
		12096 => to_signed(30037, LUT_AMPL_WIDTH),
		12097 => to_signed(30038, LUT_AMPL_WIDTH),
		12098 => to_signed(30039, LUT_AMPL_WIDTH),
		12099 => to_signed(30041, LUT_AMPL_WIDTH),
		12100 => to_signed(30042, LUT_AMPL_WIDTH),
		12101 => to_signed(30043, LUT_AMPL_WIDTH),
		12102 => to_signed(30044, LUT_AMPL_WIDTH),
		12103 => to_signed(30046, LUT_AMPL_WIDTH),
		12104 => to_signed(30047, LUT_AMPL_WIDTH),
		12105 => to_signed(30048, LUT_AMPL_WIDTH),
		12106 => to_signed(30049, LUT_AMPL_WIDTH),
		12107 => to_signed(30051, LUT_AMPL_WIDTH),
		12108 => to_signed(30052, LUT_AMPL_WIDTH),
		12109 => to_signed(30053, LUT_AMPL_WIDTH),
		12110 => to_signed(30054, LUT_AMPL_WIDTH),
		12111 => to_signed(30056, LUT_AMPL_WIDTH),
		12112 => to_signed(30057, LUT_AMPL_WIDTH),
		12113 => to_signed(30058, LUT_AMPL_WIDTH),
		12114 => to_signed(30059, LUT_AMPL_WIDTH),
		12115 => to_signed(30061, LUT_AMPL_WIDTH),
		12116 => to_signed(30062, LUT_AMPL_WIDTH),
		12117 => to_signed(30063, LUT_AMPL_WIDTH),
		12118 => to_signed(30064, LUT_AMPL_WIDTH),
		12119 => to_signed(30066, LUT_AMPL_WIDTH),
		12120 => to_signed(30067, LUT_AMPL_WIDTH),
		12121 => to_signed(30068, LUT_AMPL_WIDTH),
		12122 => to_signed(30069, LUT_AMPL_WIDTH),
		12123 => to_signed(30071, LUT_AMPL_WIDTH),
		12124 => to_signed(30072, LUT_AMPL_WIDTH),
		12125 => to_signed(30073, LUT_AMPL_WIDTH),
		12126 => to_signed(30074, LUT_AMPL_WIDTH),
		12127 => to_signed(30076, LUT_AMPL_WIDTH),
		12128 => to_signed(30077, LUT_AMPL_WIDTH),
		12129 => to_signed(30078, LUT_AMPL_WIDTH),
		12130 => to_signed(30079, LUT_AMPL_WIDTH),
		12131 => to_signed(30081, LUT_AMPL_WIDTH),
		12132 => to_signed(30082, LUT_AMPL_WIDTH),
		12133 => to_signed(30083, LUT_AMPL_WIDTH),
		12134 => to_signed(30084, LUT_AMPL_WIDTH),
		12135 => to_signed(30086, LUT_AMPL_WIDTH),
		12136 => to_signed(30087, LUT_AMPL_WIDTH),
		12137 => to_signed(30088, LUT_AMPL_WIDTH),
		12138 => to_signed(30089, LUT_AMPL_WIDTH),
		12139 => to_signed(30091, LUT_AMPL_WIDTH),
		12140 => to_signed(30092, LUT_AMPL_WIDTH),
		12141 => to_signed(30093, LUT_AMPL_WIDTH),
		12142 => to_signed(30094, LUT_AMPL_WIDTH),
		12143 => to_signed(30096, LUT_AMPL_WIDTH),
		12144 => to_signed(30097, LUT_AMPL_WIDTH),
		12145 => to_signed(30098, LUT_AMPL_WIDTH),
		12146 => to_signed(30099, LUT_AMPL_WIDTH),
		12147 => to_signed(30100, LUT_AMPL_WIDTH),
		12148 => to_signed(30102, LUT_AMPL_WIDTH),
		12149 => to_signed(30103, LUT_AMPL_WIDTH),
		12150 => to_signed(30104, LUT_AMPL_WIDTH),
		12151 => to_signed(30105, LUT_AMPL_WIDTH),
		12152 => to_signed(30107, LUT_AMPL_WIDTH),
		12153 => to_signed(30108, LUT_AMPL_WIDTH),
		12154 => to_signed(30109, LUT_AMPL_WIDTH),
		12155 => to_signed(30110, LUT_AMPL_WIDTH),
		12156 => to_signed(30112, LUT_AMPL_WIDTH),
		12157 => to_signed(30113, LUT_AMPL_WIDTH),
		12158 => to_signed(30114, LUT_AMPL_WIDTH),
		12159 => to_signed(30115, LUT_AMPL_WIDTH),
		12160 => to_signed(30117, LUT_AMPL_WIDTH),
		12161 => to_signed(30118, LUT_AMPL_WIDTH),
		12162 => to_signed(30119, LUT_AMPL_WIDTH),
		12163 => to_signed(30120, LUT_AMPL_WIDTH),
		12164 => to_signed(30122, LUT_AMPL_WIDTH),
		12165 => to_signed(30123, LUT_AMPL_WIDTH),
		12166 => to_signed(30124, LUT_AMPL_WIDTH),
		12167 => to_signed(30125, LUT_AMPL_WIDTH),
		12168 => to_signed(30126, LUT_AMPL_WIDTH),
		12169 => to_signed(30128, LUT_AMPL_WIDTH),
		12170 => to_signed(30129, LUT_AMPL_WIDTH),
		12171 => to_signed(30130, LUT_AMPL_WIDTH),
		12172 => to_signed(30131, LUT_AMPL_WIDTH),
		12173 => to_signed(30133, LUT_AMPL_WIDTH),
		12174 => to_signed(30134, LUT_AMPL_WIDTH),
		12175 => to_signed(30135, LUT_AMPL_WIDTH),
		12176 => to_signed(30136, LUT_AMPL_WIDTH),
		12177 => to_signed(30138, LUT_AMPL_WIDTH),
		12178 => to_signed(30139, LUT_AMPL_WIDTH),
		12179 => to_signed(30140, LUT_AMPL_WIDTH),
		12180 => to_signed(30141, LUT_AMPL_WIDTH),
		12181 => to_signed(30143, LUT_AMPL_WIDTH),
		12182 => to_signed(30144, LUT_AMPL_WIDTH),
		12183 => to_signed(30145, LUT_AMPL_WIDTH),
		12184 => to_signed(30146, LUT_AMPL_WIDTH),
		12185 => to_signed(30147, LUT_AMPL_WIDTH),
		12186 => to_signed(30149, LUT_AMPL_WIDTH),
		12187 => to_signed(30150, LUT_AMPL_WIDTH),
		12188 => to_signed(30151, LUT_AMPL_WIDTH),
		12189 => to_signed(30152, LUT_AMPL_WIDTH),
		12190 => to_signed(30154, LUT_AMPL_WIDTH),
		12191 => to_signed(30155, LUT_AMPL_WIDTH),
		12192 => to_signed(30156, LUT_AMPL_WIDTH),
		12193 => to_signed(30157, LUT_AMPL_WIDTH),
		12194 => to_signed(30159, LUT_AMPL_WIDTH),
		12195 => to_signed(30160, LUT_AMPL_WIDTH),
		12196 => to_signed(30161, LUT_AMPL_WIDTH),
		12197 => to_signed(30162, LUT_AMPL_WIDTH),
		12198 => to_signed(30163, LUT_AMPL_WIDTH),
		12199 => to_signed(30165, LUT_AMPL_WIDTH),
		12200 => to_signed(30166, LUT_AMPL_WIDTH),
		12201 => to_signed(30167, LUT_AMPL_WIDTH),
		12202 => to_signed(30168, LUT_AMPL_WIDTH),
		12203 => to_signed(30170, LUT_AMPL_WIDTH),
		12204 => to_signed(30171, LUT_AMPL_WIDTH),
		12205 => to_signed(30172, LUT_AMPL_WIDTH),
		12206 => to_signed(30173, LUT_AMPL_WIDTH),
		12207 => to_signed(30174, LUT_AMPL_WIDTH),
		12208 => to_signed(30176, LUT_AMPL_WIDTH),
		12209 => to_signed(30177, LUT_AMPL_WIDTH),
		12210 => to_signed(30178, LUT_AMPL_WIDTH),
		12211 => to_signed(30179, LUT_AMPL_WIDTH),
		12212 => to_signed(30181, LUT_AMPL_WIDTH),
		12213 => to_signed(30182, LUT_AMPL_WIDTH),
		12214 => to_signed(30183, LUT_AMPL_WIDTH),
		12215 => to_signed(30184, LUT_AMPL_WIDTH),
		12216 => to_signed(30185, LUT_AMPL_WIDTH),
		12217 => to_signed(30187, LUT_AMPL_WIDTH),
		12218 => to_signed(30188, LUT_AMPL_WIDTH),
		12219 => to_signed(30189, LUT_AMPL_WIDTH),
		12220 => to_signed(30190, LUT_AMPL_WIDTH),
		12221 => to_signed(30192, LUT_AMPL_WIDTH),
		12222 => to_signed(30193, LUT_AMPL_WIDTH),
		12223 => to_signed(30194, LUT_AMPL_WIDTH),
		12224 => to_signed(30195, LUT_AMPL_WIDTH),
		12225 => to_signed(30196, LUT_AMPL_WIDTH),
		12226 => to_signed(30198, LUT_AMPL_WIDTH),
		12227 => to_signed(30199, LUT_AMPL_WIDTH),
		12228 => to_signed(30200, LUT_AMPL_WIDTH),
		12229 => to_signed(30201, LUT_AMPL_WIDTH),
		12230 => to_signed(30203, LUT_AMPL_WIDTH),
		12231 => to_signed(30204, LUT_AMPL_WIDTH),
		12232 => to_signed(30205, LUT_AMPL_WIDTH),
		12233 => to_signed(30206, LUT_AMPL_WIDTH),
		12234 => to_signed(30207, LUT_AMPL_WIDTH),
		12235 => to_signed(30209, LUT_AMPL_WIDTH),
		12236 => to_signed(30210, LUT_AMPL_WIDTH),
		12237 => to_signed(30211, LUT_AMPL_WIDTH),
		12238 => to_signed(30212, LUT_AMPL_WIDTH),
		12239 => to_signed(30214, LUT_AMPL_WIDTH),
		12240 => to_signed(30215, LUT_AMPL_WIDTH),
		12241 => to_signed(30216, LUT_AMPL_WIDTH),
		12242 => to_signed(30217, LUT_AMPL_WIDTH),
		12243 => to_signed(30218, LUT_AMPL_WIDTH),
		12244 => to_signed(30220, LUT_AMPL_WIDTH),
		12245 => to_signed(30221, LUT_AMPL_WIDTH),
		12246 => to_signed(30222, LUT_AMPL_WIDTH),
		12247 => to_signed(30223, LUT_AMPL_WIDTH),
		12248 => to_signed(30224, LUT_AMPL_WIDTH),
		12249 => to_signed(30226, LUT_AMPL_WIDTH),
		12250 => to_signed(30227, LUT_AMPL_WIDTH),
		12251 => to_signed(30228, LUT_AMPL_WIDTH),
		12252 => to_signed(30229, LUT_AMPL_WIDTH),
		12253 => to_signed(30231, LUT_AMPL_WIDTH),
		12254 => to_signed(30232, LUT_AMPL_WIDTH),
		12255 => to_signed(30233, LUT_AMPL_WIDTH),
		12256 => to_signed(30234, LUT_AMPL_WIDTH),
		12257 => to_signed(30235, LUT_AMPL_WIDTH),
		12258 => to_signed(30237, LUT_AMPL_WIDTH),
		12259 => to_signed(30238, LUT_AMPL_WIDTH),
		12260 => to_signed(30239, LUT_AMPL_WIDTH),
		12261 => to_signed(30240, LUT_AMPL_WIDTH),
		12262 => to_signed(30241, LUT_AMPL_WIDTH),
		12263 => to_signed(30243, LUT_AMPL_WIDTH),
		12264 => to_signed(30244, LUT_AMPL_WIDTH),
		12265 => to_signed(30245, LUT_AMPL_WIDTH),
		12266 => to_signed(30246, LUT_AMPL_WIDTH),
		12267 => to_signed(30247, LUT_AMPL_WIDTH),
		12268 => to_signed(30249, LUT_AMPL_WIDTH),
		12269 => to_signed(30250, LUT_AMPL_WIDTH),
		12270 => to_signed(30251, LUT_AMPL_WIDTH),
		12271 => to_signed(30252, LUT_AMPL_WIDTH),
		12272 => to_signed(30253, LUT_AMPL_WIDTH),
		12273 => to_signed(30255, LUT_AMPL_WIDTH),
		12274 => to_signed(30256, LUT_AMPL_WIDTH),
		12275 => to_signed(30257, LUT_AMPL_WIDTH),
		12276 => to_signed(30258, LUT_AMPL_WIDTH),
		12277 => to_signed(30260, LUT_AMPL_WIDTH),
		12278 => to_signed(30261, LUT_AMPL_WIDTH),
		12279 => to_signed(30262, LUT_AMPL_WIDTH),
		12280 => to_signed(30263, LUT_AMPL_WIDTH),
		12281 => to_signed(30264, LUT_AMPL_WIDTH),
		12282 => to_signed(30266, LUT_AMPL_WIDTH),
		12283 => to_signed(30267, LUT_AMPL_WIDTH),
		12284 => to_signed(30268, LUT_AMPL_WIDTH),
		12285 => to_signed(30269, LUT_AMPL_WIDTH),
		12286 => to_signed(30270, LUT_AMPL_WIDTH),
		12287 => to_signed(30272, LUT_AMPL_WIDTH),
		12288 => to_signed(30273, LUT_AMPL_WIDTH),
		12289 => to_signed(30274, LUT_AMPL_WIDTH),
		12290 => to_signed(30275, LUT_AMPL_WIDTH),
		12291 => to_signed(30276, LUT_AMPL_WIDTH),
		12292 => to_signed(30278, LUT_AMPL_WIDTH),
		12293 => to_signed(30279, LUT_AMPL_WIDTH),
		12294 => to_signed(30280, LUT_AMPL_WIDTH),
		12295 => to_signed(30281, LUT_AMPL_WIDTH),
		12296 => to_signed(30282, LUT_AMPL_WIDTH),
		12297 => to_signed(30284, LUT_AMPL_WIDTH),
		12298 => to_signed(30285, LUT_AMPL_WIDTH),
		12299 => to_signed(30286, LUT_AMPL_WIDTH),
		12300 => to_signed(30287, LUT_AMPL_WIDTH),
		12301 => to_signed(30288, LUT_AMPL_WIDTH),
		12302 => to_signed(30290, LUT_AMPL_WIDTH),
		12303 => to_signed(30291, LUT_AMPL_WIDTH),
		12304 => to_signed(30292, LUT_AMPL_WIDTH),
		12305 => to_signed(30293, LUT_AMPL_WIDTH),
		12306 => to_signed(30294, LUT_AMPL_WIDTH),
		12307 => to_signed(30296, LUT_AMPL_WIDTH),
		12308 => to_signed(30297, LUT_AMPL_WIDTH),
		12309 => to_signed(30298, LUT_AMPL_WIDTH),
		12310 => to_signed(30299, LUT_AMPL_WIDTH),
		12311 => to_signed(30300, LUT_AMPL_WIDTH),
		12312 => to_signed(30302, LUT_AMPL_WIDTH),
		12313 => to_signed(30303, LUT_AMPL_WIDTH),
		12314 => to_signed(30304, LUT_AMPL_WIDTH),
		12315 => to_signed(30305, LUT_AMPL_WIDTH),
		12316 => to_signed(30306, LUT_AMPL_WIDTH),
		12317 => to_signed(30308, LUT_AMPL_WIDTH),
		12318 => to_signed(30309, LUT_AMPL_WIDTH),
		12319 => to_signed(30310, LUT_AMPL_WIDTH),
		12320 => to_signed(30311, LUT_AMPL_WIDTH),
		12321 => to_signed(30312, LUT_AMPL_WIDTH),
		12322 => to_signed(30313, LUT_AMPL_WIDTH),
		12323 => to_signed(30315, LUT_AMPL_WIDTH),
		12324 => to_signed(30316, LUT_AMPL_WIDTH),
		12325 => to_signed(30317, LUT_AMPL_WIDTH),
		12326 => to_signed(30318, LUT_AMPL_WIDTH),
		12327 => to_signed(30319, LUT_AMPL_WIDTH),
		12328 => to_signed(30321, LUT_AMPL_WIDTH),
		12329 => to_signed(30322, LUT_AMPL_WIDTH),
		12330 => to_signed(30323, LUT_AMPL_WIDTH),
		12331 => to_signed(30324, LUT_AMPL_WIDTH),
		12332 => to_signed(30325, LUT_AMPL_WIDTH),
		12333 => to_signed(30327, LUT_AMPL_WIDTH),
		12334 => to_signed(30328, LUT_AMPL_WIDTH),
		12335 => to_signed(30329, LUT_AMPL_WIDTH),
		12336 => to_signed(30330, LUT_AMPL_WIDTH),
		12337 => to_signed(30331, LUT_AMPL_WIDTH),
		12338 => to_signed(30333, LUT_AMPL_WIDTH),
		12339 => to_signed(30334, LUT_AMPL_WIDTH),
		12340 => to_signed(30335, LUT_AMPL_WIDTH),
		12341 => to_signed(30336, LUT_AMPL_WIDTH),
		12342 => to_signed(30337, LUT_AMPL_WIDTH),
		12343 => to_signed(30338, LUT_AMPL_WIDTH),
		12344 => to_signed(30340, LUT_AMPL_WIDTH),
		12345 => to_signed(30341, LUT_AMPL_WIDTH),
		12346 => to_signed(30342, LUT_AMPL_WIDTH),
		12347 => to_signed(30343, LUT_AMPL_WIDTH),
		12348 => to_signed(30344, LUT_AMPL_WIDTH),
		12349 => to_signed(30346, LUT_AMPL_WIDTH),
		12350 => to_signed(30347, LUT_AMPL_WIDTH),
		12351 => to_signed(30348, LUT_AMPL_WIDTH),
		12352 => to_signed(30349, LUT_AMPL_WIDTH),
		12353 => to_signed(30350, LUT_AMPL_WIDTH),
		12354 => to_signed(30351, LUT_AMPL_WIDTH),
		12355 => to_signed(30353, LUT_AMPL_WIDTH),
		12356 => to_signed(30354, LUT_AMPL_WIDTH),
		12357 => to_signed(30355, LUT_AMPL_WIDTH),
		12358 => to_signed(30356, LUT_AMPL_WIDTH),
		12359 => to_signed(30357, LUT_AMPL_WIDTH),
		12360 => to_signed(30359, LUT_AMPL_WIDTH),
		12361 => to_signed(30360, LUT_AMPL_WIDTH),
		12362 => to_signed(30361, LUT_AMPL_WIDTH),
		12363 => to_signed(30362, LUT_AMPL_WIDTH),
		12364 => to_signed(30363, LUT_AMPL_WIDTH),
		12365 => to_signed(30365, LUT_AMPL_WIDTH),
		12366 => to_signed(30366, LUT_AMPL_WIDTH),
		12367 => to_signed(30367, LUT_AMPL_WIDTH),
		12368 => to_signed(30368, LUT_AMPL_WIDTH),
		12369 => to_signed(30369, LUT_AMPL_WIDTH),
		12370 => to_signed(30370, LUT_AMPL_WIDTH),
		12371 => to_signed(30372, LUT_AMPL_WIDTH),
		12372 => to_signed(30373, LUT_AMPL_WIDTH),
		12373 => to_signed(30374, LUT_AMPL_WIDTH),
		12374 => to_signed(30375, LUT_AMPL_WIDTH),
		12375 => to_signed(30376, LUT_AMPL_WIDTH),
		12376 => to_signed(30377, LUT_AMPL_WIDTH),
		12377 => to_signed(30379, LUT_AMPL_WIDTH),
		12378 => to_signed(30380, LUT_AMPL_WIDTH),
		12379 => to_signed(30381, LUT_AMPL_WIDTH),
		12380 => to_signed(30382, LUT_AMPL_WIDTH),
		12381 => to_signed(30383, LUT_AMPL_WIDTH),
		12382 => to_signed(30385, LUT_AMPL_WIDTH),
		12383 => to_signed(30386, LUT_AMPL_WIDTH),
		12384 => to_signed(30387, LUT_AMPL_WIDTH),
		12385 => to_signed(30388, LUT_AMPL_WIDTH),
		12386 => to_signed(30389, LUT_AMPL_WIDTH),
		12387 => to_signed(30390, LUT_AMPL_WIDTH),
		12388 => to_signed(30392, LUT_AMPL_WIDTH),
		12389 => to_signed(30393, LUT_AMPL_WIDTH),
		12390 => to_signed(30394, LUT_AMPL_WIDTH),
		12391 => to_signed(30395, LUT_AMPL_WIDTH),
		12392 => to_signed(30396, LUT_AMPL_WIDTH),
		12393 => to_signed(30397, LUT_AMPL_WIDTH),
		12394 => to_signed(30399, LUT_AMPL_WIDTH),
		12395 => to_signed(30400, LUT_AMPL_WIDTH),
		12396 => to_signed(30401, LUT_AMPL_WIDTH),
		12397 => to_signed(30402, LUT_AMPL_WIDTH),
		12398 => to_signed(30403, LUT_AMPL_WIDTH),
		12399 => to_signed(30404, LUT_AMPL_WIDTH),
		12400 => to_signed(30406, LUT_AMPL_WIDTH),
		12401 => to_signed(30407, LUT_AMPL_WIDTH),
		12402 => to_signed(30408, LUT_AMPL_WIDTH),
		12403 => to_signed(30409, LUT_AMPL_WIDTH),
		12404 => to_signed(30410, LUT_AMPL_WIDTH),
		12405 => to_signed(30412, LUT_AMPL_WIDTH),
		12406 => to_signed(30413, LUT_AMPL_WIDTH),
		12407 => to_signed(30414, LUT_AMPL_WIDTH),
		12408 => to_signed(30415, LUT_AMPL_WIDTH),
		12409 => to_signed(30416, LUT_AMPL_WIDTH),
		12410 => to_signed(30417, LUT_AMPL_WIDTH),
		12411 => to_signed(30419, LUT_AMPL_WIDTH),
		12412 => to_signed(30420, LUT_AMPL_WIDTH),
		12413 => to_signed(30421, LUT_AMPL_WIDTH),
		12414 => to_signed(30422, LUT_AMPL_WIDTH),
		12415 => to_signed(30423, LUT_AMPL_WIDTH),
		12416 => to_signed(30424, LUT_AMPL_WIDTH),
		12417 => to_signed(30426, LUT_AMPL_WIDTH),
		12418 => to_signed(30427, LUT_AMPL_WIDTH),
		12419 => to_signed(30428, LUT_AMPL_WIDTH),
		12420 => to_signed(30429, LUT_AMPL_WIDTH),
		12421 => to_signed(30430, LUT_AMPL_WIDTH),
		12422 => to_signed(30431, LUT_AMPL_WIDTH),
		12423 => to_signed(30433, LUT_AMPL_WIDTH),
		12424 => to_signed(30434, LUT_AMPL_WIDTH),
		12425 => to_signed(30435, LUT_AMPL_WIDTH),
		12426 => to_signed(30436, LUT_AMPL_WIDTH),
		12427 => to_signed(30437, LUT_AMPL_WIDTH),
		12428 => to_signed(30438, LUT_AMPL_WIDTH),
		12429 => to_signed(30439, LUT_AMPL_WIDTH),
		12430 => to_signed(30441, LUT_AMPL_WIDTH),
		12431 => to_signed(30442, LUT_AMPL_WIDTH),
		12432 => to_signed(30443, LUT_AMPL_WIDTH),
		12433 => to_signed(30444, LUT_AMPL_WIDTH),
		12434 => to_signed(30445, LUT_AMPL_WIDTH),
		12435 => to_signed(30446, LUT_AMPL_WIDTH),
		12436 => to_signed(30448, LUT_AMPL_WIDTH),
		12437 => to_signed(30449, LUT_AMPL_WIDTH),
		12438 => to_signed(30450, LUT_AMPL_WIDTH),
		12439 => to_signed(30451, LUT_AMPL_WIDTH),
		12440 => to_signed(30452, LUT_AMPL_WIDTH),
		12441 => to_signed(30453, LUT_AMPL_WIDTH),
		12442 => to_signed(30455, LUT_AMPL_WIDTH),
		12443 => to_signed(30456, LUT_AMPL_WIDTH),
		12444 => to_signed(30457, LUT_AMPL_WIDTH),
		12445 => to_signed(30458, LUT_AMPL_WIDTH),
		12446 => to_signed(30459, LUT_AMPL_WIDTH),
		12447 => to_signed(30460, LUT_AMPL_WIDTH),
		12448 => to_signed(30462, LUT_AMPL_WIDTH),
		12449 => to_signed(30463, LUT_AMPL_WIDTH),
		12450 => to_signed(30464, LUT_AMPL_WIDTH),
		12451 => to_signed(30465, LUT_AMPL_WIDTH),
		12452 => to_signed(30466, LUT_AMPL_WIDTH),
		12453 => to_signed(30467, LUT_AMPL_WIDTH),
		12454 => to_signed(30468, LUT_AMPL_WIDTH),
		12455 => to_signed(30470, LUT_AMPL_WIDTH),
		12456 => to_signed(30471, LUT_AMPL_WIDTH),
		12457 => to_signed(30472, LUT_AMPL_WIDTH),
		12458 => to_signed(30473, LUT_AMPL_WIDTH),
		12459 => to_signed(30474, LUT_AMPL_WIDTH),
		12460 => to_signed(30475, LUT_AMPL_WIDTH),
		12461 => to_signed(30477, LUT_AMPL_WIDTH),
		12462 => to_signed(30478, LUT_AMPL_WIDTH),
		12463 => to_signed(30479, LUT_AMPL_WIDTH),
		12464 => to_signed(30480, LUT_AMPL_WIDTH),
		12465 => to_signed(30481, LUT_AMPL_WIDTH),
		12466 => to_signed(30482, LUT_AMPL_WIDTH),
		12467 => to_signed(30483, LUT_AMPL_WIDTH),
		12468 => to_signed(30485, LUT_AMPL_WIDTH),
		12469 => to_signed(30486, LUT_AMPL_WIDTH),
		12470 => to_signed(30487, LUT_AMPL_WIDTH),
		12471 => to_signed(30488, LUT_AMPL_WIDTH),
		12472 => to_signed(30489, LUT_AMPL_WIDTH),
		12473 => to_signed(30490, LUT_AMPL_WIDTH),
		12474 => to_signed(30492, LUT_AMPL_WIDTH),
		12475 => to_signed(30493, LUT_AMPL_WIDTH),
		12476 => to_signed(30494, LUT_AMPL_WIDTH),
		12477 => to_signed(30495, LUT_AMPL_WIDTH),
		12478 => to_signed(30496, LUT_AMPL_WIDTH),
		12479 => to_signed(30497, LUT_AMPL_WIDTH),
		12480 => to_signed(30498, LUT_AMPL_WIDTH),
		12481 => to_signed(30500, LUT_AMPL_WIDTH),
		12482 => to_signed(30501, LUT_AMPL_WIDTH),
		12483 => to_signed(30502, LUT_AMPL_WIDTH),
		12484 => to_signed(30503, LUT_AMPL_WIDTH),
		12485 => to_signed(30504, LUT_AMPL_WIDTH),
		12486 => to_signed(30505, LUT_AMPL_WIDTH),
		12487 => to_signed(30506, LUT_AMPL_WIDTH),
		12488 => to_signed(30508, LUT_AMPL_WIDTH),
		12489 => to_signed(30509, LUT_AMPL_WIDTH),
		12490 => to_signed(30510, LUT_AMPL_WIDTH),
		12491 => to_signed(30511, LUT_AMPL_WIDTH),
		12492 => to_signed(30512, LUT_AMPL_WIDTH),
		12493 => to_signed(30513, LUT_AMPL_WIDTH),
		12494 => to_signed(30514, LUT_AMPL_WIDTH),
		12495 => to_signed(30516, LUT_AMPL_WIDTH),
		12496 => to_signed(30517, LUT_AMPL_WIDTH),
		12497 => to_signed(30518, LUT_AMPL_WIDTH),
		12498 => to_signed(30519, LUT_AMPL_WIDTH),
		12499 => to_signed(30520, LUT_AMPL_WIDTH),
		12500 => to_signed(30521, LUT_AMPL_WIDTH),
		12501 => to_signed(30522, LUT_AMPL_WIDTH),
		12502 => to_signed(30524, LUT_AMPL_WIDTH),
		12503 => to_signed(30525, LUT_AMPL_WIDTH),
		12504 => to_signed(30526, LUT_AMPL_WIDTH),
		12505 => to_signed(30527, LUT_AMPL_WIDTH),
		12506 => to_signed(30528, LUT_AMPL_WIDTH),
		12507 => to_signed(30529, LUT_AMPL_WIDTH),
		12508 => to_signed(30530, LUT_AMPL_WIDTH),
		12509 => to_signed(30532, LUT_AMPL_WIDTH),
		12510 => to_signed(30533, LUT_AMPL_WIDTH),
		12511 => to_signed(30534, LUT_AMPL_WIDTH),
		12512 => to_signed(30535, LUT_AMPL_WIDTH),
		12513 => to_signed(30536, LUT_AMPL_WIDTH),
		12514 => to_signed(30537, LUT_AMPL_WIDTH),
		12515 => to_signed(30538, LUT_AMPL_WIDTH),
		12516 => to_signed(30540, LUT_AMPL_WIDTH),
		12517 => to_signed(30541, LUT_AMPL_WIDTH),
		12518 => to_signed(30542, LUT_AMPL_WIDTH),
		12519 => to_signed(30543, LUT_AMPL_WIDTH),
		12520 => to_signed(30544, LUT_AMPL_WIDTH),
		12521 => to_signed(30545, LUT_AMPL_WIDTH),
		12522 => to_signed(30546, LUT_AMPL_WIDTH),
		12523 => to_signed(30548, LUT_AMPL_WIDTH),
		12524 => to_signed(30549, LUT_AMPL_WIDTH),
		12525 => to_signed(30550, LUT_AMPL_WIDTH),
		12526 => to_signed(30551, LUT_AMPL_WIDTH),
		12527 => to_signed(30552, LUT_AMPL_WIDTH),
		12528 => to_signed(30553, LUT_AMPL_WIDTH),
		12529 => to_signed(30554, LUT_AMPL_WIDTH),
		12530 => to_signed(30556, LUT_AMPL_WIDTH),
		12531 => to_signed(30557, LUT_AMPL_WIDTH),
		12532 => to_signed(30558, LUT_AMPL_WIDTH),
		12533 => to_signed(30559, LUT_AMPL_WIDTH),
		12534 => to_signed(30560, LUT_AMPL_WIDTH),
		12535 => to_signed(30561, LUT_AMPL_WIDTH),
		12536 => to_signed(30562, LUT_AMPL_WIDTH),
		12537 => to_signed(30563, LUT_AMPL_WIDTH),
		12538 => to_signed(30565, LUT_AMPL_WIDTH),
		12539 => to_signed(30566, LUT_AMPL_WIDTH),
		12540 => to_signed(30567, LUT_AMPL_WIDTH),
		12541 => to_signed(30568, LUT_AMPL_WIDTH),
		12542 => to_signed(30569, LUT_AMPL_WIDTH),
		12543 => to_signed(30570, LUT_AMPL_WIDTH),
		12544 => to_signed(30571, LUT_AMPL_WIDTH),
		12545 => to_signed(30573, LUT_AMPL_WIDTH),
		12546 => to_signed(30574, LUT_AMPL_WIDTH),
		12547 => to_signed(30575, LUT_AMPL_WIDTH),
		12548 => to_signed(30576, LUT_AMPL_WIDTH),
		12549 => to_signed(30577, LUT_AMPL_WIDTH),
		12550 => to_signed(30578, LUT_AMPL_WIDTH),
		12551 => to_signed(30579, LUT_AMPL_WIDTH),
		12552 => to_signed(30580, LUT_AMPL_WIDTH),
		12553 => to_signed(30582, LUT_AMPL_WIDTH),
		12554 => to_signed(30583, LUT_AMPL_WIDTH),
		12555 => to_signed(30584, LUT_AMPL_WIDTH),
		12556 => to_signed(30585, LUT_AMPL_WIDTH),
		12557 => to_signed(30586, LUT_AMPL_WIDTH),
		12558 => to_signed(30587, LUT_AMPL_WIDTH),
		12559 => to_signed(30588, LUT_AMPL_WIDTH),
		12560 => to_signed(30589, LUT_AMPL_WIDTH),
		12561 => to_signed(30591, LUT_AMPL_WIDTH),
		12562 => to_signed(30592, LUT_AMPL_WIDTH),
		12563 => to_signed(30593, LUT_AMPL_WIDTH),
		12564 => to_signed(30594, LUT_AMPL_WIDTH),
		12565 => to_signed(30595, LUT_AMPL_WIDTH),
		12566 => to_signed(30596, LUT_AMPL_WIDTH),
		12567 => to_signed(30597, LUT_AMPL_WIDTH),
		12568 => to_signed(30598, LUT_AMPL_WIDTH),
		12569 => to_signed(30600, LUT_AMPL_WIDTH),
		12570 => to_signed(30601, LUT_AMPL_WIDTH),
		12571 => to_signed(30602, LUT_AMPL_WIDTH),
		12572 => to_signed(30603, LUT_AMPL_WIDTH),
		12573 => to_signed(30604, LUT_AMPL_WIDTH),
		12574 => to_signed(30605, LUT_AMPL_WIDTH),
		12575 => to_signed(30606, LUT_AMPL_WIDTH),
		12576 => to_signed(30607, LUT_AMPL_WIDTH),
		12577 => to_signed(30609, LUT_AMPL_WIDTH),
		12578 => to_signed(30610, LUT_AMPL_WIDTH),
		12579 => to_signed(30611, LUT_AMPL_WIDTH),
		12580 => to_signed(30612, LUT_AMPL_WIDTH),
		12581 => to_signed(30613, LUT_AMPL_WIDTH),
		12582 => to_signed(30614, LUT_AMPL_WIDTH),
		12583 => to_signed(30615, LUT_AMPL_WIDTH),
		12584 => to_signed(30616, LUT_AMPL_WIDTH),
		12585 => to_signed(30617, LUT_AMPL_WIDTH),
		12586 => to_signed(30619, LUT_AMPL_WIDTH),
		12587 => to_signed(30620, LUT_AMPL_WIDTH),
		12588 => to_signed(30621, LUT_AMPL_WIDTH),
		12589 => to_signed(30622, LUT_AMPL_WIDTH),
		12590 => to_signed(30623, LUT_AMPL_WIDTH),
		12591 => to_signed(30624, LUT_AMPL_WIDTH),
		12592 => to_signed(30625, LUT_AMPL_WIDTH),
		12593 => to_signed(30626, LUT_AMPL_WIDTH),
		12594 => to_signed(30628, LUT_AMPL_WIDTH),
		12595 => to_signed(30629, LUT_AMPL_WIDTH),
		12596 => to_signed(30630, LUT_AMPL_WIDTH),
		12597 => to_signed(30631, LUT_AMPL_WIDTH),
		12598 => to_signed(30632, LUT_AMPL_WIDTH),
		12599 => to_signed(30633, LUT_AMPL_WIDTH),
		12600 => to_signed(30634, LUT_AMPL_WIDTH),
		12601 => to_signed(30635, LUT_AMPL_WIDTH),
		12602 => to_signed(30636, LUT_AMPL_WIDTH),
		12603 => to_signed(30638, LUT_AMPL_WIDTH),
		12604 => to_signed(30639, LUT_AMPL_WIDTH),
		12605 => to_signed(30640, LUT_AMPL_WIDTH),
		12606 => to_signed(30641, LUT_AMPL_WIDTH),
		12607 => to_signed(30642, LUT_AMPL_WIDTH),
		12608 => to_signed(30643, LUT_AMPL_WIDTH),
		12609 => to_signed(30644, LUT_AMPL_WIDTH),
		12610 => to_signed(30645, LUT_AMPL_WIDTH),
		12611 => to_signed(30646, LUT_AMPL_WIDTH),
		12612 => to_signed(30648, LUT_AMPL_WIDTH),
		12613 => to_signed(30649, LUT_AMPL_WIDTH),
		12614 => to_signed(30650, LUT_AMPL_WIDTH),
		12615 => to_signed(30651, LUT_AMPL_WIDTH),
		12616 => to_signed(30652, LUT_AMPL_WIDTH),
		12617 => to_signed(30653, LUT_AMPL_WIDTH),
		12618 => to_signed(30654, LUT_AMPL_WIDTH),
		12619 => to_signed(30655, LUT_AMPL_WIDTH),
		12620 => to_signed(30656, LUT_AMPL_WIDTH),
		12621 => to_signed(30658, LUT_AMPL_WIDTH),
		12622 => to_signed(30659, LUT_AMPL_WIDTH),
		12623 => to_signed(30660, LUT_AMPL_WIDTH),
		12624 => to_signed(30661, LUT_AMPL_WIDTH),
		12625 => to_signed(30662, LUT_AMPL_WIDTH),
		12626 => to_signed(30663, LUT_AMPL_WIDTH),
		12627 => to_signed(30664, LUT_AMPL_WIDTH),
		12628 => to_signed(30665, LUT_AMPL_WIDTH),
		12629 => to_signed(30666, LUT_AMPL_WIDTH),
		12630 => to_signed(30668, LUT_AMPL_WIDTH),
		12631 => to_signed(30669, LUT_AMPL_WIDTH),
		12632 => to_signed(30670, LUT_AMPL_WIDTH),
		12633 => to_signed(30671, LUT_AMPL_WIDTH),
		12634 => to_signed(30672, LUT_AMPL_WIDTH),
		12635 => to_signed(30673, LUT_AMPL_WIDTH),
		12636 => to_signed(30674, LUT_AMPL_WIDTH),
		12637 => to_signed(30675, LUT_AMPL_WIDTH),
		12638 => to_signed(30676, LUT_AMPL_WIDTH),
		12639 => to_signed(30678, LUT_AMPL_WIDTH),
		12640 => to_signed(30679, LUT_AMPL_WIDTH),
		12641 => to_signed(30680, LUT_AMPL_WIDTH),
		12642 => to_signed(30681, LUT_AMPL_WIDTH),
		12643 => to_signed(30682, LUT_AMPL_WIDTH),
		12644 => to_signed(30683, LUT_AMPL_WIDTH),
		12645 => to_signed(30684, LUT_AMPL_WIDTH),
		12646 => to_signed(30685, LUT_AMPL_WIDTH),
		12647 => to_signed(30686, LUT_AMPL_WIDTH),
		12648 => to_signed(30687, LUT_AMPL_WIDTH),
		12649 => to_signed(30689, LUT_AMPL_WIDTH),
		12650 => to_signed(30690, LUT_AMPL_WIDTH),
		12651 => to_signed(30691, LUT_AMPL_WIDTH),
		12652 => to_signed(30692, LUT_AMPL_WIDTH),
		12653 => to_signed(30693, LUT_AMPL_WIDTH),
		12654 => to_signed(30694, LUT_AMPL_WIDTH),
		12655 => to_signed(30695, LUT_AMPL_WIDTH),
		12656 => to_signed(30696, LUT_AMPL_WIDTH),
		12657 => to_signed(30697, LUT_AMPL_WIDTH),
		12658 => to_signed(30698, LUT_AMPL_WIDTH),
		12659 => to_signed(30700, LUT_AMPL_WIDTH),
		12660 => to_signed(30701, LUT_AMPL_WIDTH),
		12661 => to_signed(30702, LUT_AMPL_WIDTH),
		12662 => to_signed(30703, LUT_AMPL_WIDTH),
		12663 => to_signed(30704, LUT_AMPL_WIDTH),
		12664 => to_signed(30705, LUT_AMPL_WIDTH),
		12665 => to_signed(30706, LUT_AMPL_WIDTH),
		12666 => to_signed(30707, LUT_AMPL_WIDTH),
		12667 => to_signed(30708, LUT_AMPL_WIDTH),
		12668 => to_signed(30709, LUT_AMPL_WIDTH),
		12669 => to_signed(30711, LUT_AMPL_WIDTH),
		12670 => to_signed(30712, LUT_AMPL_WIDTH),
		12671 => to_signed(30713, LUT_AMPL_WIDTH),
		12672 => to_signed(30714, LUT_AMPL_WIDTH),
		12673 => to_signed(30715, LUT_AMPL_WIDTH),
		12674 => to_signed(30716, LUT_AMPL_WIDTH),
		12675 => to_signed(30717, LUT_AMPL_WIDTH),
		12676 => to_signed(30718, LUT_AMPL_WIDTH),
		12677 => to_signed(30719, LUT_AMPL_WIDTH),
		12678 => to_signed(30720, LUT_AMPL_WIDTH),
		12679 => to_signed(30721, LUT_AMPL_WIDTH),
		12680 => to_signed(30723, LUT_AMPL_WIDTH),
		12681 => to_signed(30724, LUT_AMPL_WIDTH),
		12682 => to_signed(30725, LUT_AMPL_WIDTH),
		12683 => to_signed(30726, LUT_AMPL_WIDTH),
		12684 => to_signed(30727, LUT_AMPL_WIDTH),
		12685 => to_signed(30728, LUT_AMPL_WIDTH),
		12686 => to_signed(30729, LUT_AMPL_WIDTH),
		12687 => to_signed(30730, LUT_AMPL_WIDTH),
		12688 => to_signed(30731, LUT_AMPL_WIDTH),
		12689 => to_signed(30732, LUT_AMPL_WIDTH),
		12690 => to_signed(30733, LUT_AMPL_WIDTH),
		12691 => to_signed(30735, LUT_AMPL_WIDTH),
		12692 => to_signed(30736, LUT_AMPL_WIDTH),
		12693 => to_signed(30737, LUT_AMPL_WIDTH),
		12694 => to_signed(30738, LUT_AMPL_WIDTH),
		12695 => to_signed(30739, LUT_AMPL_WIDTH),
		12696 => to_signed(30740, LUT_AMPL_WIDTH),
		12697 => to_signed(30741, LUT_AMPL_WIDTH),
		12698 => to_signed(30742, LUT_AMPL_WIDTH),
		12699 => to_signed(30743, LUT_AMPL_WIDTH),
		12700 => to_signed(30744, LUT_AMPL_WIDTH),
		12701 => to_signed(30745, LUT_AMPL_WIDTH),
		12702 => to_signed(30746, LUT_AMPL_WIDTH),
		12703 => to_signed(30748, LUT_AMPL_WIDTH),
		12704 => to_signed(30749, LUT_AMPL_WIDTH),
		12705 => to_signed(30750, LUT_AMPL_WIDTH),
		12706 => to_signed(30751, LUT_AMPL_WIDTH),
		12707 => to_signed(30752, LUT_AMPL_WIDTH),
		12708 => to_signed(30753, LUT_AMPL_WIDTH),
		12709 => to_signed(30754, LUT_AMPL_WIDTH),
		12710 => to_signed(30755, LUT_AMPL_WIDTH),
		12711 => to_signed(30756, LUT_AMPL_WIDTH),
		12712 => to_signed(30757, LUT_AMPL_WIDTH),
		12713 => to_signed(30758, LUT_AMPL_WIDTH),
		12714 => to_signed(30760, LUT_AMPL_WIDTH),
		12715 => to_signed(30761, LUT_AMPL_WIDTH),
		12716 => to_signed(30762, LUT_AMPL_WIDTH),
		12717 => to_signed(30763, LUT_AMPL_WIDTH),
		12718 => to_signed(30764, LUT_AMPL_WIDTH),
		12719 => to_signed(30765, LUT_AMPL_WIDTH),
		12720 => to_signed(30766, LUT_AMPL_WIDTH),
		12721 => to_signed(30767, LUT_AMPL_WIDTH),
		12722 => to_signed(30768, LUT_AMPL_WIDTH),
		12723 => to_signed(30769, LUT_AMPL_WIDTH),
		12724 => to_signed(30770, LUT_AMPL_WIDTH),
		12725 => to_signed(30771, LUT_AMPL_WIDTH),
		12726 => to_signed(30772, LUT_AMPL_WIDTH),
		12727 => to_signed(30774, LUT_AMPL_WIDTH),
		12728 => to_signed(30775, LUT_AMPL_WIDTH),
		12729 => to_signed(30776, LUT_AMPL_WIDTH),
		12730 => to_signed(30777, LUT_AMPL_WIDTH),
		12731 => to_signed(30778, LUT_AMPL_WIDTH),
		12732 => to_signed(30779, LUT_AMPL_WIDTH),
		12733 => to_signed(30780, LUT_AMPL_WIDTH),
		12734 => to_signed(30781, LUT_AMPL_WIDTH),
		12735 => to_signed(30782, LUT_AMPL_WIDTH),
		12736 => to_signed(30783, LUT_AMPL_WIDTH),
		12737 => to_signed(30784, LUT_AMPL_WIDTH),
		12738 => to_signed(30785, LUT_AMPL_WIDTH),
		12739 => to_signed(30786, LUT_AMPL_WIDTH),
		12740 => to_signed(30788, LUT_AMPL_WIDTH),
		12741 => to_signed(30789, LUT_AMPL_WIDTH),
		12742 => to_signed(30790, LUT_AMPL_WIDTH),
		12743 => to_signed(30791, LUT_AMPL_WIDTH),
		12744 => to_signed(30792, LUT_AMPL_WIDTH),
		12745 => to_signed(30793, LUT_AMPL_WIDTH),
		12746 => to_signed(30794, LUT_AMPL_WIDTH),
		12747 => to_signed(30795, LUT_AMPL_WIDTH),
		12748 => to_signed(30796, LUT_AMPL_WIDTH),
		12749 => to_signed(30797, LUT_AMPL_WIDTH),
		12750 => to_signed(30798, LUT_AMPL_WIDTH),
		12751 => to_signed(30799, LUT_AMPL_WIDTH),
		12752 => to_signed(30800, LUT_AMPL_WIDTH),
		12753 => to_signed(30802, LUT_AMPL_WIDTH),
		12754 => to_signed(30803, LUT_AMPL_WIDTH),
		12755 => to_signed(30804, LUT_AMPL_WIDTH),
		12756 => to_signed(30805, LUT_AMPL_WIDTH),
		12757 => to_signed(30806, LUT_AMPL_WIDTH),
		12758 => to_signed(30807, LUT_AMPL_WIDTH),
		12759 => to_signed(30808, LUT_AMPL_WIDTH),
		12760 => to_signed(30809, LUT_AMPL_WIDTH),
		12761 => to_signed(30810, LUT_AMPL_WIDTH),
		12762 => to_signed(30811, LUT_AMPL_WIDTH),
		12763 => to_signed(30812, LUT_AMPL_WIDTH),
		12764 => to_signed(30813, LUT_AMPL_WIDTH),
		12765 => to_signed(30814, LUT_AMPL_WIDTH),
		12766 => to_signed(30815, LUT_AMPL_WIDTH),
		12767 => to_signed(30816, LUT_AMPL_WIDTH),
		12768 => to_signed(30818, LUT_AMPL_WIDTH),
		12769 => to_signed(30819, LUT_AMPL_WIDTH),
		12770 => to_signed(30820, LUT_AMPL_WIDTH),
		12771 => to_signed(30821, LUT_AMPL_WIDTH),
		12772 => to_signed(30822, LUT_AMPL_WIDTH),
		12773 => to_signed(30823, LUT_AMPL_WIDTH),
		12774 => to_signed(30824, LUT_AMPL_WIDTH),
		12775 => to_signed(30825, LUT_AMPL_WIDTH),
		12776 => to_signed(30826, LUT_AMPL_WIDTH),
		12777 => to_signed(30827, LUT_AMPL_WIDTH),
		12778 => to_signed(30828, LUT_AMPL_WIDTH),
		12779 => to_signed(30829, LUT_AMPL_WIDTH),
		12780 => to_signed(30830, LUT_AMPL_WIDTH),
		12781 => to_signed(30831, LUT_AMPL_WIDTH),
		12782 => to_signed(30832, LUT_AMPL_WIDTH),
		12783 => to_signed(30834, LUT_AMPL_WIDTH),
		12784 => to_signed(30835, LUT_AMPL_WIDTH),
		12785 => to_signed(30836, LUT_AMPL_WIDTH),
		12786 => to_signed(30837, LUT_AMPL_WIDTH),
		12787 => to_signed(30838, LUT_AMPL_WIDTH),
		12788 => to_signed(30839, LUT_AMPL_WIDTH),
		12789 => to_signed(30840, LUT_AMPL_WIDTH),
		12790 => to_signed(30841, LUT_AMPL_WIDTH),
		12791 => to_signed(30842, LUT_AMPL_WIDTH),
		12792 => to_signed(30843, LUT_AMPL_WIDTH),
		12793 => to_signed(30844, LUT_AMPL_WIDTH),
		12794 => to_signed(30845, LUT_AMPL_WIDTH),
		12795 => to_signed(30846, LUT_AMPL_WIDTH),
		12796 => to_signed(30847, LUT_AMPL_WIDTH),
		12797 => to_signed(30848, LUT_AMPL_WIDTH),
		12798 => to_signed(30849, LUT_AMPL_WIDTH),
		12799 => to_signed(30851, LUT_AMPL_WIDTH),
		12800 => to_signed(30852, LUT_AMPL_WIDTH),
		12801 => to_signed(30853, LUT_AMPL_WIDTH),
		12802 => to_signed(30854, LUT_AMPL_WIDTH),
		12803 => to_signed(30855, LUT_AMPL_WIDTH),
		12804 => to_signed(30856, LUT_AMPL_WIDTH),
		12805 => to_signed(30857, LUT_AMPL_WIDTH),
		12806 => to_signed(30858, LUT_AMPL_WIDTH),
		12807 => to_signed(30859, LUT_AMPL_WIDTH),
		12808 => to_signed(30860, LUT_AMPL_WIDTH),
		12809 => to_signed(30861, LUT_AMPL_WIDTH),
		12810 => to_signed(30862, LUT_AMPL_WIDTH),
		12811 => to_signed(30863, LUT_AMPL_WIDTH),
		12812 => to_signed(30864, LUT_AMPL_WIDTH),
		12813 => to_signed(30865, LUT_AMPL_WIDTH),
		12814 => to_signed(30866, LUT_AMPL_WIDTH),
		12815 => to_signed(30867, LUT_AMPL_WIDTH),
		12816 => to_signed(30868, LUT_AMPL_WIDTH),
		12817 => to_signed(30870, LUT_AMPL_WIDTH),
		12818 => to_signed(30871, LUT_AMPL_WIDTH),
		12819 => to_signed(30872, LUT_AMPL_WIDTH),
		12820 => to_signed(30873, LUT_AMPL_WIDTH),
		12821 => to_signed(30874, LUT_AMPL_WIDTH),
		12822 => to_signed(30875, LUT_AMPL_WIDTH),
		12823 => to_signed(30876, LUT_AMPL_WIDTH),
		12824 => to_signed(30877, LUT_AMPL_WIDTH),
		12825 => to_signed(30878, LUT_AMPL_WIDTH),
		12826 => to_signed(30879, LUT_AMPL_WIDTH),
		12827 => to_signed(30880, LUT_AMPL_WIDTH),
		12828 => to_signed(30881, LUT_AMPL_WIDTH),
		12829 => to_signed(30882, LUT_AMPL_WIDTH),
		12830 => to_signed(30883, LUT_AMPL_WIDTH),
		12831 => to_signed(30884, LUT_AMPL_WIDTH),
		12832 => to_signed(30885, LUT_AMPL_WIDTH),
		12833 => to_signed(30886, LUT_AMPL_WIDTH),
		12834 => to_signed(30887, LUT_AMPL_WIDTH),
		12835 => to_signed(30888, LUT_AMPL_WIDTH),
		12836 => to_signed(30889, LUT_AMPL_WIDTH),
		12837 => to_signed(30891, LUT_AMPL_WIDTH),
		12838 => to_signed(30892, LUT_AMPL_WIDTH),
		12839 => to_signed(30893, LUT_AMPL_WIDTH),
		12840 => to_signed(30894, LUT_AMPL_WIDTH),
		12841 => to_signed(30895, LUT_AMPL_WIDTH),
		12842 => to_signed(30896, LUT_AMPL_WIDTH),
		12843 => to_signed(30897, LUT_AMPL_WIDTH),
		12844 => to_signed(30898, LUT_AMPL_WIDTH),
		12845 => to_signed(30899, LUT_AMPL_WIDTH),
		12846 => to_signed(30900, LUT_AMPL_WIDTH),
		12847 => to_signed(30901, LUT_AMPL_WIDTH),
		12848 => to_signed(30902, LUT_AMPL_WIDTH),
		12849 => to_signed(30903, LUT_AMPL_WIDTH),
		12850 => to_signed(30904, LUT_AMPL_WIDTH),
		12851 => to_signed(30905, LUT_AMPL_WIDTH),
		12852 => to_signed(30906, LUT_AMPL_WIDTH),
		12853 => to_signed(30907, LUT_AMPL_WIDTH),
		12854 => to_signed(30908, LUT_AMPL_WIDTH),
		12855 => to_signed(30909, LUT_AMPL_WIDTH),
		12856 => to_signed(30910, LUT_AMPL_WIDTH),
		12857 => to_signed(30911, LUT_AMPL_WIDTH),
		12858 => to_signed(30912, LUT_AMPL_WIDTH),
		12859 => to_signed(30914, LUT_AMPL_WIDTH),
		12860 => to_signed(30915, LUT_AMPL_WIDTH),
		12861 => to_signed(30916, LUT_AMPL_WIDTH),
		12862 => to_signed(30917, LUT_AMPL_WIDTH),
		12863 => to_signed(30918, LUT_AMPL_WIDTH),
		12864 => to_signed(30919, LUT_AMPL_WIDTH),
		12865 => to_signed(30920, LUT_AMPL_WIDTH),
		12866 => to_signed(30921, LUT_AMPL_WIDTH),
		12867 => to_signed(30922, LUT_AMPL_WIDTH),
		12868 => to_signed(30923, LUT_AMPL_WIDTH),
		12869 => to_signed(30924, LUT_AMPL_WIDTH),
		12870 => to_signed(30925, LUT_AMPL_WIDTH),
		12871 => to_signed(30926, LUT_AMPL_WIDTH),
		12872 => to_signed(30927, LUT_AMPL_WIDTH),
		12873 => to_signed(30928, LUT_AMPL_WIDTH),
		12874 => to_signed(30929, LUT_AMPL_WIDTH),
		12875 => to_signed(30930, LUT_AMPL_WIDTH),
		12876 => to_signed(30931, LUT_AMPL_WIDTH),
		12877 => to_signed(30932, LUT_AMPL_WIDTH),
		12878 => to_signed(30933, LUT_AMPL_WIDTH),
		12879 => to_signed(30934, LUT_AMPL_WIDTH),
		12880 => to_signed(30935, LUT_AMPL_WIDTH),
		12881 => to_signed(30936, LUT_AMPL_WIDTH),
		12882 => to_signed(30937, LUT_AMPL_WIDTH),
		12883 => to_signed(30938, LUT_AMPL_WIDTH),
		12884 => to_signed(30939, LUT_AMPL_WIDTH),
		12885 => to_signed(30941, LUT_AMPL_WIDTH),
		12886 => to_signed(30942, LUT_AMPL_WIDTH),
		12887 => to_signed(30943, LUT_AMPL_WIDTH),
		12888 => to_signed(30944, LUT_AMPL_WIDTH),
		12889 => to_signed(30945, LUT_AMPL_WIDTH),
		12890 => to_signed(30946, LUT_AMPL_WIDTH),
		12891 => to_signed(30947, LUT_AMPL_WIDTH),
		12892 => to_signed(30948, LUT_AMPL_WIDTH),
		12893 => to_signed(30949, LUT_AMPL_WIDTH),
		12894 => to_signed(30950, LUT_AMPL_WIDTH),
		12895 => to_signed(30951, LUT_AMPL_WIDTH),
		12896 => to_signed(30952, LUT_AMPL_WIDTH),
		12897 => to_signed(30953, LUT_AMPL_WIDTH),
		12898 => to_signed(30954, LUT_AMPL_WIDTH),
		12899 => to_signed(30955, LUT_AMPL_WIDTH),
		12900 => to_signed(30956, LUT_AMPL_WIDTH),
		12901 => to_signed(30957, LUT_AMPL_WIDTH),
		12902 => to_signed(30958, LUT_AMPL_WIDTH),
		12903 => to_signed(30959, LUT_AMPL_WIDTH),
		12904 => to_signed(30960, LUT_AMPL_WIDTH),
		12905 => to_signed(30961, LUT_AMPL_WIDTH),
		12906 => to_signed(30962, LUT_AMPL_WIDTH),
		12907 => to_signed(30963, LUT_AMPL_WIDTH),
		12908 => to_signed(30964, LUT_AMPL_WIDTH),
		12909 => to_signed(30965, LUT_AMPL_WIDTH),
		12910 => to_signed(30966, LUT_AMPL_WIDTH),
		12911 => to_signed(30967, LUT_AMPL_WIDTH),
		12912 => to_signed(30968, LUT_AMPL_WIDTH),
		12913 => to_signed(30969, LUT_AMPL_WIDTH),
		12914 => to_signed(30970, LUT_AMPL_WIDTH),
		12915 => to_signed(30971, LUT_AMPL_WIDTH),
		12916 => to_signed(30972, LUT_AMPL_WIDTH),
		12917 => to_signed(30973, LUT_AMPL_WIDTH),
		12918 => to_signed(30974, LUT_AMPL_WIDTH),
		12919 => to_signed(30976, LUT_AMPL_WIDTH),
		12920 => to_signed(30977, LUT_AMPL_WIDTH),
		12921 => to_signed(30978, LUT_AMPL_WIDTH),
		12922 => to_signed(30979, LUT_AMPL_WIDTH),
		12923 => to_signed(30980, LUT_AMPL_WIDTH),
		12924 => to_signed(30981, LUT_AMPL_WIDTH),
		12925 => to_signed(30982, LUT_AMPL_WIDTH),
		12926 => to_signed(30983, LUT_AMPL_WIDTH),
		12927 => to_signed(30984, LUT_AMPL_WIDTH),
		12928 => to_signed(30985, LUT_AMPL_WIDTH),
		12929 => to_signed(30986, LUT_AMPL_WIDTH),
		12930 => to_signed(30987, LUT_AMPL_WIDTH),
		12931 => to_signed(30988, LUT_AMPL_WIDTH),
		12932 => to_signed(30989, LUT_AMPL_WIDTH),
		12933 => to_signed(30990, LUT_AMPL_WIDTH),
		12934 => to_signed(30991, LUT_AMPL_WIDTH),
		12935 => to_signed(30992, LUT_AMPL_WIDTH),
		12936 => to_signed(30993, LUT_AMPL_WIDTH),
		12937 => to_signed(30994, LUT_AMPL_WIDTH),
		12938 => to_signed(30995, LUT_AMPL_WIDTH),
		12939 => to_signed(30996, LUT_AMPL_WIDTH),
		12940 => to_signed(30997, LUT_AMPL_WIDTH),
		12941 => to_signed(30998, LUT_AMPL_WIDTH),
		12942 => to_signed(30999, LUT_AMPL_WIDTH),
		12943 => to_signed(31000, LUT_AMPL_WIDTH),
		12944 => to_signed(31001, LUT_AMPL_WIDTH),
		12945 => to_signed(31002, LUT_AMPL_WIDTH),
		12946 => to_signed(31003, LUT_AMPL_WIDTH),
		12947 => to_signed(31004, LUT_AMPL_WIDTH),
		12948 => to_signed(31005, LUT_AMPL_WIDTH),
		12949 => to_signed(31006, LUT_AMPL_WIDTH),
		12950 => to_signed(31007, LUT_AMPL_WIDTH),
		12951 => to_signed(31008, LUT_AMPL_WIDTH),
		12952 => to_signed(31009, LUT_AMPL_WIDTH),
		12953 => to_signed(31010, LUT_AMPL_WIDTH),
		12954 => to_signed(31011, LUT_AMPL_WIDTH),
		12955 => to_signed(31012, LUT_AMPL_WIDTH),
		12956 => to_signed(31013, LUT_AMPL_WIDTH),
		12957 => to_signed(31014, LUT_AMPL_WIDTH),
		12958 => to_signed(31015, LUT_AMPL_WIDTH),
		12959 => to_signed(31016, LUT_AMPL_WIDTH),
		12960 => to_signed(31017, LUT_AMPL_WIDTH),
		12961 => to_signed(31018, LUT_AMPL_WIDTH),
		12962 => to_signed(31019, LUT_AMPL_WIDTH),
		12963 => to_signed(31020, LUT_AMPL_WIDTH),
		12964 => to_signed(31021, LUT_AMPL_WIDTH),
		12965 => to_signed(31022, LUT_AMPL_WIDTH),
		12966 => to_signed(31023, LUT_AMPL_WIDTH),
		12967 => to_signed(31024, LUT_AMPL_WIDTH),
		12968 => to_signed(31025, LUT_AMPL_WIDTH),
		12969 => to_signed(31026, LUT_AMPL_WIDTH),
		12970 => to_signed(31027, LUT_AMPL_WIDTH),
		12971 => to_signed(31028, LUT_AMPL_WIDTH),
		12972 => to_signed(31029, LUT_AMPL_WIDTH),
		12973 => to_signed(31030, LUT_AMPL_WIDTH),
		12974 => to_signed(31031, LUT_AMPL_WIDTH),
		12975 => to_signed(31032, LUT_AMPL_WIDTH),
		12976 => to_signed(31033, LUT_AMPL_WIDTH),
		12977 => to_signed(31034, LUT_AMPL_WIDTH),
		12978 => to_signed(31035, LUT_AMPL_WIDTH),
		12979 => to_signed(31036, LUT_AMPL_WIDTH),
		12980 => to_signed(31037, LUT_AMPL_WIDTH),
		12981 => to_signed(31038, LUT_AMPL_WIDTH),
		12982 => to_signed(31039, LUT_AMPL_WIDTH),
		12983 => to_signed(31040, LUT_AMPL_WIDTH),
		12984 => to_signed(31041, LUT_AMPL_WIDTH),
		12985 => to_signed(31043, LUT_AMPL_WIDTH),
		12986 => to_signed(31044, LUT_AMPL_WIDTH),
		12987 => to_signed(31045, LUT_AMPL_WIDTH),
		12988 => to_signed(31046, LUT_AMPL_WIDTH),
		12989 => to_signed(31047, LUT_AMPL_WIDTH),
		12990 => to_signed(31048, LUT_AMPL_WIDTH),
		12991 => to_signed(31049, LUT_AMPL_WIDTH),
		12992 => to_signed(31050, LUT_AMPL_WIDTH),
		12993 => to_signed(31051, LUT_AMPL_WIDTH),
		12994 => to_signed(31052, LUT_AMPL_WIDTH),
		12995 => to_signed(31053, LUT_AMPL_WIDTH),
		12996 => to_signed(31054, LUT_AMPL_WIDTH),
		12997 => to_signed(31055, LUT_AMPL_WIDTH),
		12998 => to_signed(31056, LUT_AMPL_WIDTH),
		12999 => to_signed(31057, LUT_AMPL_WIDTH),
		13000 => to_signed(31058, LUT_AMPL_WIDTH),
		13001 => to_signed(31059, LUT_AMPL_WIDTH),
		13002 => to_signed(31060, LUT_AMPL_WIDTH),
		13003 => to_signed(31061, LUT_AMPL_WIDTH),
		13004 => to_signed(31062, LUT_AMPL_WIDTH),
		13005 => to_signed(31063, LUT_AMPL_WIDTH),
		13006 => to_signed(31064, LUT_AMPL_WIDTH),
		13007 => to_signed(31065, LUT_AMPL_WIDTH),
		13008 => to_signed(31066, LUT_AMPL_WIDTH),
		13009 => to_signed(31067, LUT_AMPL_WIDTH),
		13010 => to_signed(31068, LUT_AMPL_WIDTH),
		13011 => to_signed(31069, LUT_AMPL_WIDTH),
		13012 => to_signed(31070, LUT_AMPL_WIDTH),
		13013 => to_signed(31071, LUT_AMPL_WIDTH),
		13014 => to_signed(31072, LUT_AMPL_WIDTH),
		13015 => to_signed(31073, LUT_AMPL_WIDTH),
		13016 => to_signed(31074, LUT_AMPL_WIDTH),
		13017 => to_signed(31075, LUT_AMPL_WIDTH),
		13018 => to_signed(31076, LUT_AMPL_WIDTH),
		13019 => to_signed(31077, LUT_AMPL_WIDTH),
		13020 => to_signed(31078, LUT_AMPL_WIDTH),
		13021 => to_signed(31079, LUT_AMPL_WIDTH),
		13022 => to_signed(31080, LUT_AMPL_WIDTH),
		13023 => to_signed(31081, LUT_AMPL_WIDTH),
		13024 => to_signed(31082, LUT_AMPL_WIDTH),
		13025 => to_signed(31083, LUT_AMPL_WIDTH),
		13026 => to_signed(31083, LUT_AMPL_WIDTH),
		13027 => to_signed(31084, LUT_AMPL_WIDTH),
		13028 => to_signed(31085, LUT_AMPL_WIDTH),
		13029 => to_signed(31086, LUT_AMPL_WIDTH),
		13030 => to_signed(31087, LUT_AMPL_WIDTH),
		13031 => to_signed(31088, LUT_AMPL_WIDTH),
		13032 => to_signed(31089, LUT_AMPL_WIDTH),
		13033 => to_signed(31090, LUT_AMPL_WIDTH),
		13034 => to_signed(31091, LUT_AMPL_WIDTH),
		13035 => to_signed(31092, LUT_AMPL_WIDTH),
		13036 => to_signed(31093, LUT_AMPL_WIDTH),
		13037 => to_signed(31094, LUT_AMPL_WIDTH),
		13038 => to_signed(31095, LUT_AMPL_WIDTH),
		13039 => to_signed(31096, LUT_AMPL_WIDTH),
		13040 => to_signed(31097, LUT_AMPL_WIDTH),
		13041 => to_signed(31098, LUT_AMPL_WIDTH),
		13042 => to_signed(31099, LUT_AMPL_WIDTH),
		13043 => to_signed(31100, LUT_AMPL_WIDTH),
		13044 => to_signed(31101, LUT_AMPL_WIDTH),
		13045 => to_signed(31102, LUT_AMPL_WIDTH),
		13046 => to_signed(31103, LUT_AMPL_WIDTH),
		13047 => to_signed(31104, LUT_AMPL_WIDTH),
		13048 => to_signed(31105, LUT_AMPL_WIDTH),
		13049 => to_signed(31106, LUT_AMPL_WIDTH),
		13050 => to_signed(31107, LUT_AMPL_WIDTH),
		13051 => to_signed(31108, LUT_AMPL_WIDTH),
		13052 => to_signed(31109, LUT_AMPL_WIDTH),
		13053 => to_signed(31110, LUT_AMPL_WIDTH),
		13054 => to_signed(31111, LUT_AMPL_WIDTH),
		13055 => to_signed(31112, LUT_AMPL_WIDTH),
		13056 => to_signed(31113, LUT_AMPL_WIDTH),
		13057 => to_signed(31114, LUT_AMPL_WIDTH),
		13058 => to_signed(31115, LUT_AMPL_WIDTH),
		13059 => to_signed(31116, LUT_AMPL_WIDTH),
		13060 => to_signed(31117, LUT_AMPL_WIDTH),
		13061 => to_signed(31118, LUT_AMPL_WIDTH),
		13062 => to_signed(31119, LUT_AMPL_WIDTH),
		13063 => to_signed(31120, LUT_AMPL_WIDTH),
		13064 => to_signed(31121, LUT_AMPL_WIDTH),
		13065 => to_signed(31122, LUT_AMPL_WIDTH),
		13066 => to_signed(31123, LUT_AMPL_WIDTH),
		13067 => to_signed(31124, LUT_AMPL_WIDTH),
		13068 => to_signed(31125, LUT_AMPL_WIDTH),
		13069 => to_signed(31126, LUT_AMPL_WIDTH),
		13070 => to_signed(31127, LUT_AMPL_WIDTH),
		13071 => to_signed(31128, LUT_AMPL_WIDTH),
		13072 => to_signed(31129, LUT_AMPL_WIDTH),
		13073 => to_signed(31130, LUT_AMPL_WIDTH),
		13074 => to_signed(31131, LUT_AMPL_WIDTH),
		13075 => to_signed(31132, LUT_AMPL_WIDTH),
		13076 => to_signed(31133, LUT_AMPL_WIDTH),
		13077 => to_signed(31134, LUT_AMPL_WIDTH),
		13078 => to_signed(31135, LUT_AMPL_WIDTH),
		13079 => to_signed(31136, LUT_AMPL_WIDTH),
		13080 => to_signed(31137, LUT_AMPL_WIDTH),
		13081 => to_signed(31138, LUT_AMPL_WIDTH),
		13082 => to_signed(31139, LUT_AMPL_WIDTH),
		13083 => to_signed(31140, LUT_AMPL_WIDTH),
		13084 => to_signed(31141, LUT_AMPL_WIDTH),
		13085 => to_signed(31142, LUT_AMPL_WIDTH),
		13086 => to_signed(31143, LUT_AMPL_WIDTH),
		13087 => to_signed(31144, LUT_AMPL_WIDTH),
		13088 => to_signed(31145, LUT_AMPL_WIDTH),
		13089 => to_signed(31146, LUT_AMPL_WIDTH),
		13090 => to_signed(31147, LUT_AMPL_WIDTH),
		13091 => to_signed(31148, LUT_AMPL_WIDTH),
		13092 => to_signed(31148, LUT_AMPL_WIDTH),
		13093 => to_signed(31149, LUT_AMPL_WIDTH),
		13094 => to_signed(31150, LUT_AMPL_WIDTH),
		13095 => to_signed(31151, LUT_AMPL_WIDTH),
		13096 => to_signed(31152, LUT_AMPL_WIDTH),
		13097 => to_signed(31153, LUT_AMPL_WIDTH),
		13098 => to_signed(31154, LUT_AMPL_WIDTH),
		13099 => to_signed(31155, LUT_AMPL_WIDTH),
		13100 => to_signed(31156, LUT_AMPL_WIDTH),
		13101 => to_signed(31157, LUT_AMPL_WIDTH),
		13102 => to_signed(31158, LUT_AMPL_WIDTH),
		13103 => to_signed(31159, LUT_AMPL_WIDTH),
		13104 => to_signed(31160, LUT_AMPL_WIDTH),
		13105 => to_signed(31161, LUT_AMPL_WIDTH),
		13106 => to_signed(31162, LUT_AMPL_WIDTH),
		13107 => to_signed(31163, LUT_AMPL_WIDTH),
		13108 => to_signed(31164, LUT_AMPL_WIDTH),
		13109 => to_signed(31165, LUT_AMPL_WIDTH),
		13110 => to_signed(31166, LUT_AMPL_WIDTH),
		13111 => to_signed(31167, LUT_AMPL_WIDTH),
		13112 => to_signed(31168, LUT_AMPL_WIDTH),
		13113 => to_signed(31169, LUT_AMPL_WIDTH),
		13114 => to_signed(31170, LUT_AMPL_WIDTH),
		13115 => to_signed(31171, LUT_AMPL_WIDTH),
		13116 => to_signed(31172, LUT_AMPL_WIDTH),
		13117 => to_signed(31173, LUT_AMPL_WIDTH),
		13118 => to_signed(31174, LUT_AMPL_WIDTH),
		13119 => to_signed(31175, LUT_AMPL_WIDTH),
		13120 => to_signed(31176, LUT_AMPL_WIDTH),
		13121 => to_signed(31177, LUT_AMPL_WIDTH),
		13122 => to_signed(31178, LUT_AMPL_WIDTH),
		13123 => to_signed(31179, LUT_AMPL_WIDTH),
		13124 => to_signed(31180, LUT_AMPL_WIDTH),
		13125 => to_signed(31181, LUT_AMPL_WIDTH),
		13126 => to_signed(31181, LUT_AMPL_WIDTH),
		13127 => to_signed(31182, LUT_AMPL_WIDTH),
		13128 => to_signed(31183, LUT_AMPL_WIDTH),
		13129 => to_signed(31184, LUT_AMPL_WIDTH),
		13130 => to_signed(31185, LUT_AMPL_WIDTH),
		13131 => to_signed(31186, LUT_AMPL_WIDTH),
		13132 => to_signed(31187, LUT_AMPL_WIDTH),
		13133 => to_signed(31188, LUT_AMPL_WIDTH),
		13134 => to_signed(31189, LUT_AMPL_WIDTH),
		13135 => to_signed(31190, LUT_AMPL_WIDTH),
		13136 => to_signed(31191, LUT_AMPL_WIDTH),
		13137 => to_signed(31192, LUT_AMPL_WIDTH),
		13138 => to_signed(31193, LUT_AMPL_WIDTH),
		13139 => to_signed(31194, LUT_AMPL_WIDTH),
		13140 => to_signed(31195, LUT_AMPL_WIDTH),
		13141 => to_signed(31196, LUT_AMPL_WIDTH),
		13142 => to_signed(31197, LUT_AMPL_WIDTH),
		13143 => to_signed(31198, LUT_AMPL_WIDTH),
		13144 => to_signed(31199, LUT_AMPL_WIDTH),
		13145 => to_signed(31200, LUT_AMPL_WIDTH),
		13146 => to_signed(31201, LUT_AMPL_WIDTH),
		13147 => to_signed(31202, LUT_AMPL_WIDTH),
		13148 => to_signed(31203, LUT_AMPL_WIDTH),
		13149 => to_signed(31204, LUT_AMPL_WIDTH),
		13150 => to_signed(31205, LUT_AMPL_WIDTH),
		13151 => to_signed(31206, LUT_AMPL_WIDTH),
		13152 => to_signed(31206, LUT_AMPL_WIDTH),
		13153 => to_signed(31207, LUT_AMPL_WIDTH),
		13154 => to_signed(31208, LUT_AMPL_WIDTH),
		13155 => to_signed(31209, LUT_AMPL_WIDTH),
		13156 => to_signed(31210, LUT_AMPL_WIDTH),
		13157 => to_signed(31211, LUT_AMPL_WIDTH),
		13158 => to_signed(31212, LUT_AMPL_WIDTH),
		13159 => to_signed(31213, LUT_AMPL_WIDTH),
		13160 => to_signed(31214, LUT_AMPL_WIDTH),
		13161 => to_signed(31215, LUT_AMPL_WIDTH),
		13162 => to_signed(31216, LUT_AMPL_WIDTH),
		13163 => to_signed(31217, LUT_AMPL_WIDTH),
		13164 => to_signed(31218, LUT_AMPL_WIDTH),
		13165 => to_signed(31219, LUT_AMPL_WIDTH),
		13166 => to_signed(31220, LUT_AMPL_WIDTH),
		13167 => to_signed(31221, LUT_AMPL_WIDTH),
		13168 => to_signed(31222, LUT_AMPL_WIDTH),
		13169 => to_signed(31223, LUT_AMPL_WIDTH),
		13170 => to_signed(31224, LUT_AMPL_WIDTH),
		13171 => to_signed(31225, LUT_AMPL_WIDTH),
		13172 => to_signed(31226, LUT_AMPL_WIDTH),
		13173 => to_signed(31227, LUT_AMPL_WIDTH),
		13174 => to_signed(31227, LUT_AMPL_WIDTH),
		13175 => to_signed(31228, LUT_AMPL_WIDTH),
		13176 => to_signed(31229, LUT_AMPL_WIDTH),
		13177 => to_signed(31230, LUT_AMPL_WIDTH),
		13178 => to_signed(31231, LUT_AMPL_WIDTH),
		13179 => to_signed(31232, LUT_AMPL_WIDTH),
		13180 => to_signed(31233, LUT_AMPL_WIDTH),
		13181 => to_signed(31234, LUT_AMPL_WIDTH),
		13182 => to_signed(31235, LUT_AMPL_WIDTH),
		13183 => to_signed(31236, LUT_AMPL_WIDTH),
		13184 => to_signed(31237, LUT_AMPL_WIDTH),
		13185 => to_signed(31238, LUT_AMPL_WIDTH),
		13186 => to_signed(31239, LUT_AMPL_WIDTH),
		13187 => to_signed(31240, LUT_AMPL_WIDTH),
		13188 => to_signed(31241, LUT_AMPL_WIDTH),
		13189 => to_signed(31242, LUT_AMPL_WIDTH),
		13190 => to_signed(31243, LUT_AMPL_WIDTH),
		13191 => to_signed(31244, LUT_AMPL_WIDTH),
		13192 => to_signed(31245, LUT_AMPL_WIDTH),
		13193 => to_signed(31246, LUT_AMPL_WIDTH),
		13194 => to_signed(31246, LUT_AMPL_WIDTH),
		13195 => to_signed(31247, LUT_AMPL_WIDTH),
		13196 => to_signed(31248, LUT_AMPL_WIDTH),
		13197 => to_signed(31249, LUT_AMPL_WIDTH),
		13198 => to_signed(31250, LUT_AMPL_WIDTH),
		13199 => to_signed(31251, LUT_AMPL_WIDTH),
		13200 => to_signed(31252, LUT_AMPL_WIDTH),
		13201 => to_signed(31253, LUT_AMPL_WIDTH),
		13202 => to_signed(31254, LUT_AMPL_WIDTH),
		13203 => to_signed(31255, LUT_AMPL_WIDTH),
		13204 => to_signed(31256, LUT_AMPL_WIDTH),
		13205 => to_signed(31257, LUT_AMPL_WIDTH),
		13206 => to_signed(31258, LUT_AMPL_WIDTH),
		13207 => to_signed(31259, LUT_AMPL_WIDTH),
		13208 => to_signed(31260, LUT_AMPL_WIDTH),
		13209 => to_signed(31261, LUT_AMPL_WIDTH),
		13210 => to_signed(31262, LUT_AMPL_WIDTH),
		13211 => to_signed(31262, LUT_AMPL_WIDTH),
		13212 => to_signed(31263, LUT_AMPL_WIDTH),
		13213 => to_signed(31264, LUT_AMPL_WIDTH),
		13214 => to_signed(31265, LUT_AMPL_WIDTH),
		13215 => to_signed(31266, LUT_AMPL_WIDTH),
		13216 => to_signed(31267, LUT_AMPL_WIDTH),
		13217 => to_signed(31268, LUT_AMPL_WIDTH),
		13218 => to_signed(31269, LUT_AMPL_WIDTH),
		13219 => to_signed(31270, LUT_AMPL_WIDTH),
		13220 => to_signed(31271, LUT_AMPL_WIDTH),
		13221 => to_signed(31272, LUT_AMPL_WIDTH),
		13222 => to_signed(31273, LUT_AMPL_WIDTH),
		13223 => to_signed(31274, LUT_AMPL_WIDTH),
		13224 => to_signed(31275, LUT_AMPL_WIDTH),
		13225 => to_signed(31276, LUT_AMPL_WIDTH),
		13226 => to_signed(31277, LUT_AMPL_WIDTH),
		13227 => to_signed(31278, LUT_AMPL_WIDTH),
		13228 => to_signed(31278, LUT_AMPL_WIDTH),
		13229 => to_signed(31279, LUT_AMPL_WIDTH),
		13230 => to_signed(31280, LUT_AMPL_WIDTH),
		13231 => to_signed(31281, LUT_AMPL_WIDTH),
		13232 => to_signed(31282, LUT_AMPL_WIDTH),
		13233 => to_signed(31283, LUT_AMPL_WIDTH),
		13234 => to_signed(31284, LUT_AMPL_WIDTH),
		13235 => to_signed(31285, LUT_AMPL_WIDTH),
		13236 => to_signed(31286, LUT_AMPL_WIDTH),
		13237 => to_signed(31287, LUT_AMPL_WIDTH),
		13238 => to_signed(31288, LUT_AMPL_WIDTH),
		13239 => to_signed(31289, LUT_AMPL_WIDTH),
		13240 => to_signed(31290, LUT_AMPL_WIDTH),
		13241 => to_signed(31291, LUT_AMPL_WIDTH),
		13242 => to_signed(31292, LUT_AMPL_WIDTH),
		13243 => to_signed(31292, LUT_AMPL_WIDTH),
		13244 => to_signed(31293, LUT_AMPL_WIDTH),
		13245 => to_signed(31294, LUT_AMPL_WIDTH),
		13246 => to_signed(31295, LUT_AMPL_WIDTH),
		13247 => to_signed(31296, LUT_AMPL_WIDTH),
		13248 => to_signed(31297, LUT_AMPL_WIDTH),
		13249 => to_signed(31298, LUT_AMPL_WIDTH),
		13250 => to_signed(31299, LUT_AMPL_WIDTH),
		13251 => to_signed(31300, LUT_AMPL_WIDTH),
		13252 => to_signed(31301, LUT_AMPL_WIDTH),
		13253 => to_signed(31302, LUT_AMPL_WIDTH),
		13254 => to_signed(31303, LUT_AMPL_WIDTH),
		13255 => to_signed(31304, LUT_AMPL_WIDTH),
		13256 => to_signed(31305, LUT_AMPL_WIDTH),
		13257 => to_signed(31305, LUT_AMPL_WIDTH),
		13258 => to_signed(31306, LUT_AMPL_WIDTH),
		13259 => to_signed(31307, LUT_AMPL_WIDTH),
		13260 => to_signed(31308, LUT_AMPL_WIDTH),
		13261 => to_signed(31309, LUT_AMPL_WIDTH),
		13262 => to_signed(31310, LUT_AMPL_WIDTH),
		13263 => to_signed(31311, LUT_AMPL_WIDTH),
		13264 => to_signed(31312, LUT_AMPL_WIDTH),
		13265 => to_signed(31313, LUT_AMPL_WIDTH),
		13266 => to_signed(31314, LUT_AMPL_WIDTH),
		13267 => to_signed(31315, LUT_AMPL_WIDTH),
		13268 => to_signed(31316, LUT_AMPL_WIDTH),
		13269 => to_signed(31317, LUT_AMPL_WIDTH),
		13270 => to_signed(31318, LUT_AMPL_WIDTH),
		13271 => to_signed(31318, LUT_AMPL_WIDTH),
		13272 => to_signed(31319, LUT_AMPL_WIDTH),
		13273 => to_signed(31320, LUT_AMPL_WIDTH),
		13274 => to_signed(31321, LUT_AMPL_WIDTH),
		13275 => to_signed(31322, LUT_AMPL_WIDTH),
		13276 => to_signed(31323, LUT_AMPL_WIDTH),
		13277 => to_signed(31324, LUT_AMPL_WIDTH),
		13278 => to_signed(31325, LUT_AMPL_WIDTH),
		13279 => to_signed(31326, LUT_AMPL_WIDTH),
		13280 => to_signed(31327, LUT_AMPL_WIDTH),
		13281 => to_signed(31328, LUT_AMPL_WIDTH),
		13282 => to_signed(31329, LUT_AMPL_WIDTH),
		13283 => to_signed(31329, LUT_AMPL_WIDTH),
		13284 => to_signed(31330, LUT_AMPL_WIDTH),
		13285 => to_signed(31331, LUT_AMPL_WIDTH),
		13286 => to_signed(31332, LUT_AMPL_WIDTH),
		13287 => to_signed(31333, LUT_AMPL_WIDTH),
		13288 => to_signed(31334, LUT_AMPL_WIDTH),
		13289 => to_signed(31335, LUT_AMPL_WIDTH),
		13290 => to_signed(31336, LUT_AMPL_WIDTH),
		13291 => to_signed(31337, LUT_AMPL_WIDTH),
		13292 => to_signed(31338, LUT_AMPL_WIDTH),
		13293 => to_signed(31339, LUT_AMPL_WIDTH),
		13294 => to_signed(31340, LUT_AMPL_WIDTH),
		13295 => to_signed(31341, LUT_AMPL_WIDTH),
		13296 => to_signed(31341, LUT_AMPL_WIDTH),
		13297 => to_signed(31342, LUT_AMPL_WIDTH),
		13298 => to_signed(31343, LUT_AMPL_WIDTH),
		13299 => to_signed(31344, LUT_AMPL_WIDTH),
		13300 => to_signed(31345, LUT_AMPL_WIDTH),
		13301 => to_signed(31346, LUT_AMPL_WIDTH),
		13302 => to_signed(31347, LUT_AMPL_WIDTH),
		13303 => to_signed(31348, LUT_AMPL_WIDTH),
		13304 => to_signed(31349, LUT_AMPL_WIDTH),
		13305 => to_signed(31350, LUT_AMPL_WIDTH),
		13306 => to_signed(31351, LUT_AMPL_WIDTH),
		13307 => to_signed(31352, LUT_AMPL_WIDTH),
		13308 => to_signed(31352, LUT_AMPL_WIDTH),
		13309 => to_signed(31353, LUT_AMPL_WIDTH),
		13310 => to_signed(31354, LUT_AMPL_WIDTH),
		13311 => to_signed(31355, LUT_AMPL_WIDTH),
		13312 => to_signed(31356, LUT_AMPL_WIDTH),
		13313 => to_signed(31357, LUT_AMPL_WIDTH),
		13314 => to_signed(31358, LUT_AMPL_WIDTH),
		13315 => to_signed(31359, LUT_AMPL_WIDTH),
		13316 => to_signed(31360, LUT_AMPL_WIDTH),
		13317 => to_signed(31361, LUT_AMPL_WIDTH),
		13318 => to_signed(31362, LUT_AMPL_WIDTH),
		13319 => to_signed(31362, LUT_AMPL_WIDTH),
		13320 => to_signed(31363, LUT_AMPL_WIDTH),
		13321 => to_signed(31364, LUT_AMPL_WIDTH),
		13322 => to_signed(31365, LUT_AMPL_WIDTH),
		13323 => to_signed(31366, LUT_AMPL_WIDTH),
		13324 => to_signed(31367, LUT_AMPL_WIDTH),
		13325 => to_signed(31368, LUT_AMPL_WIDTH),
		13326 => to_signed(31369, LUT_AMPL_WIDTH),
		13327 => to_signed(31370, LUT_AMPL_WIDTH),
		13328 => to_signed(31371, LUT_AMPL_WIDTH),
		13329 => to_signed(31372, LUT_AMPL_WIDTH),
		13330 => to_signed(31372, LUT_AMPL_WIDTH),
		13331 => to_signed(31373, LUT_AMPL_WIDTH),
		13332 => to_signed(31374, LUT_AMPL_WIDTH),
		13333 => to_signed(31375, LUT_AMPL_WIDTH),
		13334 => to_signed(31376, LUT_AMPL_WIDTH),
		13335 => to_signed(31377, LUT_AMPL_WIDTH),
		13336 => to_signed(31378, LUT_AMPL_WIDTH),
		13337 => to_signed(31379, LUT_AMPL_WIDTH),
		13338 => to_signed(31380, LUT_AMPL_WIDTH),
		13339 => to_signed(31381, LUT_AMPL_WIDTH),
		13340 => to_signed(31381, LUT_AMPL_WIDTH),
		13341 => to_signed(31382, LUT_AMPL_WIDTH),
		13342 => to_signed(31383, LUT_AMPL_WIDTH),
		13343 => to_signed(31384, LUT_AMPL_WIDTH),
		13344 => to_signed(31385, LUT_AMPL_WIDTH),
		13345 => to_signed(31386, LUT_AMPL_WIDTH),
		13346 => to_signed(31387, LUT_AMPL_WIDTH),
		13347 => to_signed(31388, LUT_AMPL_WIDTH),
		13348 => to_signed(31389, LUT_AMPL_WIDTH),
		13349 => to_signed(31390, LUT_AMPL_WIDTH),
		13350 => to_signed(31391, LUT_AMPL_WIDTH),
		13351 => to_signed(31391, LUT_AMPL_WIDTH),
		13352 => to_signed(31392, LUT_AMPL_WIDTH),
		13353 => to_signed(31393, LUT_AMPL_WIDTH),
		13354 => to_signed(31394, LUT_AMPL_WIDTH),
		13355 => to_signed(31395, LUT_AMPL_WIDTH),
		13356 => to_signed(31396, LUT_AMPL_WIDTH),
		13357 => to_signed(31397, LUT_AMPL_WIDTH),
		13358 => to_signed(31398, LUT_AMPL_WIDTH),
		13359 => to_signed(31399, LUT_AMPL_WIDTH),
		13360 => to_signed(31400, LUT_AMPL_WIDTH),
		13361 => to_signed(31400, LUT_AMPL_WIDTH),
		13362 => to_signed(31401, LUT_AMPL_WIDTH),
		13363 => to_signed(31402, LUT_AMPL_WIDTH),
		13364 => to_signed(31403, LUT_AMPL_WIDTH),
		13365 => to_signed(31404, LUT_AMPL_WIDTH),
		13366 => to_signed(31405, LUT_AMPL_WIDTH),
		13367 => to_signed(31406, LUT_AMPL_WIDTH),
		13368 => to_signed(31407, LUT_AMPL_WIDTH),
		13369 => to_signed(31408, LUT_AMPL_WIDTH),
		13370 => to_signed(31408, LUT_AMPL_WIDTH),
		13371 => to_signed(31409, LUT_AMPL_WIDTH),
		13372 => to_signed(31410, LUT_AMPL_WIDTH),
		13373 => to_signed(31411, LUT_AMPL_WIDTH),
		13374 => to_signed(31412, LUT_AMPL_WIDTH),
		13375 => to_signed(31413, LUT_AMPL_WIDTH),
		13376 => to_signed(31414, LUT_AMPL_WIDTH),
		13377 => to_signed(31415, LUT_AMPL_WIDTH),
		13378 => to_signed(31416, LUT_AMPL_WIDTH),
		13379 => to_signed(31417, LUT_AMPL_WIDTH),
		13380 => to_signed(31417, LUT_AMPL_WIDTH),
		13381 => to_signed(31418, LUT_AMPL_WIDTH),
		13382 => to_signed(31419, LUT_AMPL_WIDTH),
		13383 => to_signed(31420, LUT_AMPL_WIDTH),
		13384 => to_signed(31421, LUT_AMPL_WIDTH),
		13385 => to_signed(31422, LUT_AMPL_WIDTH),
		13386 => to_signed(31423, LUT_AMPL_WIDTH),
		13387 => to_signed(31424, LUT_AMPL_WIDTH),
		13388 => to_signed(31425, LUT_AMPL_WIDTH),
		13389 => to_signed(31425, LUT_AMPL_WIDTH),
		13390 => to_signed(31426, LUT_AMPL_WIDTH),
		13391 => to_signed(31427, LUT_AMPL_WIDTH),
		13392 => to_signed(31428, LUT_AMPL_WIDTH),
		13393 => to_signed(31429, LUT_AMPL_WIDTH),
		13394 => to_signed(31430, LUT_AMPL_WIDTH),
		13395 => to_signed(31431, LUT_AMPL_WIDTH),
		13396 => to_signed(31432, LUT_AMPL_WIDTH),
		13397 => to_signed(31433, LUT_AMPL_WIDTH),
		13398 => to_signed(31433, LUT_AMPL_WIDTH),
		13399 => to_signed(31434, LUT_AMPL_WIDTH),
		13400 => to_signed(31435, LUT_AMPL_WIDTH),
		13401 => to_signed(31436, LUT_AMPL_WIDTH),
		13402 => to_signed(31437, LUT_AMPL_WIDTH),
		13403 => to_signed(31438, LUT_AMPL_WIDTH),
		13404 => to_signed(31439, LUT_AMPL_WIDTH),
		13405 => to_signed(31440, LUT_AMPL_WIDTH),
		13406 => to_signed(31441, LUT_AMPL_WIDTH),
		13407 => to_signed(31441, LUT_AMPL_WIDTH),
		13408 => to_signed(31442, LUT_AMPL_WIDTH),
		13409 => to_signed(31443, LUT_AMPL_WIDTH),
		13410 => to_signed(31444, LUT_AMPL_WIDTH),
		13411 => to_signed(31445, LUT_AMPL_WIDTH),
		13412 => to_signed(31446, LUT_AMPL_WIDTH),
		13413 => to_signed(31447, LUT_AMPL_WIDTH),
		13414 => to_signed(31448, LUT_AMPL_WIDTH),
		13415 => to_signed(31448, LUT_AMPL_WIDTH),
		13416 => to_signed(31449, LUT_AMPL_WIDTH),
		13417 => to_signed(31450, LUT_AMPL_WIDTH),
		13418 => to_signed(31451, LUT_AMPL_WIDTH),
		13419 => to_signed(31452, LUT_AMPL_WIDTH),
		13420 => to_signed(31453, LUT_AMPL_WIDTH),
		13421 => to_signed(31454, LUT_AMPL_WIDTH),
		13422 => to_signed(31455, LUT_AMPL_WIDTH),
		13423 => to_signed(31456, LUT_AMPL_WIDTH),
		13424 => to_signed(31456, LUT_AMPL_WIDTH),
		13425 => to_signed(31457, LUT_AMPL_WIDTH),
		13426 => to_signed(31458, LUT_AMPL_WIDTH),
		13427 => to_signed(31459, LUT_AMPL_WIDTH),
		13428 => to_signed(31460, LUT_AMPL_WIDTH),
		13429 => to_signed(31461, LUT_AMPL_WIDTH),
		13430 => to_signed(31462, LUT_AMPL_WIDTH),
		13431 => to_signed(31463, LUT_AMPL_WIDTH),
		13432 => to_signed(31463, LUT_AMPL_WIDTH),
		13433 => to_signed(31464, LUT_AMPL_WIDTH),
		13434 => to_signed(31465, LUT_AMPL_WIDTH),
		13435 => to_signed(31466, LUT_AMPL_WIDTH),
		13436 => to_signed(31467, LUT_AMPL_WIDTH),
		13437 => to_signed(31468, LUT_AMPL_WIDTH),
		13438 => to_signed(31469, LUT_AMPL_WIDTH),
		13439 => to_signed(31470, LUT_AMPL_WIDTH),
		13440 => to_signed(31470, LUT_AMPL_WIDTH),
		13441 => to_signed(31471, LUT_AMPL_WIDTH),
		13442 => to_signed(31472, LUT_AMPL_WIDTH),
		13443 => to_signed(31473, LUT_AMPL_WIDTH),
		13444 => to_signed(31474, LUT_AMPL_WIDTH),
		13445 => to_signed(31475, LUT_AMPL_WIDTH),
		13446 => to_signed(31476, LUT_AMPL_WIDTH),
		13447 => to_signed(31477, LUT_AMPL_WIDTH),
		13448 => to_signed(31477, LUT_AMPL_WIDTH),
		13449 => to_signed(31478, LUT_AMPL_WIDTH),
		13450 => to_signed(31479, LUT_AMPL_WIDTH),
		13451 => to_signed(31480, LUT_AMPL_WIDTH),
		13452 => to_signed(31481, LUT_AMPL_WIDTH),
		13453 => to_signed(31482, LUT_AMPL_WIDTH),
		13454 => to_signed(31483, LUT_AMPL_WIDTH),
		13455 => to_signed(31484, LUT_AMPL_WIDTH),
		13456 => to_signed(31484, LUT_AMPL_WIDTH),
		13457 => to_signed(31485, LUT_AMPL_WIDTH),
		13458 => to_signed(31486, LUT_AMPL_WIDTH),
		13459 => to_signed(31487, LUT_AMPL_WIDTH),
		13460 => to_signed(31488, LUT_AMPL_WIDTH),
		13461 => to_signed(31489, LUT_AMPL_WIDTH),
		13462 => to_signed(31490, LUT_AMPL_WIDTH),
		13463 => to_signed(31490, LUT_AMPL_WIDTH),
		13464 => to_signed(31491, LUT_AMPL_WIDTH),
		13465 => to_signed(31492, LUT_AMPL_WIDTH),
		13466 => to_signed(31493, LUT_AMPL_WIDTH),
		13467 => to_signed(31494, LUT_AMPL_WIDTH),
		13468 => to_signed(31495, LUT_AMPL_WIDTH),
		13469 => to_signed(31496, LUT_AMPL_WIDTH),
		13470 => to_signed(31497, LUT_AMPL_WIDTH),
		13471 => to_signed(31497, LUT_AMPL_WIDTH),
		13472 => to_signed(31498, LUT_AMPL_WIDTH),
		13473 => to_signed(31499, LUT_AMPL_WIDTH),
		13474 => to_signed(31500, LUT_AMPL_WIDTH),
		13475 => to_signed(31501, LUT_AMPL_WIDTH),
		13476 => to_signed(31502, LUT_AMPL_WIDTH),
		13477 => to_signed(31503, LUT_AMPL_WIDTH),
		13478 => to_signed(31503, LUT_AMPL_WIDTH),
		13479 => to_signed(31504, LUT_AMPL_WIDTH),
		13480 => to_signed(31505, LUT_AMPL_WIDTH),
		13481 => to_signed(31506, LUT_AMPL_WIDTH),
		13482 => to_signed(31507, LUT_AMPL_WIDTH),
		13483 => to_signed(31508, LUT_AMPL_WIDTH),
		13484 => to_signed(31509, LUT_AMPL_WIDTH),
		13485 => to_signed(31510, LUT_AMPL_WIDTH),
		13486 => to_signed(31510, LUT_AMPL_WIDTH),
		13487 => to_signed(31511, LUT_AMPL_WIDTH),
		13488 => to_signed(31512, LUT_AMPL_WIDTH),
		13489 => to_signed(31513, LUT_AMPL_WIDTH),
		13490 => to_signed(31514, LUT_AMPL_WIDTH),
		13491 => to_signed(31515, LUT_AMPL_WIDTH),
		13492 => to_signed(31516, LUT_AMPL_WIDTH),
		13493 => to_signed(31516, LUT_AMPL_WIDTH),
		13494 => to_signed(31517, LUT_AMPL_WIDTH),
		13495 => to_signed(31518, LUT_AMPL_WIDTH),
		13496 => to_signed(31519, LUT_AMPL_WIDTH),
		13497 => to_signed(31520, LUT_AMPL_WIDTH),
		13498 => to_signed(31521, LUT_AMPL_WIDTH),
		13499 => to_signed(31522, LUT_AMPL_WIDTH),
		13500 => to_signed(31522, LUT_AMPL_WIDTH),
		13501 => to_signed(31523, LUT_AMPL_WIDTH),
		13502 => to_signed(31524, LUT_AMPL_WIDTH),
		13503 => to_signed(31525, LUT_AMPL_WIDTH),
		13504 => to_signed(31526, LUT_AMPL_WIDTH),
		13505 => to_signed(31527, LUT_AMPL_WIDTH),
		13506 => to_signed(31528, LUT_AMPL_WIDTH),
		13507 => to_signed(31528, LUT_AMPL_WIDTH),
		13508 => to_signed(31529, LUT_AMPL_WIDTH),
		13509 => to_signed(31530, LUT_AMPL_WIDTH),
		13510 => to_signed(31531, LUT_AMPL_WIDTH),
		13511 => to_signed(31532, LUT_AMPL_WIDTH),
		13512 => to_signed(31533, LUT_AMPL_WIDTH),
		13513 => to_signed(31534, LUT_AMPL_WIDTH),
		13514 => to_signed(31534, LUT_AMPL_WIDTH),
		13515 => to_signed(31535, LUT_AMPL_WIDTH),
		13516 => to_signed(31536, LUT_AMPL_WIDTH),
		13517 => to_signed(31537, LUT_AMPL_WIDTH),
		13518 => to_signed(31538, LUT_AMPL_WIDTH),
		13519 => to_signed(31539, LUT_AMPL_WIDTH),
		13520 => to_signed(31539, LUT_AMPL_WIDTH),
		13521 => to_signed(31540, LUT_AMPL_WIDTH),
		13522 => to_signed(31541, LUT_AMPL_WIDTH),
		13523 => to_signed(31542, LUT_AMPL_WIDTH),
		13524 => to_signed(31543, LUT_AMPL_WIDTH),
		13525 => to_signed(31544, LUT_AMPL_WIDTH),
		13526 => to_signed(31545, LUT_AMPL_WIDTH),
		13527 => to_signed(31545, LUT_AMPL_WIDTH),
		13528 => to_signed(31546, LUT_AMPL_WIDTH),
		13529 => to_signed(31547, LUT_AMPL_WIDTH),
		13530 => to_signed(31548, LUT_AMPL_WIDTH),
		13531 => to_signed(31549, LUT_AMPL_WIDTH),
		13532 => to_signed(31550, LUT_AMPL_WIDTH),
		13533 => to_signed(31551, LUT_AMPL_WIDTH),
		13534 => to_signed(31551, LUT_AMPL_WIDTH),
		13535 => to_signed(31552, LUT_AMPL_WIDTH),
		13536 => to_signed(31553, LUT_AMPL_WIDTH),
		13537 => to_signed(31554, LUT_AMPL_WIDTH),
		13538 => to_signed(31555, LUT_AMPL_WIDTH),
		13539 => to_signed(31556, LUT_AMPL_WIDTH),
		13540 => to_signed(31556, LUT_AMPL_WIDTH),
		13541 => to_signed(31557, LUT_AMPL_WIDTH),
		13542 => to_signed(31558, LUT_AMPL_WIDTH),
		13543 => to_signed(31559, LUT_AMPL_WIDTH),
		13544 => to_signed(31560, LUT_AMPL_WIDTH),
		13545 => to_signed(31561, LUT_AMPL_WIDTH),
		13546 => to_signed(31562, LUT_AMPL_WIDTH),
		13547 => to_signed(31562, LUT_AMPL_WIDTH),
		13548 => to_signed(31563, LUT_AMPL_WIDTH),
		13549 => to_signed(31564, LUT_AMPL_WIDTH),
		13550 => to_signed(31565, LUT_AMPL_WIDTH),
		13551 => to_signed(31566, LUT_AMPL_WIDTH),
		13552 => to_signed(31567, LUT_AMPL_WIDTH),
		13553 => to_signed(31567, LUT_AMPL_WIDTH),
		13554 => to_signed(31568, LUT_AMPL_WIDTH),
		13555 => to_signed(31569, LUT_AMPL_WIDTH),
		13556 => to_signed(31570, LUT_AMPL_WIDTH),
		13557 => to_signed(31571, LUT_AMPL_WIDTH),
		13558 => to_signed(31572, LUT_AMPL_WIDTH),
		13559 => to_signed(31572, LUT_AMPL_WIDTH),
		13560 => to_signed(31573, LUT_AMPL_WIDTH),
		13561 => to_signed(31574, LUT_AMPL_WIDTH),
		13562 => to_signed(31575, LUT_AMPL_WIDTH),
		13563 => to_signed(31576, LUT_AMPL_WIDTH),
		13564 => to_signed(31577, LUT_AMPL_WIDTH),
		13565 => to_signed(31578, LUT_AMPL_WIDTH),
		13566 => to_signed(31578, LUT_AMPL_WIDTH),
		13567 => to_signed(31579, LUT_AMPL_WIDTH),
		13568 => to_signed(31580, LUT_AMPL_WIDTH),
		13569 => to_signed(31581, LUT_AMPL_WIDTH),
		13570 => to_signed(31582, LUT_AMPL_WIDTH),
		13571 => to_signed(31583, LUT_AMPL_WIDTH),
		13572 => to_signed(31583, LUT_AMPL_WIDTH),
		13573 => to_signed(31584, LUT_AMPL_WIDTH),
		13574 => to_signed(31585, LUT_AMPL_WIDTH),
		13575 => to_signed(31586, LUT_AMPL_WIDTH),
		13576 => to_signed(31587, LUT_AMPL_WIDTH),
		13577 => to_signed(31588, LUT_AMPL_WIDTH),
		13578 => to_signed(31588, LUT_AMPL_WIDTH),
		13579 => to_signed(31589, LUT_AMPL_WIDTH),
		13580 => to_signed(31590, LUT_AMPL_WIDTH),
		13581 => to_signed(31591, LUT_AMPL_WIDTH),
		13582 => to_signed(31592, LUT_AMPL_WIDTH),
		13583 => to_signed(31593, LUT_AMPL_WIDTH),
		13584 => to_signed(31593, LUT_AMPL_WIDTH),
		13585 => to_signed(31594, LUT_AMPL_WIDTH),
		13586 => to_signed(31595, LUT_AMPL_WIDTH),
		13587 => to_signed(31596, LUT_AMPL_WIDTH),
		13588 => to_signed(31597, LUT_AMPL_WIDTH),
		13589 => to_signed(31598, LUT_AMPL_WIDTH),
		13590 => to_signed(31598, LUT_AMPL_WIDTH),
		13591 => to_signed(31599, LUT_AMPL_WIDTH),
		13592 => to_signed(31600, LUT_AMPL_WIDTH),
		13593 => to_signed(31601, LUT_AMPL_WIDTH),
		13594 => to_signed(31602, LUT_AMPL_WIDTH),
		13595 => to_signed(31603, LUT_AMPL_WIDTH),
		13596 => to_signed(31603, LUT_AMPL_WIDTH),
		13597 => to_signed(31604, LUT_AMPL_WIDTH),
		13598 => to_signed(31605, LUT_AMPL_WIDTH),
		13599 => to_signed(31606, LUT_AMPL_WIDTH),
		13600 => to_signed(31607, LUT_AMPL_WIDTH),
		13601 => to_signed(31608, LUT_AMPL_WIDTH),
		13602 => to_signed(31608, LUT_AMPL_WIDTH),
		13603 => to_signed(31609, LUT_AMPL_WIDTH),
		13604 => to_signed(31610, LUT_AMPL_WIDTH),
		13605 => to_signed(31611, LUT_AMPL_WIDTH),
		13606 => to_signed(31612, LUT_AMPL_WIDTH),
		13607 => to_signed(31613, LUT_AMPL_WIDTH),
		13608 => to_signed(31613, LUT_AMPL_WIDTH),
		13609 => to_signed(31614, LUT_AMPL_WIDTH),
		13610 => to_signed(31615, LUT_AMPL_WIDTH),
		13611 => to_signed(31616, LUT_AMPL_WIDTH),
		13612 => to_signed(31617, LUT_AMPL_WIDTH),
		13613 => to_signed(31617, LUT_AMPL_WIDTH),
		13614 => to_signed(31618, LUT_AMPL_WIDTH),
		13615 => to_signed(31619, LUT_AMPL_WIDTH),
		13616 => to_signed(31620, LUT_AMPL_WIDTH),
		13617 => to_signed(31621, LUT_AMPL_WIDTH),
		13618 => to_signed(31622, LUT_AMPL_WIDTH),
		13619 => to_signed(31622, LUT_AMPL_WIDTH),
		13620 => to_signed(31623, LUT_AMPL_WIDTH),
		13621 => to_signed(31624, LUT_AMPL_WIDTH),
		13622 => to_signed(31625, LUT_AMPL_WIDTH),
		13623 => to_signed(31626, LUT_AMPL_WIDTH),
		13624 => to_signed(31627, LUT_AMPL_WIDTH),
		13625 => to_signed(31627, LUT_AMPL_WIDTH),
		13626 => to_signed(31628, LUT_AMPL_WIDTH),
		13627 => to_signed(31629, LUT_AMPL_WIDTH),
		13628 => to_signed(31630, LUT_AMPL_WIDTH),
		13629 => to_signed(31631, LUT_AMPL_WIDTH),
		13630 => to_signed(31631, LUT_AMPL_WIDTH),
		13631 => to_signed(31632, LUT_AMPL_WIDTH),
		13632 => to_signed(31633, LUT_AMPL_WIDTH),
		13633 => to_signed(31634, LUT_AMPL_WIDTH),
		13634 => to_signed(31635, LUT_AMPL_WIDTH),
		13635 => to_signed(31636, LUT_AMPL_WIDTH),
		13636 => to_signed(31636, LUT_AMPL_WIDTH),
		13637 => to_signed(31637, LUT_AMPL_WIDTH),
		13638 => to_signed(31638, LUT_AMPL_WIDTH),
		13639 => to_signed(31639, LUT_AMPL_WIDTH),
		13640 => to_signed(31640, LUT_AMPL_WIDTH),
		13641 => to_signed(31640, LUT_AMPL_WIDTH),
		13642 => to_signed(31641, LUT_AMPL_WIDTH),
		13643 => to_signed(31642, LUT_AMPL_WIDTH),
		13644 => to_signed(31643, LUT_AMPL_WIDTH),
		13645 => to_signed(31644, LUT_AMPL_WIDTH),
		13646 => to_signed(31645, LUT_AMPL_WIDTH),
		13647 => to_signed(31645, LUT_AMPL_WIDTH),
		13648 => to_signed(31646, LUT_AMPL_WIDTH),
		13649 => to_signed(31647, LUT_AMPL_WIDTH),
		13650 => to_signed(31648, LUT_AMPL_WIDTH),
		13651 => to_signed(31649, LUT_AMPL_WIDTH),
		13652 => to_signed(31649, LUT_AMPL_WIDTH),
		13653 => to_signed(31650, LUT_AMPL_WIDTH),
		13654 => to_signed(31651, LUT_AMPL_WIDTH),
		13655 => to_signed(31652, LUT_AMPL_WIDTH),
		13656 => to_signed(31653, LUT_AMPL_WIDTH),
		13657 => to_signed(31653, LUT_AMPL_WIDTH),
		13658 => to_signed(31654, LUT_AMPL_WIDTH),
		13659 => to_signed(31655, LUT_AMPL_WIDTH),
		13660 => to_signed(31656, LUT_AMPL_WIDTH),
		13661 => to_signed(31657, LUT_AMPL_WIDTH),
		13662 => to_signed(31658, LUT_AMPL_WIDTH),
		13663 => to_signed(31658, LUT_AMPL_WIDTH),
		13664 => to_signed(31659, LUT_AMPL_WIDTH),
		13665 => to_signed(31660, LUT_AMPL_WIDTH),
		13666 => to_signed(31661, LUT_AMPL_WIDTH),
		13667 => to_signed(31662, LUT_AMPL_WIDTH),
		13668 => to_signed(31662, LUT_AMPL_WIDTH),
		13669 => to_signed(31663, LUT_AMPL_WIDTH),
		13670 => to_signed(31664, LUT_AMPL_WIDTH),
		13671 => to_signed(31665, LUT_AMPL_WIDTH),
		13672 => to_signed(31666, LUT_AMPL_WIDTH),
		13673 => to_signed(31666, LUT_AMPL_WIDTH),
		13674 => to_signed(31667, LUT_AMPL_WIDTH),
		13675 => to_signed(31668, LUT_AMPL_WIDTH),
		13676 => to_signed(31669, LUT_AMPL_WIDTH),
		13677 => to_signed(31670, LUT_AMPL_WIDTH),
		13678 => to_signed(31670, LUT_AMPL_WIDTH),
		13679 => to_signed(31671, LUT_AMPL_WIDTH),
		13680 => to_signed(31672, LUT_AMPL_WIDTH),
		13681 => to_signed(31673, LUT_AMPL_WIDTH),
		13682 => to_signed(31674, LUT_AMPL_WIDTH),
		13683 => to_signed(31674, LUT_AMPL_WIDTH),
		13684 => to_signed(31675, LUT_AMPL_WIDTH),
		13685 => to_signed(31676, LUT_AMPL_WIDTH),
		13686 => to_signed(31677, LUT_AMPL_WIDTH),
		13687 => to_signed(31678, LUT_AMPL_WIDTH),
		13688 => to_signed(31679, LUT_AMPL_WIDTH),
		13689 => to_signed(31679, LUT_AMPL_WIDTH),
		13690 => to_signed(31680, LUT_AMPL_WIDTH),
		13691 => to_signed(31681, LUT_AMPL_WIDTH),
		13692 => to_signed(31682, LUT_AMPL_WIDTH),
		13693 => to_signed(31683, LUT_AMPL_WIDTH),
		13694 => to_signed(31683, LUT_AMPL_WIDTH),
		13695 => to_signed(31684, LUT_AMPL_WIDTH),
		13696 => to_signed(31685, LUT_AMPL_WIDTH),
		13697 => to_signed(31686, LUT_AMPL_WIDTH),
		13698 => to_signed(31687, LUT_AMPL_WIDTH),
		13699 => to_signed(31687, LUT_AMPL_WIDTH),
		13700 => to_signed(31688, LUT_AMPL_WIDTH),
		13701 => to_signed(31689, LUT_AMPL_WIDTH),
		13702 => to_signed(31690, LUT_AMPL_WIDTH),
		13703 => to_signed(31691, LUT_AMPL_WIDTH),
		13704 => to_signed(31691, LUT_AMPL_WIDTH),
		13705 => to_signed(31692, LUT_AMPL_WIDTH),
		13706 => to_signed(31693, LUT_AMPL_WIDTH),
		13707 => to_signed(31694, LUT_AMPL_WIDTH),
		13708 => to_signed(31695, LUT_AMPL_WIDTH),
		13709 => to_signed(31695, LUT_AMPL_WIDTH),
		13710 => to_signed(31696, LUT_AMPL_WIDTH),
		13711 => to_signed(31697, LUT_AMPL_WIDTH),
		13712 => to_signed(31698, LUT_AMPL_WIDTH),
		13713 => to_signed(31698, LUT_AMPL_WIDTH),
		13714 => to_signed(31699, LUT_AMPL_WIDTH),
		13715 => to_signed(31700, LUT_AMPL_WIDTH),
		13716 => to_signed(31701, LUT_AMPL_WIDTH),
		13717 => to_signed(31702, LUT_AMPL_WIDTH),
		13718 => to_signed(31702, LUT_AMPL_WIDTH),
		13719 => to_signed(31703, LUT_AMPL_WIDTH),
		13720 => to_signed(31704, LUT_AMPL_WIDTH),
		13721 => to_signed(31705, LUT_AMPL_WIDTH),
		13722 => to_signed(31706, LUT_AMPL_WIDTH),
		13723 => to_signed(31706, LUT_AMPL_WIDTH),
		13724 => to_signed(31707, LUT_AMPL_WIDTH),
		13725 => to_signed(31708, LUT_AMPL_WIDTH),
		13726 => to_signed(31709, LUT_AMPL_WIDTH),
		13727 => to_signed(31710, LUT_AMPL_WIDTH),
		13728 => to_signed(31710, LUT_AMPL_WIDTH),
		13729 => to_signed(31711, LUT_AMPL_WIDTH),
		13730 => to_signed(31712, LUT_AMPL_WIDTH),
		13731 => to_signed(31713, LUT_AMPL_WIDTH),
		13732 => to_signed(31714, LUT_AMPL_WIDTH),
		13733 => to_signed(31714, LUT_AMPL_WIDTH),
		13734 => to_signed(31715, LUT_AMPL_WIDTH),
		13735 => to_signed(31716, LUT_AMPL_WIDTH),
		13736 => to_signed(31717, LUT_AMPL_WIDTH),
		13737 => to_signed(31718, LUT_AMPL_WIDTH),
		13738 => to_signed(31718, LUT_AMPL_WIDTH),
		13739 => to_signed(31719, LUT_AMPL_WIDTH),
		13740 => to_signed(31720, LUT_AMPL_WIDTH),
		13741 => to_signed(31721, LUT_AMPL_WIDTH),
		13742 => to_signed(31721, LUT_AMPL_WIDTH),
		13743 => to_signed(31722, LUT_AMPL_WIDTH),
		13744 => to_signed(31723, LUT_AMPL_WIDTH),
		13745 => to_signed(31724, LUT_AMPL_WIDTH),
		13746 => to_signed(31725, LUT_AMPL_WIDTH),
		13747 => to_signed(31725, LUT_AMPL_WIDTH),
		13748 => to_signed(31726, LUT_AMPL_WIDTH),
		13749 => to_signed(31727, LUT_AMPL_WIDTH),
		13750 => to_signed(31728, LUT_AMPL_WIDTH),
		13751 => to_signed(31729, LUT_AMPL_WIDTH),
		13752 => to_signed(31729, LUT_AMPL_WIDTH),
		13753 => to_signed(31730, LUT_AMPL_WIDTH),
		13754 => to_signed(31731, LUT_AMPL_WIDTH),
		13755 => to_signed(31732, LUT_AMPL_WIDTH),
		13756 => to_signed(31732, LUT_AMPL_WIDTH),
		13757 => to_signed(31733, LUT_AMPL_WIDTH),
		13758 => to_signed(31734, LUT_AMPL_WIDTH),
		13759 => to_signed(31735, LUT_AMPL_WIDTH),
		13760 => to_signed(31736, LUT_AMPL_WIDTH),
		13761 => to_signed(31736, LUT_AMPL_WIDTH),
		13762 => to_signed(31737, LUT_AMPL_WIDTH),
		13763 => to_signed(31738, LUT_AMPL_WIDTH),
		13764 => to_signed(31739, LUT_AMPL_WIDTH),
		13765 => to_signed(31739, LUT_AMPL_WIDTH),
		13766 => to_signed(31740, LUT_AMPL_WIDTH),
		13767 => to_signed(31741, LUT_AMPL_WIDTH),
		13768 => to_signed(31742, LUT_AMPL_WIDTH),
		13769 => to_signed(31743, LUT_AMPL_WIDTH),
		13770 => to_signed(31743, LUT_AMPL_WIDTH),
		13771 => to_signed(31744, LUT_AMPL_WIDTH),
		13772 => to_signed(31745, LUT_AMPL_WIDTH),
		13773 => to_signed(31746, LUT_AMPL_WIDTH),
		13774 => to_signed(31746, LUT_AMPL_WIDTH),
		13775 => to_signed(31747, LUT_AMPL_WIDTH),
		13776 => to_signed(31748, LUT_AMPL_WIDTH),
		13777 => to_signed(31749, LUT_AMPL_WIDTH),
		13778 => to_signed(31750, LUT_AMPL_WIDTH),
		13779 => to_signed(31750, LUT_AMPL_WIDTH),
		13780 => to_signed(31751, LUT_AMPL_WIDTH),
		13781 => to_signed(31752, LUT_AMPL_WIDTH),
		13782 => to_signed(31753, LUT_AMPL_WIDTH),
		13783 => to_signed(31753, LUT_AMPL_WIDTH),
		13784 => to_signed(31754, LUT_AMPL_WIDTH),
		13785 => to_signed(31755, LUT_AMPL_WIDTH),
		13786 => to_signed(31756, LUT_AMPL_WIDTH),
		13787 => to_signed(31757, LUT_AMPL_WIDTH),
		13788 => to_signed(31757, LUT_AMPL_WIDTH),
		13789 => to_signed(31758, LUT_AMPL_WIDTH),
		13790 => to_signed(31759, LUT_AMPL_WIDTH),
		13791 => to_signed(31760, LUT_AMPL_WIDTH),
		13792 => to_signed(31760, LUT_AMPL_WIDTH),
		13793 => to_signed(31761, LUT_AMPL_WIDTH),
		13794 => to_signed(31762, LUT_AMPL_WIDTH),
		13795 => to_signed(31763, LUT_AMPL_WIDTH),
		13796 => to_signed(31764, LUT_AMPL_WIDTH),
		13797 => to_signed(31764, LUT_AMPL_WIDTH),
		13798 => to_signed(31765, LUT_AMPL_WIDTH),
		13799 => to_signed(31766, LUT_AMPL_WIDTH),
		13800 => to_signed(31767, LUT_AMPL_WIDTH),
		13801 => to_signed(31767, LUT_AMPL_WIDTH),
		13802 => to_signed(31768, LUT_AMPL_WIDTH),
		13803 => to_signed(31769, LUT_AMPL_WIDTH),
		13804 => to_signed(31770, LUT_AMPL_WIDTH),
		13805 => to_signed(31770, LUT_AMPL_WIDTH),
		13806 => to_signed(31771, LUT_AMPL_WIDTH),
		13807 => to_signed(31772, LUT_AMPL_WIDTH),
		13808 => to_signed(31773, LUT_AMPL_WIDTH),
		13809 => to_signed(31774, LUT_AMPL_WIDTH),
		13810 => to_signed(31774, LUT_AMPL_WIDTH),
		13811 => to_signed(31775, LUT_AMPL_WIDTH),
		13812 => to_signed(31776, LUT_AMPL_WIDTH),
		13813 => to_signed(31777, LUT_AMPL_WIDTH),
		13814 => to_signed(31777, LUT_AMPL_WIDTH),
		13815 => to_signed(31778, LUT_AMPL_WIDTH),
		13816 => to_signed(31779, LUT_AMPL_WIDTH),
		13817 => to_signed(31780, LUT_AMPL_WIDTH),
		13818 => to_signed(31780, LUT_AMPL_WIDTH),
		13819 => to_signed(31781, LUT_AMPL_WIDTH),
		13820 => to_signed(31782, LUT_AMPL_WIDTH),
		13821 => to_signed(31783, LUT_AMPL_WIDTH),
		13822 => to_signed(31783, LUT_AMPL_WIDTH),
		13823 => to_signed(31784, LUT_AMPL_WIDTH),
		13824 => to_signed(31785, LUT_AMPL_WIDTH),
		13825 => to_signed(31786, LUT_AMPL_WIDTH),
		13826 => to_signed(31787, LUT_AMPL_WIDTH),
		13827 => to_signed(31787, LUT_AMPL_WIDTH),
		13828 => to_signed(31788, LUT_AMPL_WIDTH),
		13829 => to_signed(31789, LUT_AMPL_WIDTH),
		13830 => to_signed(31790, LUT_AMPL_WIDTH),
		13831 => to_signed(31790, LUT_AMPL_WIDTH),
		13832 => to_signed(31791, LUT_AMPL_WIDTH),
		13833 => to_signed(31792, LUT_AMPL_WIDTH),
		13834 => to_signed(31793, LUT_AMPL_WIDTH),
		13835 => to_signed(31793, LUT_AMPL_WIDTH),
		13836 => to_signed(31794, LUT_AMPL_WIDTH),
		13837 => to_signed(31795, LUT_AMPL_WIDTH),
		13838 => to_signed(31796, LUT_AMPL_WIDTH),
		13839 => to_signed(31796, LUT_AMPL_WIDTH),
		13840 => to_signed(31797, LUT_AMPL_WIDTH),
		13841 => to_signed(31798, LUT_AMPL_WIDTH),
		13842 => to_signed(31799, LUT_AMPL_WIDTH),
		13843 => to_signed(31799, LUT_AMPL_WIDTH),
		13844 => to_signed(31800, LUT_AMPL_WIDTH),
		13845 => to_signed(31801, LUT_AMPL_WIDTH),
		13846 => to_signed(31802, LUT_AMPL_WIDTH),
		13847 => to_signed(31802, LUT_AMPL_WIDTH),
		13848 => to_signed(31803, LUT_AMPL_WIDTH),
		13849 => to_signed(31804, LUT_AMPL_WIDTH),
		13850 => to_signed(31805, LUT_AMPL_WIDTH),
		13851 => to_signed(31806, LUT_AMPL_WIDTH),
		13852 => to_signed(31806, LUT_AMPL_WIDTH),
		13853 => to_signed(31807, LUT_AMPL_WIDTH),
		13854 => to_signed(31808, LUT_AMPL_WIDTH),
		13855 => to_signed(31809, LUT_AMPL_WIDTH),
		13856 => to_signed(31809, LUT_AMPL_WIDTH),
		13857 => to_signed(31810, LUT_AMPL_WIDTH),
		13858 => to_signed(31811, LUT_AMPL_WIDTH),
		13859 => to_signed(31812, LUT_AMPL_WIDTH),
		13860 => to_signed(31812, LUT_AMPL_WIDTH),
		13861 => to_signed(31813, LUT_AMPL_WIDTH),
		13862 => to_signed(31814, LUT_AMPL_WIDTH),
		13863 => to_signed(31815, LUT_AMPL_WIDTH),
		13864 => to_signed(31815, LUT_AMPL_WIDTH),
		13865 => to_signed(31816, LUT_AMPL_WIDTH),
		13866 => to_signed(31817, LUT_AMPL_WIDTH),
		13867 => to_signed(31818, LUT_AMPL_WIDTH),
		13868 => to_signed(31818, LUT_AMPL_WIDTH),
		13869 => to_signed(31819, LUT_AMPL_WIDTH),
		13870 => to_signed(31820, LUT_AMPL_WIDTH),
		13871 => to_signed(31821, LUT_AMPL_WIDTH),
		13872 => to_signed(31821, LUT_AMPL_WIDTH),
		13873 => to_signed(31822, LUT_AMPL_WIDTH),
		13874 => to_signed(31823, LUT_AMPL_WIDTH),
		13875 => to_signed(31824, LUT_AMPL_WIDTH),
		13876 => to_signed(31824, LUT_AMPL_WIDTH),
		13877 => to_signed(31825, LUT_AMPL_WIDTH),
		13878 => to_signed(31826, LUT_AMPL_WIDTH),
		13879 => to_signed(31827, LUT_AMPL_WIDTH),
		13880 => to_signed(31827, LUT_AMPL_WIDTH),
		13881 => to_signed(31828, LUT_AMPL_WIDTH),
		13882 => to_signed(31829, LUT_AMPL_WIDTH),
		13883 => to_signed(31830, LUT_AMPL_WIDTH),
		13884 => to_signed(31830, LUT_AMPL_WIDTH),
		13885 => to_signed(31831, LUT_AMPL_WIDTH),
		13886 => to_signed(31832, LUT_AMPL_WIDTH),
		13887 => to_signed(31833, LUT_AMPL_WIDTH),
		13888 => to_signed(31833, LUT_AMPL_WIDTH),
		13889 => to_signed(31834, LUT_AMPL_WIDTH),
		13890 => to_signed(31835, LUT_AMPL_WIDTH),
		13891 => to_signed(31836, LUT_AMPL_WIDTH),
		13892 => to_signed(31836, LUT_AMPL_WIDTH),
		13893 => to_signed(31837, LUT_AMPL_WIDTH),
		13894 => to_signed(31838, LUT_AMPL_WIDTH),
		13895 => to_signed(31838, LUT_AMPL_WIDTH),
		13896 => to_signed(31839, LUT_AMPL_WIDTH),
		13897 => to_signed(31840, LUT_AMPL_WIDTH),
		13898 => to_signed(31841, LUT_AMPL_WIDTH),
		13899 => to_signed(31841, LUT_AMPL_WIDTH),
		13900 => to_signed(31842, LUT_AMPL_WIDTH),
		13901 => to_signed(31843, LUT_AMPL_WIDTH),
		13902 => to_signed(31844, LUT_AMPL_WIDTH),
		13903 => to_signed(31844, LUT_AMPL_WIDTH),
		13904 => to_signed(31845, LUT_AMPL_WIDTH),
		13905 => to_signed(31846, LUT_AMPL_WIDTH),
		13906 => to_signed(31847, LUT_AMPL_WIDTH),
		13907 => to_signed(31847, LUT_AMPL_WIDTH),
		13908 => to_signed(31848, LUT_AMPL_WIDTH),
		13909 => to_signed(31849, LUT_AMPL_WIDTH),
		13910 => to_signed(31850, LUT_AMPL_WIDTH),
		13911 => to_signed(31850, LUT_AMPL_WIDTH),
		13912 => to_signed(31851, LUT_AMPL_WIDTH),
		13913 => to_signed(31852, LUT_AMPL_WIDTH),
		13914 => to_signed(31853, LUT_AMPL_WIDTH),
		13915 => to_signed(31853, LUT_AMPL_WIDTH),
		13916 => to_signed(31854, LUT_AMPL_WIDTH),
		13917 => to_signed(31855, LUT_AMPL_WIDTH),
		13918 => to_signed(31855, LUT_AMPL_WIDTH),
		13919 => to_signed(31856, LUT_AMPL_WIDTH),
		13920 => to_signed(31857, LUT_AMPL_WIDTH),
		13921 => to_signed(31858, LUT_AMPL_WIDTH),
		13922 => to_signed(31858, LUT_AMPL_WIDTH),
		13923 => to_signed(31859, LUT_AMPL_WIDTH),
		13924 => to_signed(31860, LUT_AMPL_WIDTH),
		13925 => to_signed(31861, LUT_AMPL_WIDTH),
		13926 => to_signed(31861, LUT_AMPL_WIDTH),
		13927 => to_signed(31862, LUT_AMPL_WIDTH),
		13928 => to_signed(31863, LUT_AMPL_WIDTH),
		13929 => to_signed(31864, LUT_AMPL_WIDTH),
		13930 => to_signed(31864, LUT_AMPL_WIDTH),
		13931 => to_signed(31865, LUT_AMPL_WIDTH),
		13932 => to_signed(31866, LUT_AMPL_WIDTH),
		13933 => to_signed(31866, LUT_AMPL_WIDTH),
		13934 => to_signed(31867, LUT_AMPL_WIDTH),
		13935 => to_signed(31868, LUT_AMPL_WIDTH),
		13936 => to_signed(31869, LUT_AMPL_WIDTH),
		13937 => to_signed(31869, LUT_AMPL_WIDTH),
		13938 => to_signed(31870, LUT_AMPL_WIDTH),
		13939 => to_signed(31871, LUT_AMPL_WIDTH),
		13940 => to_signed(31872, LUT_AMPL_WIDTH),
		13941 => to_signed(31872, LUT_AMPL_WIDTH),
		13942 => to_signed(31873, LUT_AMPL_WIDTH),
		13943 => to_signed(31874, LUT_AMPL_WIDTH),
		13944 => to_signed(31875, LUT_AMPL_WIDTH),
		13945 => to_signed(31875, LUT_AMPL_WIDTH),
		13946 => to_signed(31876, LUT_AMPL_WIDTH),
		13947 => to_signed(31877, LUT_AMPL_WIDTH),
		13948 => to_signed(31877, LUT_AMPL_WIDTH),
		13949 => to_signed(31878, LUT_AMPL_WIDTH),
		13950 => to_signed(31879, LUT_AMPL_WIDTH),
		13951 => to_signed(31880, LUT_AMPL_WIDTH),
		13952 => to_signed(31880, LUT_AMPL_WIDTH),
		13953 => to_signed(31881, LUT_AMPL_WIDTH),
		13954 => to_signed(31882, LUT_AMPL_WIDTH),
		13955 => to_signed(31882, LUT_AMPL_WIDTH),
		13956 => to_signed(31883, LUT_AMPL_WIDTH),
		13957 => to_signed(31884, LUT_AMPL_WIDTH),
		13958 => to_signed(31885, LUT_AMPL_WIDTH),
		13959 => to_signed(31885, LUT_AMPL_WIDTH),
		13960 => to_signed(31886, LUT_AMPL_WIDTH),
		13961 => to_signed(31887, LUT_AMPL_WIDTH),
		13962 => to_signed(31888, LUT_AMPL_WIDTH),
		13963 => to_signed(31888, LUT_AMPL_WIDTH),
		13964 => to_signed(31889, LUT_AMPL_WIDTH),
		13965 => to_signed(31890, LUT_AMPL_WIDTH),
		13966 => to_signed(31890, LUT_AMPL_WIDTH),
		13967 => to_signed(31891, LUT_AMPL_WIDTH),
		13968 => to_signed(31892, LUT_AMPL_WIDTH),
		13969 => to_signed(31893, LUT_AMPL_WIDTH),
		13970 => to_signed(31893, LUT_AMPL_WIDTH),
		13971 => to_signed(31894, LUT_AMPL_WIDTH),
		13972 => to_signed(31895, LUT_AMPL_WIDTH),
		13973 => to_signed(31896, LUT_AMPL_WIDTH),
		13974 => to_signed(31896, LUT_AMPL_WIDTH),
		13975 => to_signed(31897, LUT_AMPL_WIDTH),
		13976 => to_signed(31898, LUT_AMPL_WIDTH),
		13977 => to_signed(31898, LUT_AMPL_WIDTH),
		13978 => to_signed(31899, LUT_AMPL_WIDTH),
		13979 => to_signed(31900, LUT_AMPL_WIDTH),
		13980 => to_signed(31901, LUT_AMPL_WIDTH),
		13981 => to_signed(31901, LUT_AMPL_WIDTH),
		13982 => to_signed(31902, LUT_AMPL_WIDTH),
		13983 => to_signed(31903, LUT_AMPL_WIDTH),
		13984 => to_signed(31903, LUT_AMPL_WIDTH),
		13985 => to_signed(31904, LUT_AMPL_WIDTH),
		13986 => to_signed(31905, LUT_AMPL_WIDTH),
		13987 => to_signed(31906, LUT_AMPL_WIDTH),
		13988 => to_signed(31906, LUT_AMPL_WIDTH),
		13989 => to_signed(31907, LUT_AMPL_WIDTH),
		13990 => to_signed(31908, LUT_AMPL_WIDTH),
		13991 => to_signed(31908, LUT_AMPL_WIDTH),
		13992 => to_signed(31909, LUT_AMPL_WIDTH),
		13993 => to_signed(31910, LUT_AMPL_WIDTH),
		13994 => to_signed(31911, LUT_AMPL_WIDTH),
		13995 => to_signed(31911, LUT_AMPL_WIDTH),
		13996 => to_signed(31912, LUT_AMPL_WIDTH),
		13997 => to_signed(31913, LUT_AMPL_WIDTH),
		13998 => to_signed(31913, LUT_AMPL_WIDTH),
		13999 => to_signed(31914, LUT_AMPL_WIDTH),
		14000 => to_signed(31915, LUT_AMPL_WIDTH),
		14001 => to_signed(31916, LUT_AMPL_WIDTH),
		14002 => to_signed(31916, LUT_AMPL_WIDTH),
		14003 => to_signed(31917, LUT_AMPL_WIDTH),
		14004 => to_signed(31918, LUT_AMPL_WIDTH),
		14005 => to_signed(31918, LUT_AMPL_WIDTH),
		14006 => to_signed(31919, LUT_AMPL_WIDTH),
		14007 => to_signed(31920, LUT_AMPL_WIDTH),
		14008 => to_signed(31921, LUT_AMPL_WIDTH),
		14009 => to_signed(31921, LUT_AMPL_WIDTH),
		14010 => to_signed(31922, LUT_AMPL_WIDTH),
		14011 => to_signed(31923, LUT_AMPL_WIDTH),
		14012 => to_signed(31923, LUT_AMPL_WIDTH),
		14013 => to_signed(31924, LUT_AMPL_WIDTH),
		14014 => to_signed(31925, LUT_AMPL_WIDTH),
		14015 => to_signed(31925, LUT_AMPL_WIDTH),
		14016 => to_signed(31926, LUT_AMPL_WIDTH),
		14017 => to_signed(31927, LUT_AMPL_WIDTH),
		14018 => to_signed(31928, LUT_AMPL_WIDTH),
		14019 => to_signed(31928, LUT_AMPL_WIDTH),
		14020 => to_signed(31929, LUT_AMPL_WIDTH),
		14021 => to_signed(31930, LUT_AMPL_WIDTH),
		14022 => to_signed(31930, LUT_AMPL_WIDTH),
		14023 => to_signed(31931, LUT_AMPL_WIDTH),
		14024 => to_signed(31932, LUT_AMPL_WIDTH),
		14025 => to_signed(31933, LUT_AMPL_WIDTH),
		14026 => to_signed(31933, LUT_AMPL_WIDTH),
		14027 => to_signed(31934, LUT_AMPL_WIDTH),
		14028 => to_signed(31935, LUT_AMPL_WIDTH),
		14029 => to_signed(31935, LUT_AMPL_WIDTH),
		14030 => to_signed(31936, LUT_AMPL_WIDTH),
		14031 => to_signed(31937, LUT_AMPL_WIDTH),
		14032 => to_signed(31937, LUT_AMPL_WIDTH),
		14033 => to_signed(31938, LUT_AMPL_WIDTH),
		14034 => to_signed(31939, LUT_AMPL_WIDTH),
		14035 => to_signed(31940, LUT_AMPL_WIDTH),
		14036 => to_signed(31940, LUT_AMPL_WIDTH),
		14037 => to_signed(31941, LUT_AMPL_WIDTH),
		14038 => to_signed(31942, LUT_AMPL_WIDTH),
		14039 => to_signed(31942, LUT_AMPL_WIDTH),
		14040 => to_signed(31943, LUT_AMPL_WIDTH),
		14041 => to_signed(31944, LUT_AMPL_WIDTH),
		14042 => to_signed(31944, LUT_AMPL_WIDTH),
		14043 => to_signed(31945, LUT_AMPL_WIDTH),
		14044 => to_signed(31946, LUT_AMPL_WIDTH),
		14045 => to_signed(31947, LUT_AMPL_WIDTH),
		14046 => to_signed(31947, LUT_AMPL_WIDTH),
		14047 => to_signed(31948, LUT_AMPL_WIDTH),
		14048 => to_signed(31949, LUT_AMPL_WIDTH),
		14049 => to_signed(31949, LUT_AMPL_WIDTH),
		14050 => to_signed(31950, LUT_AMPL_WIDTH),
		14051 => to_signed(31951, LUT_AMPL_WIDTH),
		14052 => to_signed(31951, LUT_AMPL_WIDTH),
		14053 => to_signed(31952, LUT_AMPL_WIDTH),
		14054 => to_signed(31953, LUT_AMPL_WIDTH),
		14055 => to_signed(31954, LUT_AMPL_WIDTH),
		14056 => to_signed(31954, LUT_AMPL_WIDTH),
		14057 => to_signed(31955, LUT_AMPL_WIDTH),
		14058 => to_signed(31956, LUT_AMPL_WIDTH),
		14059 => to_signed(31956, LUT_AMPL_WIDTH),
		14060 => to_signed(31957, LUT_AMPL_WIDTH),
		14061 => to_signed(31958, LUT_AMPL_WIDTH),
		14062 => to_signed(31958, LUT_AMPL_WIDTH),
		14063 => to_signed(31959, LUT_AMPL_WIDTH),
		14064 => to_signed(31960, LUT_AMPL_WIDTH),
		14065 => to_signed(31960, LUT_AMPL_WIDTH),
		14066 => to_signed(31961, LUT_AMPL_WIDTH),
		14067 => to_signed(31962, LUT_AMPL_WIDTH),
		14068 => to_signed(31963, LUT_AMPL_WIDTH),
		14069 => to_signed(31963, LUT_AMPL_WIDTH),
		14070 => to_signed(31964, LUT_AMPL_WIDTH),
		14071 => to_signed(31965, LUT_AMPL_WIDTH),
		14072 => to_signed(31965, LUT_AMPL_WIDTH),
		14073 => to_signed(31966, LUT_AMPL_WIDTH),
		14074 => to_signed(31967, LUT_AMPL_WIDTH),
		14075 => to_signed(31967, LUT_AMPL_WIDTH),
		14076 => to_signed(31968, LUT_AMPL_WIDTH),
		14077 => to_signed(31969, LUT_AMPL_WIDTH),
		14078 => to_signed(31969, LUT_AMPL_WIDTH),
		14079 => to_signed(31970, LUT_AMPL_WIDTH),
		14080 => to_signed(31971, LUT_AMPL_WIDTH),
		14081 => to_signed(31972, LUT_AMPL_WIDTH),
		14082 => to_signed(31972, LUT_AMPL_WIDTH),
		14083 => to_signed(31973, LUT_AMPL_WIDTH),
		14084 => to_signed(31974, LUT_AMPL_WIDTH),
		14085 => to_signed(31974, LUT_AMPL_WIDTH),
		14086 => to_signed(31975, LUT_AMPL_WIDTH),
		14087 => to_signed(31976, LUT_AMPL_WIDTH),
		14088 => to_signed(31976, LUT_AMPL_WIDTH),
		14089 => to_signed(31977, LUT_AMPL_WIDTH),
		14090 => to_signed(31978, LUT_AMPL_WIDTH),
		14091 => to_signed(31978, LUT_AMPL_WIDTH),
		14092 => to_signed(31979, LUT_AMPL_WIDTH),
		14093 => to_signed(31980, LUT_AMPL_WIDTH),
		14094 => to_signed(31980, LUT_AMPL_WIDTH),
		14095 => to_signed(31981, LUT_AMPL_WIDTH),
		14096 => to_signed(31982, LUT_AMPL_WIDTH),
		14097 => to_signed(31982, LUT_AMPL_WIDTH),
		14098 => to_signed(31983, LUT_AMPL_WIDTH),
		14099 => to_signed(31984, LUT_AMPL_WIDTH),
		14100 => to_signed(31985, LUT_AMPL_WIDTH),
		14101 => to_signed(31985, LUT_AMPL_WIDTH),
		14102 => to_signed(31986, LUT_AMPL_WIDTH),
		14103 => to_signed(31987, LUT_AMPL_WIDTH),
		14104 => to_signed(31987, LUT_AMPL_WIDTH),
		14105 => to_signed(31988, LUT_AMPL_WIDTH),
		14106 => to_signed(31989, LUT_AMPL_WIDTH),
		14107 => to_signed(31989, LUT_AMPL_WIDTH),
		14108 => to_signed(31990, LUT_AMPL_WIDTH),
		14109 => to_signed(31991, LUT_AMPL_WIDTH),
		14110 => to_signed(31991, LUT_AMPL_WIDTH),
		14111 => to_signed(31992, LUT_AMPL_WIDTH),
		14112 => to_signed(31993, LUT_AMPL_WIDTH),
		14113 => to_signed(31993, LUT_AMPL_WIDTH),
		14114 => to_signed(31994, LUT_AMPL_WIDTH),
		14115 => to_signed(31995, LUT_AMPL_WIDTH),
		14116 => to_signed(31995, LUT_AMPL_WIDTH),
		14117 => to_signed(31996, LUT_AMPL_WIDTH),
		14118 => to_signed(31997, LUT_AMPL_WIDTH),
		14119 => to_signed(31997, LUT_AMPL_WIDTH),
		14120 => to_signed(31998, LUT_AMPL_WIDTH),
		14121 => to_signed(31999, LUT_AMPL_WIDTH),
		14122 => to_signed(31999, LUT_AMPL_WIDTH),
		14123 => to_signed(32000, LUT_AMPL_WIDTH),
		14124 => to_signed(32001, LUT_AMPL_WIDTH),
		14125 => to_signed(32002, LUT_AMPL_WIDTH),
		14126 => to_signed(32002, LUT_AMPL_WIDTH),
		14127 => to_signed(32003, LUT_AMPL_WIDTH),
		14128 => to_signed(32004, LUT_AMPL_WIDTH),
		14129 => to_signed(32004, LUT_AMPL_WIDTH),
		14130 => to_signed(32005, LUT_AMPL_WIDTH),
		14131 => to_signed(32006, LUT_AMPL_WIDTH),
		14132 => to_signed(32006, LUT_AMPL_WIDTH),
		14133 => to_signed(32007, LUT_AMPL_WIDTH),
		14134 => to_signed(32008, LUT_AMPL_WIDTH),
		14135 => to_signed(32008, LUT_AMPL_WIDTH),
		14136 => to_signed(32009, LUT_AMPL_WIDTH),
		14137 => to_signed(32010, LUT_AMPL_WIDTH),
		14138 => to_signed(32010, LUT_AMPL_WIDTH),
		14139 => to_signed(32011, LUT_AMPL_WIDTH),
		14140 => to_signed(32012, LUT_AMPL_WIDTH),
		14141 => to_signed(32012, LUT_AMPL_WIDTH),
		14142 => to_signed(32013, LUT_AMPL_WIDTH),
		14143 => to_signed(32014, LUT_AMPL_WIDTH),
		14144 => to_signed(32014, LUT_AMPL_WIDTH),
		14145 => to_signed(32015, LUT_AMPL_WIDTH),
		14146 => to_signed(32016, LUT_AMPL_WIDTH),
		14147 => to_signed(32016, LUT_AMPL_WIDTH),
		14148 => to_signed(32017, LUT_AMPL_WIDTH),
		14149 => to_signed(32018, LUT_AMPL_WIDTH),
		14150 => to_signed(32018, LUT_AMPL_WIDTH),
		14151 => to_signed(32019, LUT_AMPL_WIDTH),
		14152 => to_signed(32020, LUT_AMPL_WIDTH),
		14153 => to_signed(32020, LUT_AMPL_WIDTH),
		14154 => to_signed(32021, LUT_AMPL_WIDTH),
		14155 => to_signed(32022, LUT_AMPL_WIDTH),
		14156 => to_signed(32022, LUT_AMPL_WIDTH),
		14157 => to_signed(32023, LUT_AMPL_WIDTH),
		14158 => to_signed(32024, LUT_AMPL_WIDTH),
		14159 => to_signed(32024, LUT_AMPL_WIDTH),
		14160 => to_signed(32025, LUT_AMPL_WIDTH),
		14161 => to_signed(32026, LUT_AMPL_WIDTH),
		14162 => to_signed(32026, LUT_AMPL_WIDTH),
		14163 => to_signed(32027, LUT_AMPL_WIDTH),
		14164 => to_signed(32028, LUT_AMPL_WIDTH),
		14165 => to_signed(32028, LUT_AMPL_WIDTH),
		14166 => to_signed(32029, LUT_AMPL_WIDTH),
		14167 => to_signed(32030, LUT_AMPL_WIDTH),
		14168 => to_signed(32030, LUT_AMPL_WIDTH),
		14169 => to_signed(32031, LUT_AMPL_WIDTH),
		14170 => to_signed(32032, LUT_AMPL_WIDTH),
		14171 => to_signed(32032, LUT_AMPL_WIDTH),
		14172 => to_signed(32033, LUT_AMPL_WIDTH),
		14173 => to_signed(32034, LUT_AMPL_WIDTH),
		14174 => to_signed(32034, LUT_AMPL_WIDTH),
		14175 => to_signed(32035, LUT_AMPL_WIDTH),
		14176 => to_signed(32036, LUT_AMPL_WIDTH),
		14177 => to_signed(32036, LUT_AMPL_WIDTH),
		14178 => to_signed(32037, LUT_AMPL_WIDTH),
		14179 => to_signed(32038, LUT_AMPL_WIDTH),
		14180 => to_signed(32038, LUT_AMPL_WIDTH),
		14181 => to_signed(32039, LUT_AMPL_WIDTH),
		14182 => to_signed(32040, LUT_AMPL_WIDTH),
		14183 => to_signed(32040, LUT_AMPL_WIDTH),
		14184 => to_signed(32041, LUT_AMPL_WIDTH),
		14185 => to_signed(32041, LUT_AMPL_WIDTH),
		14186 => to_signed(32042, LUT_AMPL_WIDTH),
		14187 => to_signed(32043, LUT_AMPL_WIDTH),
		14188 => to_signed(32043, LUT_AMPL_WIDTH),
		14189 => to_signed(32044, LUT_AMPL_WIDTH),
		14190 => to_signed(32045, LUT_AMPL_WIDTH),
		14191 => to_signed(32045, LUT_AMPL_WIDTH),
		14192 => to_signed(32046, LUT_AMPL_WIDTH),
		14193 => to_signed(32047, LUT_AMPL_WIDTH),
		14194 => to_signed(32047, LUT_AMPL_WIDTH),
		14195 => to_signed(32048, LUT_AMPL_WIDTH),
		14196 => to_signed(32049, LUT_AMPL_WIDTH),
		14197 => to_signed(32049, LUT_AMPL_WIDTH),
		14198 => to_signed(32050, LUT_AMPL_WIDTH),
		14199 => to_signed(32051, LUT_AMPL_WIDTH),
		14200 => to_signed(32051, LUT_AMPL_WIDTH),
		14201 => to_signed(32052, LUT_AMPL_WIDTH),
		14202 => to_signed(32053, LUT_AMPL_WIDTH),
		14203 => to_signed(32053, LUT_AMPL_WIDTH),
		14204 => to_signed(32054, LUT_AMPL_WIDTH),
		14205 => to_signed(32055, LUT_AMPL_WIDTH),
		14206 => to_signed(32055, LUT_AMPL_WIDTH),
		14207 => to_signed(32056, LUT_AMPL_WIDTH),
		14208 => to_signed(32057, LUT_AMPL_WIDTH),
		14209 => to_signed(32057, LUT_AMPL_WIDTH),
		14210 => to_signed(32058, LUT_AMPL_WIDTH),
		14211 => to_signed(32058, LUT_AMPL_WIDTH),
		14212 => to_signed(32059, LUT_AMPL_WIDTH),
		14213 => to_signed(32060, LUT_AMPL_WIDTH),
		14214 => to_signed(32060, LUT_AMPL_WIDTH),
		14215 => to_signed(32061, LUT_AMPL_WIDTH),
		14216 => to_signed(32062, LUT_AMPL_WIDTH),
		14217 => to_signed(32062, LUT_AMPL_WIDTH),
		14218 => to_signed(32063, LUT_AMPL_WIDTH),
		14219 => to_signed(32064, LUT_AMPL_WIDTH),
		14220 => to_signed(32064, LUT_AMPL_WIDTH),
		14221 => to_signed(32065, LUT_AMPL_WIDTH),
		14222 => to_signed(32066, LUT_AMPL_WIDTH),
		14223 => to_signed(32066, LUT_AMPL_WIDTH),
		14224 => to_signed(32067, LUT_AMPL_WIDTH),
		14225 => to_signed(32068, LUT_AMPL_WIDTH),
		14226 => to_signed(32068, LUT_AMPL_WIDTH),
		14227 => to_signed(32069, LUT_AMPL_WIDTH),
		14228 => to_signed(32069, LUT_AMPL_WIDTH),
		14229 => to_signed(32070, LUT_AMPL_WIDTH),
		14230 => to_signed(32071, LUT_AMPL_WIDTH),
		14231 => to_signed(32071, LUT_AMPL_WIDTH),
		14232 => to_signed(32072, LUT_AMPL_WIDTH),
		14233 => to_signed(32073, LUT_AMPL_WIDTH),
		14234 => to_signed(32073, LUT_AMPL_WIDTH),
		14235 => to_signed(32074, LUT_AMPL_WIDTH),
		14236 => to_signed(32075, LUT_AMPL_WIDTH),
		14237 => to_signed(32075, LUT_AMPL_WIDTH),
		14238 => to_signed(32076, LUT_AMPL_WIDTH),
		14239 => to_signed(32077, LUT_AMPL_WIDTH),
		14240 => to_signed(32077, LUT_AMPL_WIDTH),
		14241 => to_signed(32078, LUT_AMPL_WIDTH),
		14242 => to_signed(32078, LUT_AMPL_WIDTH),
		14243 => to_signed(32079, LUT_AMPL_WIDTH),
		14244 => to_signed(32080, LUT_AMPL_WIDTH),
		14245 => to_signed(32080, LUT_AMPL_WIDTH),
		14246 => to_signed(32081, LUT_AMPL_WIDTH),
		14247 => to_signed(32082, LUT_AMPL_WIDTH),
		14248 => to_signed(32082, LUT_AMPL_WIDTH),
		14249 => to_signed(32083, LUT_AMPL_WIDTH),
		14250 => to_signed(32084, LUT_AMPL_WIDTH),
		14251 => to_signed(32084, LUT_AMPL_WIDTH),
		14252 => to_signed(32085, LUT_AMPL_WIDTH),
		14253 => to_signed(32086, LUT_AMPL_WIDTH),
		14254 => to_signed(32086, LUT_AMPL_WIDTH),
		14255 => to_signed(32087, LUT_AMPL_WIDTH),
		14256 => to_signed(32087, LUT_AMPL_WIDTH),
		14257 => to_signed(32088, LUT_AMPL_WIDTH),
		14258 => to_signed(32089, LUT_AMPL_WIDTH),
		14259 => to_signed(32089, LUT_AMPL_WIDTH),
		14260 => to_signed(32090, LUT_AMPL_WIDTH),
		14261 => to_signed(32091, LUT_AMPL_WIDTH),
		14262 => to_signed(32091, LUT_AMPL_WIDTH),
		14263 => to_signed(32092, LUT_AMPL_WIDTH),
		14264 => to_signed(32092, LUT_AMPL_WIDTH),
		14265 => to_signed(32093, LUT_AMPL_WIDTH),
		14266 => to_signed(32094, LUT_AMPL_WIDTH),
		14267 => to_signed(32094, LUT_AMPL_WIDTH),
		14268 => to_signed(32095, LUT_AMPL_WIDTH),
		14269 => to_signed(32096, LUT_AMPL_WIDTH),
		14270 => to_signed(32096, LUT_AMPL_WIDTH),
		14271 => to_signed(32097, LUT_AMPL_WIDTH),
		14272 => to_signed(32098, LUT_AMPL_WIDTH),
		14273 => to_signed(32098, LUT_AMPL_WIDTH),
		14274 => to_signed(32099, LUT_AMPL_WIDTH),
		14275 => to_signed(32099, LUT_AMPL_WIDTH),
		14276 => to_signed(32100, LUT_AMPL_WIDTH),
		14277 => to_signed(32101, LUT_AMPL_WIDTH),
		14278 => to_signed(32101, LUT_AMPL_WIDTH),
		14279 => to_signed(32102, LUT_AMPL_WIDTH),
		14280 => to_signed(32103, LUT_AMPL_WIDTH),
		14281 => to_signed(32103, LUT_AMPL_WIDTH),
		14282 => to_signed(32104, LUT_AMPL_WIDTH),
		14283 => to_signed(32104, LUT_AMPL_WIDTH),
		14284 => to_signed(32105, LUT_AMPL_WIDTH),
		14285 => to_signed(32106, LUT_AMPL_WIDTH),
		14286 => to_signed(32106, LUT_AMPL_WIDTH),
		14287 => to_signed(32107, LUT_AMPL_WIDTH),
		14288 => to_signed(32108, LUT_AMPL_WIDTH),
		14289 => to_signed(32108, LUT_AMPL_WIDTH),
		14290 => to_signed(32109, LUT_AMPL_WIDTH),
		14291 => to_signed(32110, LUT_AMPL_WIDTH),
		14292 => to_signed(32110, LUT_AMPL_WIDTH),
		14293 => to_signed(32111, LUT_AMPL_WIDTH),
		14294 => to_signed(32111, LUT_AMPL_WIDTH),
		14295 => to_signed(32112, LUT_AMPL_WIDTH),
		14296 => to_signed(32113, LUT_AMPL_WIDTH),
		14297 => to_signed(32113, LUT_AMPL_WIDTH),
		14298 => to_signed(32114, LUT_AMPL_WIDTH),
		14299 => to_signed(32115, LUT_AMPL_WIDTH),
		14300 => to_signed(32115, LUT_AMPL_WIDTH),
		14301 => to_signed(32116, LUT_AMPL_WIDTH),
		14302 => to_signed(32116, LUT_AMPL_WIDTH),
		14303 => to_signed(32117, LUT_AMPL_WIDTH),
		14304 => to_signed(32118, LUT_AMPL_WIDTH),
		14305 => to_signed(32118, LUT_AMPL_WIDTH),
		14306 => to_signed(32119, LUT_AMPL_WIDTH),
		14307 => to_signed(32119, LUT_AMPL_WIDTH),
		14308 => to_signed(32120, LUT_AMPL_WIDTH),
		14309 => to_signed(32121, LUT_AMPL_WIDTH),
		14310 => to_signed(32121, LUT_AMPL_WIDTH),
		14311 => to_signed(32122, LUT_AMPL_WIDTH),
		14312 => to_signed(32123, LUT_AMPL_WIDTH),
		14313 => to_signed(32123, LUT_AMPL_WIDTH),
		14314 => to_signed(32124, LUT_AMPL_WIDTH),
		14315 => to_signed(32124, LUT_AMPL_WIDTH),
		14316 => to_signed(32125, LUT_AMPL_WIDTH),
		14317 => to_signed(32126, LUT_AMPL_WIDTH),
		14318 => to_signed(32126, LUT_AMPL_WIDTH),
		14319 => to_signed(32127, LUT_AMPL_WIDTH),
		14320 => to_signed(32128, LUT_AMPL_WIDTH),
		14321 => to_signed(32128, LUT_AMPL_WIDTH),
		14322 => to_signed(32129, LUT_AMPL_WIDTH),
		14323 => to_signed(32129, LUT_AMPL_WIDTH),
		14324 => to_signed(32130, LUT_AMPL_WIDTH),
		14325 => to_signed(32131, LUT_AMPL_WIDTH),
		14326 => to_signed(32131, LUT_AMPL_WIDTH),
		14327 => to_signed(32132, LUT_AMPL_WIDTH),
		14328 => to_signed(32132, LUT_AMPL_WIDTH),
		14329 => to_signed(32133, LUT_AMPL_WIDTH),
		14330 => to_signed(32134, LUT_AMPL_WIDTH),
		14331 => to_signed(32134, LUT_AMPL_WIDTH),
		14332 => to_signed(32135, LUT_AMPL_WIDTH),
		14333 => to_signed(32136, LUT_AMPL_WIDTH),
		14334 => to_signed(32136, LUT_AMPL_WIDTH),
		14335 => to_signed(32137, LUT_AMPL_WIDTH),
		14336 => to_signed(32137, LUT_AMPL_WIDTH),
		14337 => to_signed(32138, LUT_AMPL_WIDTH),
		14338 => to_signed(32139, LUT_AMPL_WIDTH),
		14339 => to_signed(32139, LUT_AMPL_WIDTH),
		14340 => to_signed(32140, LUT_AMPL_WIDTH),
		14341 => to_signed(32140, LUT_AMPL_WIDTH),
		14342 => to_signed(32141, LUT_AMPL_WIDTH),
		14343 => to_signed(32142, LUT_AMPL_WIDTH),
		14344 => to_signed(32142, LUT_AMPL_WIDTH),
		14345 => to_signed(32143, LUT_AMPL_WIDTH),
		14346 => to_signed(32144, LUT_AMPL_WIDTH),
		14347 => to_signed(32144, LUT_AMPL_WIDTH),
		14348 => to_signed(32145, LUT_AMPL_WIDTH),
		14349 => to_signed(32145, LUT_AMPL_WIDTH),
		14350 => to_signed(32146, LUT_AMPL_WIDTH),
		14351 => to_signed(32147, LUT_AMPL_WIDTH),
		14352 => to_signed(32147, LUT_AMPL_WIDTH),
		14353 => to_signed(32148, LUT_AMPL_WIDTH),
		14354 => to_signed(32148, LUT_AMPL_WIDTH),
		14355 => to_signed(32149, LUT_AMPL_WIDTH),
		14356 => to_signed(32150, LUT_AMPL_WIDTH),
		14357 => to_signed(32150, LUT_AMPL_WIDTH),
		14358 => to_signed(32151, LUT_AMPL_WIDTH),
		14359 => to_signed(32151, LUT_AMPL_WIDTH),
		14360 => to_signed(32152, LUT_AMPL_WIDTH),
		14361 => to_signed(32153, LUT_AMPL_WIDTH),
		14362 => to_signed(32153, LUT_AMPL_WIDTH),
		14363 => to_signed(32154, LUT_AMPL_WIDTH),
		14364 => to_signed(32154, LUT_AMPL_WIDTH),
		14365 => to_signed(32155, LUT_AMPL_WIDTH),
		14366 => to_signed(32156, LUT_AMPL_WIDTH),
		14367 => to_signed(32156, LUT_AMPL_WIDTH),
		14368 => to_signed(32157, LUT_AMPL_WIDTH),
		14369 => to_signed(32157, LUT_AMPL_WIDTH),
		14370 => to_signed(32158, LUT_AMPL_WIDTH),
		14371 => to_signed(32159, LUT_AMPL_WIDTH),
		14372 => to_signed(32159, LUT_AMPL_WIDTH),
		14373 => to_signed(32160, LUT_AMPL_WIDTH),
		14374 => to_signed(32160, LUT_AMPL_WIDTH),
		14375 => to_signed(32161, LUT_AMPL_WIDTH),
		14376 => to_signed(32162, LUT_AMPL_WIDTH),
		14377 => to_signed(32162, LUT_AMPL_WIDTH),
		14378 => to_signed(32163, LUT_AMPL_WIDTH),
		14379 => to_signed(32163, LUT_AMPL_WIDTH),
		14380 => to_signed(32164, LUT_AMPL_WIDTH),
		14381 => to_signed(32165, LUT_AMPL_WIDTH),
		14382 => to_signed(32165, LUT_AMPL_WIDTH),
		14383 => to_signed(32166, LUT_AMPL_WIDTH),
		14384 => to_signed(32166, LUT_AMPL_WIDTH),
		14385 => to_signed(32167, LUT_AMPL_WIDTH),
		14386 => to_signed(32168, LUT_AMPL_WIDTH),
		14387 => to_signed(32168, LUT_AMPL_WIDTH),
		14388 => to_signed(32169, LUT_AMPL_WIDTH),
		14389 => to_signed(32169, LUT_AMPL_WIDTH),
		14390 => to_signed(32170, LUT_AMPL_WIDTH),
		14391 => to_signed(32171, LUT_AMPL_WIDTH),
		14392 => to_signed(32171, LUT_AMPL_WIDTH),
		14393 => to_signed(32172, LUT_AMPL_WIDTH),
		14394 => to_signed(32172, LUT_AMPL_WIDTH),
		14395 => to_signed(32173, LUT_AMPL_WIDTH),
		14396 => to_signed(32174, LUT_AMPL_WIDTH),
		14397 => to_signed(32174, LUT_AMPL_WIDTH),
		14398 => to_signed(32175, LUT_AMPL_WIDTH),
		14399 => to_signed(32175, LUT_AMPL_WIDTH),
		14400 => to_signed(32176, LUT_AMPL_WIDTH),
		14401 => to_signed(32177, LUT_AMPL_WIDTH),
		14402 => to_signed(32177, LUT_AMPL_WIDTH),
		14403 => to_signed(32178, LUT_AMPL_WIDTH),
		14404 => to_signed(32178, LUT_AMPL_WIDTH),
		14405 => to_signed(32179, LUT_AMPL_WIDTH),
		14406 => to_signed(32180, LUT_AMPL_WIDTH),
		14407 => to_signed(32180, LUT_AMPL_WIDTH),
		14408 => to_signed(32181, LUT_AMPL_WIDTH),
		14409 => to_signed(32181, LUT_AMPL_WIDTH),
		14410 => to_signed(32182, LUT_AMPL_WIDTH),
		14411 => to_signed(32183, LUT_AMPL_WIDTH),
		14412 => to_signed(32183, LUT_AMPL_WIDTH),
		14413 => to_signed(32184, LUT_AMPL_WIDTH),
		14414 => to_signed(32184, LUT_AMPL_WIDTH),
		14415 => to_signed(32185, LUT_AMPL_WIDTH),
		14416 => to_signed(32185, LUT_AMPL_WIDTH),
		14417 => to_signed(32186, LUT_AMPL_WIDTH),
		14418 => to_signed(32187, LUT_AMPL_WIDTH),
		14419 => to_signed(32187, LUT_AMPL_WIDTH),
		14420 => to_signed(32188, LUT_AMPL_WIDTH),
		14421 => to_signed(32188, LUT_AMPL_WIDTH),
		14422 => to_signed(32189, LUT_AMPL_WIDTH),
		14423 => to_signed(32190, LUT_AMPL_WIDTH),
		14424 => to_signed(32190, LUT_AMPL_WIDTH),
		14425 => to_signed(32191, LUT_AMPL_WIDTH),
		14426 => to_signed(32191, LUT_AMPL_WIDTH),
		14427 => to_signed(32192, LUT_AMPL_WIDTH),
		14428 => to_signed(32193, LUT_AMPL_WIDTH),
		14429 => to_signed(32193, LUT_AMPL_WIDTH),
		14430 => to_signed(32194, LUT_AMPL_WIDTH),
		14431 => to_signed(32194, LUT_AMPL_WIDTH),
		14432 => to_signed(32195, LUT_AMPL_WIDTH),
		14433 => to_signed(32195, LUT_AMPL_WIDTH),
		14434 => to_signed(32196, LUT_AMPL_WIDTH),
		14435 => to_signed(32197, LUT_AMPL_WIDTH),
		14436 => to_signed(32197, LUT_AMPL_WIDTH),
		14437 => to_signed(32198, LUT_AMPL_WIDTH),
		14438 => to_signed(32198, LUT_AMPL_WIDTH),
		14439 => to_signed(32199, LUT_AMPL_WIDTH),
		14440 => to_signed(32200, LUT_AMPL_WIDTH),
		14441 => to_signed(32200, LUT_AMPL_WIDTH),
		14442 => to_signed(32201, LUT_AMPL_WIDTH),
		14443 => to_signed(32201, LUT_AMPL_WIDTH),
		14444 => to_signed(32202, LUT_AMPL_WIDTH),
		14445 => to_signed(32202, LUT_AMPL_WIDTH),
		14446 => to_signed(32203, LUT_AMPL_WIDTH),
		14447 => to_signed(32204, LUT_AMPL_WIDTH),
		14448 => to_signed(32204, LUT_AMPL_WIDTH),
		14449 => to_signed(32205, LUT_AMPL_WIDTH),
		14450 => to_signed(32205, LUT_AMPL_WIDTH),
		14451 => to_signed(32206, LUT_AMPL_WIDTH),
		14452 => to_signed(32206, LUT_AMPL_WIDTH),
		14453 => to_signed(32207, LUT_AMPL_WIDTH),
		14454 => to_signed(32208, LUT_AMPL_WIDTH),
		14455 => to_signed(32208, LUT_AMPL_WIDTH),
		14456 => to_signed(32209, LUT_AMPL_WIDTH),
		14457 => to_signed(32209, LUT_AMPL_WIDTH),
		14458 => to_signed(32210, LUT_AMPL_WIDTH),
		14459 => to_signed(32211, LUT_AMPL_WIDTH),
		14460 => to_signed(32211, LUT_AMPL_WIDTH),
		14461 => to_signed(32212, LUT_AMPL_WIDTH),
		14462 => to_signed(32212, LUT_AMPL_WIDTH),
		14463 => to_signed(32213, LUT_AMPL_WIDTH),
		14464 => to_signed(32213, LUT_AMPL_WIDTH),
		14465 => to_signed(32214, LUT_AMPL_WIDTH),
		14466 => to_signed(32215, LUT_AMPL_WIDTH),
		14467 => to_signed(32215, LUT_AMPL_WIDTH),
		14468 => to_signed(32216, LUT_AMPL_WIDTH),
		14469 => to_signed(32216, LUT_AMPL_WIDTH),
		14470 => to_signed(32217, LUT_AMPL_WIDTH),
		14471 => to_signed(32217, LUT_AMPL_WIDTH),
		14472 => to_signed(32218, LUT_AMPL_WIDTH),
		14473 => to_signed(32219, LUT_AMPL_WIDTH),
		14474 => to_signed(32219, LUT_AMPL_WIDTH),
		14475 => to_signed(32220, LUT_AMPL_WIDTH),
		14476 => to_signed(32220, LUT_AMPL_WIDTH),
		14477 => to_signed(32221, LUT_AMPL_WIDTH),
		14478 => to_signed(32221, LUT_AMPL_WIDTH),
		14479 => to_signed(32222, LUT_AMPL_WIDTH),
		14480 => to_signed(32223, LUT_AMPL_WIDTH),
		14481 => to_signed(32223, LUT_AMPL_WIDTH),
		14482 => to_signed(32224, LUT_AMPL_WIDTH),
		14483 => to_signed(32224, LUT_AMPL_WIDTH),
		14484 => to_signed(32225, LUT_AMPL_WIDTH),
		14485 => to_signed(32225, LUT_AMPL_WIDTH),
		14486 => to_signed(32226, LUT_AMPL_WIDTH),
		14487 => to_signed(32227, LUT_AMPL_WIDTH),
		14488 => to_signed(32227, LUT_AMPL_WIDTH),
		14489 => to_signed(32228, LUT_AMPL_WIDTH),
		14490 => to_signed(32228, LUT_AMPL_WIDTH),
		14491 => to_signed(32229, LUT_AMPL_WIDTH),
		14492 => to_signed(32229, LUT_AMPL_WIDTH),
		14493 => to_signed(32230, LUT_AMPL_WIDTH),
		14494 => to_signed(32231, LUT_AMPL_WIDTH),
		14495 => to_signed(32231, LUT_AMPL_WIDTH),
		14496 => to_signed(32232, LUT_AMPL_WIDTH),
		14497 => to_signed(32232, LUT_AMPL_WIDTH),
		14498 => to_signed(32233, LUT_AMPL_WIDTH),
		14499 => to_signed(32233, LUT_AMPL_WIDTH),
		14500 => to_signed(32234, LUT_AMPL_WIDTH),
		14501 => to_signed(32234, LUT_AMPL_WIDTH),
		14502 => to_signed(32235, LUT_AMPL_WIDTH),
		14503 => to_signed(32236, LUT_AMPL_WIDTH),
		14504 => to_signed(32236, LUT_AMPL_WIDTH),
		14505 => to_signed(32237, LUT_AMPL_WIDTH),
		14506 => to_signed(32237, LUT_AMPL_WIDTH),
		14507 => to_signed(32238, LUT_AMPL_WIDTH),
		14508 => to_signed(32238, LUT_AMPL_WIDTH),
		14509 => to_signed(32239, LUT_AMPL_WIDTH),
		14510 => to_signed(32240, LUT_AMPL_WIDTH),
		14511 => to_signed(32240, LUT_AMPL_WIDTH),
		14512 => to_signed(32241, LUT_AMPL_WIDTH),
		14513 => to_signed(32241, LUT_AMPL_WIDTH),
		14514 => to_signed(32242, LUT_AMPL_WIDTH),
		14515 => to_signed(32242, LUT_AMPL_WIDTH),
		14516 => to_signed(32243, LUT_AMPL_WIDTH),
		14517 => to_signed(32243, LUT_AMPL_WIDTH),
		14518 => to_signed(32244, LUT_AMPL_WIDTH),
		14519 => to_signed(32245, LUT_AMPL_WIDTH),
		14520 => to_signed(32245, LUT_AMPL_WIDTH),
		14521 => to_signed(32246, LUT_AMPL_WIDTH),
		14522 => to_signed(32246, LUT_AMPL_WIDTH),
		14523 => to_signed(32247, LUT_AMPL_WIDTH),
		14524 => to_signed(32247, LUT_AMPL_WIDTH),
		14525 => to_signed(32248, LUT_AMPL_WIDTH),
		14526 => to_signed(32248, LUT_AMPL_WIDTH),
		14527 => to_signed(32249, LUT_AMPL_WIDTH),
		14528 => to_signed(32250, LUT_AMPL_WIDTH),
		14529 => to_signed(32250, LUT_AMPL_WIDTH),
		14530 => to_signed(32251, LUT_AMPL_WIDTH),
		14531 => to_signed(32251, LUT_AMPL_WIDTH),
		14532 => to_signed(32252, LUT_AMPL_WIDTH),
		14533 => to_signed(32252, LUT_AMPL_WIDTH),
		14534 => to_signed(32253, LUT_AMPL_WIDTH),
		14535 => to_signed(32253, LUT_AMPL_WIDTH),
		14536 => to_signed(32254, LUT_AMPL_WIDTH),
		14537 => to_signed(32255, LUT_AMPL_WIDTH),
		14538 => to_signed(32255, LUT_AMPL_WIDTH),
		14539 => to_signed(32256, LUT_AMPL_WIDTH),
		14540 => to_signed(32256, LUT_AMPL_WIDTH),
		14541 => to_signed(32257, LUT_AMPL_WIDTH),
		14542 => to_signed(32257, LUT_AMPL_WIDTH),
		14543 => to_signed(32258, LUT_AMPL_WIDTH),
		14544 => to_signed(32258, LUT_AMPL_WIDTH),
		14545 => to_signed(32259, LUT_AMPL_WIDTH),
		14546 => to_signed(32260, LUT_AMPL_WIDTH),
		14547 => to_signed(32260, LUT_AMPL_WIDTH),
		14548 => to_signed(32261, LUT_AMPL_WIDTH),
		14549 => to_signed(32261, LUT_AMPL_WIDTH),
		14550 => to_signed(32262, LUT_AMPL_WIDTH),
		14551 => to_signed(32262, LUT_AMPL_WIDTH),
		14552 => to_signed(32263, LUT_AMPL_WIDTH),
		14553 => to_signed(32263, LUT_AMPL_WIDTH),
		14554 => to_signed(32264, LUT_AMPL_WIDTH),
		14555 => to_signed(32265, LUT_AMPL_WIDTH),
		14556 => to_signed(32265, LUT_AMPL_WIDTH),
		14557 => to_signed(32266, LUT_AMPL_WIDTH),
		14558 => to_signed(32266, LUT_AMPL_WIDTH),
		14559 => to_signed(32267, LUT_AMPL_WIDTH),
		14560 => to_signed(32267, LUT_AMPL_WIDTH),
		14561 => to_signed(32268, LUT_AMPL_WIDTH),
		14562 => to_signed(32268, LUT_AMPL_WIDTH),
		14563 => to_signed(32269, LUT_AMPL_WIDTH),
		14564 => to_signed(32269, LUT_AMPL_WIDTH),
		14565 => to_signed(32270, LUT_AMPL_WIDTH),
		14566 => to_signed(32271, LUT_AMPL_WIDTH),
		14567 => to_signed(32271, LUT_AMPL_WIDTH),
		14568 => to_signed(32272, LUT_AMPL_WIDTH),
		14569 => to_signed(32272, LUT_AMPL_WIDTH),
		14570 => to_signed(32273, LUT_AMPL_WIDTH),
		14571 => to_signed(32273, LUT_AMPL_WIDTH),
		14572 => to_signed(32274, LUT_AMPL_WIDTH),
		14573 => to_signed(32274, LUT_AMPL_WIDTH),
		14574 => to_signed(32275, LUT_AMPL_WIDTH),
		14575 => to_signed(32275, LUT_AMPL_WIDTH),
		14576 => to_signed(32276, LUT_AMPL_WIDTH),
		14577 => to_signed(32277, LUT_AMPL_WIDTH),
		14578 => to_signed(32277, LUT_AMPL_WIDTH),
		14579 => to_signed(32278, LUT_AMPL_WIDTH),
		14580 => to_signed(32278, LUT_AMPL_WIDTH),
		14581 => to_signed(32279, LUT_AMPL_WIDTH),
		14582 => to_signed(32279, LUT_AMPL_WIDTH),
		14583 => to_signed(32280, LUT_AMPL_WIDTH),
		14584 => to_signed(32280, LUT_AMPL_WIDTH),
		14585 => to_signed(32281, LUT_AMPL_WIDTH),
		14586 => to_signed(32281, LUT_AMPL_WIDTH),
		14587 => to_signed(32282, LUT_AMPL_WIDTH),
		14588 => to_signed(32282, LUT_AMPL_WIDTH),
		14589 => to_signed(32283, LUT_AMPL_WIDTH),
		14590 => to_signed(32284, LUT_AMPL_WIDTH),
		14591 => to_signed(32284, LUT_AMPL_WIDTH),
		14592 => to_signed(32285, LUT_AMPL_WIDTH),
		14593 => to_signed(32285, LUT_AMPL_WIDTH),
		14594 => to_signed(32286, LUT_AMPL_WIDTH),
		14595 => to_signed(32286, LUT_AMPL_WIDTH),
		14596 => to_signed(32287, LUT_AMPL_WIDTH),
		14597 => to_signed(32287, LUT_AMPL_WIDTH),
		14598 => to_signed(32288, LUT_AMPL_WIDTH),
		14599 => to_signed(32288, LUT_AMPL_WIDTH),
		14600 => to_signed(32289, LUT_AMPL_WIDTH),
		14601 => to_signed(32289, LUT_AMPL_WIDTH),
		14602 => to_signed(32290, LUT_AMPL_WIDTH),
		14603 => to_signed(32290, LUT_AMPL_WIDTH),
		14604 => to_signed(32291, LUT_AMPL_WIDTH),
		14605 => to_signed(32292, LUT_AMPL_WIDTH),
		14606 => to_signed(32292, LUT_AMPL_WIDTH),
		14607 => to_signed(32293, LUT_AMPL_WIDTH),
		14608 => to_signed(32293, LUT_AMPL_WIDTH),
		14609 => to_signed(32294, LUT_AMPL_WIDTH),
		14610 => to_signed(32294, LUT_AMPL_WIDTH),
		14611 => to_signed(32295, LUT_AMPL_WIDTH),
		14612 => to_signed(32295, LUT_AMPL_WIDTH),
		14613 => to_signed(32296, LUT_AMPL_WIDTH),
		14614 => to_signed(32296, LUT_AMPL_WIDTH),
		14615 => to_signed(32297, LUT_AMPL_WIDTH),
		14616 => to_signed(32297, LUT_AMPL_WIDTH),
		14617 => to_signed(32298, LUT_AMPL_WIDTH),
		14618 => to_signed(32298, LUT_AMPL_WIDTH),
		14619 => to_signed(32299, LUT_AMPL_WIDTH),
		14620 => to_signed(32300, LUT_AMPL_WIDTH),
		14621 => to_signed(32300, LUT_AMPL_WIDTH),
		14622 => to_signed(32301, LUT_AMPL_WIDTH),
		14623 => to_signed(32301, LUT_AMPL_WIDTH),
		14624 => to_signed(32302, LUT_AMPL_WIDTH),
		14625 => to_signed(32302, LUT_AMPL_WIDTH),
		14626 => to_signed(32303, LUT_AMPL_WIDTH),
		14627 => to_signed(32303, LUT_AMPL_WIDTH),
		14628 => to_signed(32304, LUT_AMPL_WIDTH),
		14629 => to_signed(32304, LUT_AMPL_WIDTH),
		14630 => to_signed(32305, LUT_AMPL_WIDTH),
		14631 => to_signed(32305, LUT_AMPL_WIDTH),
		14632 => to_signed(32306, LUT_AMPL_WIDTH),
		14633 => to_signed(32306, LUT_AMPL_WIDTH),
		14634 => to_signed(32307, LUT_AMPL_WIDTH),
		14635 => to_signed(32307, LUT_AMPL_WIDTH),
		14636 => to_signed(32308, LUT_AMPL_WIDTH),
		14637 => to_signed(32308, LUT_AMPL_WIDTH),
		14638 => to_signed(32309, LUT_AMPL_WIDTH),
		14639 => to_signed(32310, LUT_AMPL_WIDTH),
		14640 => to_signed(32310, LUT_AMPL_WIDTH),
		14641 => to_signed(32311, LUT_AMPL_WIDTH),
		14642 => to_signed(32311, LUT_AMPL_WIDTH),
		14643 => to_signed(32312, LUT_AMPL_WIDTH),
		14644 => to_signed(32312, LUT_AMPL_WIDTH),
		14645 => to_signed(32313, LUT_AMPL_WIDTH),
		14646 => to_signed(32313, LUT_AMPL_WIDTH),
		14647 => to_signed(32314, LUT_AMPL_WIDTH),
		14648 => to_signed(32314, LUT_AMPL_WIDTH),
		14649 => to_signed(32315, LUT_AMPL_WIDTH),
		14650 => to_signed(32315, LUT_AMPL_WIDTH),
		14651 => to_signed(32316, LUT_AMPL_WIDTH),
		14652 => to_signed(32316, LUT_AMPL_WIDTH),
		14653 => to_signed(32317, LUT_AMPL_WIDTH),
		14654 => to_signed(32317, LUT_AMPL_WIDTH),
		14655 => to_signed(32318, LUT_AMPL_WIDTH),
		14656 => to_signed(32318, LUT_AMPL_WIDTH),
		14657 => to_signed(32319, LUT_AMPL_WIDTH),
		14658 => to_signed(32319, LUT_AMPL_WIDTH),
		14659 => to_signed(32320, LUT_AMPL_WIDTH),
		14660 => to_signed(32320, LUT_AMPL_WIDTH),
		14661 => to_signed(32321, LUT_AMPL_WIDTH),
		14662 => to_signed(32321, LUT_AMPL_WIDTH),
		14663 => to_signed(32322, LUT_AMPL_WIDTH),
		14664 => to_signed(32322, LUT_AMPL_WIDTH),
		14665 => to_signed(32323, LUT_AMPL_WIDTH),
		14666 => to_signed(32324, LUT_AMPL_WIDTH),
		14667 => to_signed(32324, LUT_AMPL_WIDTH),
		14668 => to_signed(32325, LUT_AMPL_WIDTH),
		14669 => to_signed(32325, LUT_AMPL_WIDTH),
		14670 => to_signed(32326, LUT_AMPL_WIDTH),
		14671 => to_signed(32326, LUT_AMPL_WIDTH),
		14672 => to_signed(32327, LUT_AMPL_WIDTH),
		14673 => to_signed(32327, LUT_AMPL_WIDTH),
		14674 => to_signed(32328, LUT_AMPL_WIDTH),
		14675 => to_signed(32328, LUT_AMPL_WIDTH),
		14676 => to_signed(32329, LUT_AMPL_WIDTH),
		14677 => to_signed(32329, LUT_AMPL_WIDTH),
		14678 => to_signed(32330, LUT_AMPL_WIDTH),
		14679 => to_signed(32330, LUT_AMPL_WIDTH),
		14680 => to_signed(32331, LUT_AMPL_WIDTH),
		14681 => to_signed(32331, LUT_AMPL_WIDTH),
		14682 => to_signed(32332, LUT_AMPL_WIDTH),
		14683 => to_signed(32332, LUT_AMPL_WIDTH),
		14684 => to_signed(32333, LUT_AMPL_WIDTH),
		14685 => to_signed(32333, LUT_AMPL_WIDTH),
		14686 => to_signed(32334, LUT_AMPL_WIDTH),
		14687 => to_signed(32334, LUT_AMPL_WIDTH),
		14688 => to_signed(32335, LUT_AMPL_WIDTH),
		14689 => to_signed(32335, LUT_AMPL_WIDTH),
		14690 => to_signed(32336, LUT_AMPL_WIDTH),
		14691 => to_signed(32336, LUT_AMPL_WIDTH),
		14692 => to_signed(32337, LUT_AMPL_WIDTH),
		14693 => to_signed(32337, LUT_AMPL_WIDTH),
		14694 => to_signed(32338, LUT_AMPL_WIDTH),
		14695 => to_signed(32338, LUT_AMPL_WIDTH),
		14696 => to_signed(32339, LUT_AMPL_WIDTH),
		14697 => to_signed(32339, LUT_AMPL_WIDTH),
		14698 => to_signed(32340, LUT_AMPL_WIDTH),
		14699 => to_signed(32340, LUT_AMPL_WIDTH),
		14700 => to_signed(32341, LUT_AMPL_WIDTH),
		14701 => to_signed(32341, LUT_AMPL_WIDTH),
		14702 => to_signed(32342, LUT_AMPL_WIDTH),
		14703 => to_signed(32342, LUT_AMPL_WIDTH),
		14704 => to_signed(32343, LUT_AMPL_WIDTH),
		14705 => to_signed(32343, LUT_AMPL_WIDTH),
		14706 => to_signed(32344, LUT_AMPL_WIDTH),
		14707 => to_signed(32344, LUT_AMPL_WIDTH),
		14708 => to_signed(32345, LUT_AMPL_WIDTH),
		14709 => to_signed(32345, LUT_AMPL_WIDTH),
		14710 => to_signed(32346, LUT_AMPL_WIDTH),
		14711 => to_signed(32346, LUT_AMPL_WIDTH),
		14712 => to_signed(32347, LUT_AMPL_WIDTH),
		14713 => to_signed(32347, LUT_AMPL_WIDTH),
		14714 => to_signed(32348, LUT_AMPL_WIDTH),
		14715 => to_signed(32348, LUT_AMPL_WIDTH),
		14716 => to_signed(32349, LUT_AMPL_WIDTH),
		14717 => to_signed(32349, LUT_AMPL_WIDTH),
		14718 => to_signed(32350, LUT_AMPL_WIDTH),
		14719 => to_signed(32350, LUT_AMPL_WIDTH),
		14720 => to_signed(32351, LUT_AMPL_WIDTH),
		14721 => to_signed(32351, LUT_AMPL_WIDTH),
		14722 => to_signed(32352, LUT_AMPL_WIDTH),
		14723 => to_signed(32352, LUT_AMPL_WIDTH),
		14724 => to_signed(32353, LUT_AMPL_WIDTH),
		14725 => to_signed(32353, LUT_AMPL_WIDTH),
		14726 => to_signed(32354, LUT_AMPL_WIDTH),
		14727 => to_signed(32354, LUT_AMPL_WIDTH),
		14728 => to_signed(32355, LUT_AMPL_WIDTH),
		14729 => to_signed(32355, LUT_AMPL_WIDTH),
		14730 => to_signed(32356, LUT_AMPL_WIDTH),
		14731 => to_signed(32356, LUT_AMPL_WIDTH),
		14732 => to_signed(32357, LUT_AMPL_WIDTH),
		14733 => to_signed(32357, LUT_AMPL_WIDTH),
		14734 => to_signed(32358, LUT_AMPL_WIDTH),
		14735 => to_signed(32358, LUT_AMPL_WIDTH),
		14736 => to_signed(32359, LUT_AMPL_WIDTH),
		14737 => to_signed(32359, LUT_AMPL_WIDTH),
		14738 => to_signed(32360, LUT_AMPL_WIDTH),
		14739 => to_signed(32360, LUT_AMPL_WIDTH),
		14740 => to_signed(32361, LUT_AMPL_WIDTH),
		14741 => to_signed(32361, LUT_AMPL_WIDTH),
		14742 => to_signed(32362, LUT_AMPL_WIDTH),
		14743 => to_signed(32362, LUT_AMPL_WIDTH),
		14744 => to_signed(32363, LUT_AMPL_WIDTH),
		14745 => to_signed(32363, LUT_AMPL_WIDTH),
		14746 => to_signed(32364, LUT_AMPL_WIDTH),
		14747 => to_signed(32364, LUT_AMPL_WIDTH),
		14748 => to_signed(32365, LUT_AMPL_WIDTH),
		14749 => to_signed(32365, LUT_AMPL_WIDTH),
		14750 => to_signed(32366, LUT_AMPL_WIDTH),
		14751 => to_signed(32366, LUT_AMPL_WIDTH),
		14752 => to_signed(32367, LUT_AMPL_WIDTH),
		14753 => to_signed(32367, LUT_AMPL_WIDTH),
		14754 => to_signed(32368, LUT_AMPL_WIDTH),
		14755 => to_signed(32368, LUT_AMPL_WIDTH),
		14756 => to_signed(32369, LUT_AMPL_WIDTH),
		14757 => to_signed(32369, LUT_AMPL_WIDTH),
		14758 => to_signed(32370, LUT_AMPL_WIDTH),
		14759 => to_signed(32370, LUT_AMPL_WIDTH),
		14760 => to_signed(32371, LUT_AMPL_WIDTH),
		14761 => to_signed(32371, LUT_AMPL_WIDTH),
		14762 => to_signed(32372, LUT_AMPL_WIDTH),
		14763 => to_signed(32372, LUT_AMPL_WIDTH),
		14764 => to_signed(32373, LUT_AMPL_WIDTH),
		14765 => to_signed(32373, LUT_AMPL_WIDTH),
		14766 => to_signed(32374, LUT_AMPL_WIDTH),
		14767 => to_signed(32374, LUT_AMPL_WIDTH),
		14768 => to_signed(32375, LUT_AMPL_WIDTH),
		14769 => to_signed(32375, LUT_AMPL_WIDTH),
		14770 => to_signed(32375, LUT_AMPL_WIDTH),
		14771 => to_signed(32376, LUT_AMPL_WIDTH),
		14772 => to_signed(32376, LUT_AMPL_WIDTH),
		14773 => to_signed(32377, LUT_AMPL_WIDTH),
		14774 => to_signed(32377, LUT_AMPL_WIDTH),
		14775 => to_signed(32378, LUT_AMPL_WIDTH),
		14776 => to_signed(32378, LUT_AMPL_WIDTH),
		14777 => to_signed(32379, LUT_AMPL_WIDTH),
		14778 => to_signed(32379, LUT_AMPL_WIDTH),
		14779 => to_signed(32380, LUT_AMPL_WIDTH),
		14780 => to_signed(32380, LUT_AMPL_WIDTH),
		14781 => to_signed(32381, LUT_AMPL_WIDTH),
		14782 => to_signed(32381, LUT_AMPL_WIDTH),
		14783 => to_signed(32382, LUT_AMPL_WIDTH),
		14784 => to_signed(32382, LUT_AMPL_WIDTH),
		14785 => to_signed(32383, LUT_AMPL_WIDTH),
		14786 => to_signed(32383, LUT_AMPL_WIDTH),
		14787 => to_signed(32384, LUT_AMPL_WIDTH),
		14788 => to_signed(32384, LUT_AMPL_WIDTH),
		14789 => to_signed(32385, LUT_AMPL_WIDTH),
		14790 => to_signed(32385, LUT_AMPL_WIDTH),
		14791 => to_signed(32386, LUT_AMPL_WIDTH),
		14792 => to_signed(32386, LUT_AMPL_WIDTH),
		14793 => to_signed(32387, LUT_AMPL_WIDTH),
		14794 => to_signed(32387, LUT_AMPL_WIDTH),
		14795 => to_signed(32387, LUT_AMPL_WIDTH),
		14796 => to_signed(32388, LUT_AMPL_WIDTH),
		14797 => to_signed(32388, LUT_AMPL_WIDTH),
		14798 => to_signed(32389, LUT_AMPL_WIDTH),
		14799 => to_signed(32389, LUT_AMPL_WIDTH),
		14800 => to_signed(32390, LUT_AMPL_WIDTH),
		14801 => to_signed(32390, LUT_AMPL_WIDTH),
		14802 => to_signed(32391, LUT_AMPL_WIDTH),
		14803 => to_signed(32391, LUT_AMPL_WIDTH),
		14804 => to_signed(32392, LUT_AMPL_WIDTH),
		14805 => to_signed(32392, LUT_AMPL_WIDTH),
		14806 => to_signed(32393, LUT_AMPL_WIDTH),
		14807 => to_signed(32393, LUT_AMPL_WIDTH),
		14808 => to_signed(32394, LUT_AMPL_WIDTH),
		14809 => to_signed(32394, LUT_AMPL_WIDTH),
		14810 => to_signed(32395, LUT_AMPL_WIDTH),
		14811 => to_signed(32395, LUT_AMPL_WIDTH),
		14812 => to_signed(32396, LUT_AMPL_WIDTH),
		14813 => to_signed(32396, LUT_AMPL_WIDTH),
		14814 => to_signed(32397, LUT_AMPL_WIDTH),
		14815 => to_signed(32397, LUT_AMPL_WIDTH),
		14816 => to_signed(32397, LUT_AMPL_WIDTH),
		14817 => to_signed(32398, LUT_AMPL_WIDTH),
		14818 => to_signed(32398, LUT_AMPL_WIDTH),
		14819 => to_signed(32399, LUT_AMPL_WIDTH),
		14820 => to_signed(32399, LUT_AMPL_WIDTH),
		14821 => to_signed(32400, LUT_AMPL_WIDTH),
		14822 => to_signed(32400, LUT_AMPL_WIDTH),
		14823 => to_signed(32401, LUT_AMPL_WIDTH),
		14824 => to_signed(32401, LUT_AMPL_WIDTH),
		14825 => to_signed(32402, LUT_AMPL_WIDTH),
		14826 => to_signed(32402, LUT_AMPL_WIDTH),
		14827 => to_signed(32403, LUT_AMPL_WIDTH),
		14828 => to_signed(32403, LUT_AMPL_WIDTH),
		14829 => to_signed(32404, LUT_AMPL_WIDTH),
		14830 => to_signed(32404, LUT_AMPL_WIDTH),
		14831 => to_signed(32404, LUT_AMPL_WIDTH),
		14832 => to_signed(32405, LUT_AMPL_WIDTH),
		14833 => to_signed(32405, LUT_AMPL_WIDTH),
		14834 => to_signed(32406, LUT_AMPL_WIDTH),
		14835 => to_signed(32406, LUT_AMPL_WIDTH),
		14836 => to_signed(32407, LUT_AMPL_WIDTH),
		14837 => to_signed(32407, LUT_AMPL_WIDTH),
		14838 => to_signed(32408, LUT_AMPL_WIDTH),
		14839 => to_signed(32408, LUT_AMPL_WIDTH),
		14840 => to_signed(32409, LUT_AMPL_WIDTH),
		14841 => to_signed(32409, LUT_AMPL_WIDTH),
		14842 => to_signed(32410, LUT_AMPL_WIDTH),
		14843 => to_signed(32410, LUT_AMPL_WIDTH),
		14844 => to_signed(32411, LUT_AMPL_WIDTH),
		14845 => to_signed(32411, LUT_AMPL_WIDTH),
		14846 => to_signed(32411, LUT_AMPL_WIDTH),
		14847 => to_signed(32412, LUT_AMPL_WIDTH),
		14848 => to_signed(32412, LUT_AMPL_WIDTH),
		14849 => to_signed(32413, LUT_AMPL_WIDTH),
		14850 => to_signed(32413, LUT_AMPL_WIDTH),
		14851 => to_signed(32414, LUT_AMPL_WIDTH),
		14852 => to_signed(32414, LUT_AMPL_WIDTH),
		14853 => to_signed(32415, LUT_AMPL_WIDTH),
		14854 => to_signed(32415, LUT_AMPL_WIDTH),
		14855 => to_signed(32416, LUT_AMPL_WIDTH),
		14856 => to_signed(32416, LUT_AMPL_WIDTH),
		14857 => to_signed(32416, LUT_AMPL_WIDTH),
		14858 => to_signed(32417, LUT_AMPL_WIDTH),
		14859 => to_signed(32417, LUT_AMPL_WIDTH),
		14860 => to_signed(32418, LUT_AMPL_WIDTH),
		14861 => to_signed(32418, LUT_AMPL_WIDTH),
		14862 => to_signed(32419, LUT_AMPL_WIDTH),
		14863 => to_signed(32419, LUT_AMPL_WIDTH),
		14864 => to_signed(32420, LUT_AMPL_WIDTH),
		14865 => to_signed(32420, LUT_AMPL_WIDTH),
		14866 => to_signed(32421, LUT_AMPL_WIDTH),
		14867 => to_signed(32421, LUT_AMPL_WIDTH),
		14868 => to_signed(32422, LUT_AMPL_WIDTH),
		14869 => to_signed(32422, LUT_AMPL_WIDTH),
		14870 => to_signed(32422, LUT_AMPL_WIDTH),
		14871 => to_signed(32423, LUT_AMPL_WIDTH),
		14872 => to_signed(32423, LUT_AMPL_WIDTH),
		14873 => to_signed(32424, LUT_AMPL_WIDTH),
		14874 => to_signed(32424, LUT_AMPL_WIDTH),
		14875 => to_signed(32425, LUT_AMPL_WIDTH),
		14876 => to_signed(32425, LUT_AMPL_WIDTH),
		14877 => to_signed(32426, LUT_AMPL_WIDTH),
		14878 => to_signed(32426, LUT_AMPL_WIDTH),
		14879 => to_signed(32426, LUT_AMPL_WIDTH),
		14880 => to_signed(32427, LUT_AMPL_WIDTH),
		14881 => to_signed(32427, LUT_AMPL_WIDTH),
		14882 => to_signed(32428, LUT_AMPL_WIDTH),
		14883 => to_signed(32428, LUT_AMPL_WIDTH),
		14884 => to_signed(32429, LUT_AMPL_WIDTH),
		14885 => to_signed(32429, LUT_AMPL_WIDTH),
		14886 => to_signed(32430, LUT_AMPL_WIDTH),
		14887 => to_signed(32430, LUT_AMPL_WIDTH),
		14888 => to_signed(32431, LUT_AMPL_WIDTH),
		14889 => to_signed(32431, LUT_AMPL_WIDTH),
		14890 => to_signed(32431, LUT_AMPL_WIDTH),
		14891 => to_signed(32432, LUT_AMPL_WIDTH),
		14892 => to_signed(32432, LUT_AMPL_WIDTH),
		14893 => to_signed(32433, LUT_AMPL_WIDTH),
		14894 => to_signed(32433, LUT_AMPL_WIDTH),
		14895 => to_signed(32434, LUT_AMPL_WIDTH),
		14896 => to_signed(32434, LUT_AMPL_WIDTH),
		14897 => to_signed(32435, LUT_AMPL_WIDTH),
		14898 => to_signed(32435, LUT_AMPL_WIDTH),
		14899 => to_signed(32435, LUT_AMPL_WIDTH),
		14900 => to_signed(32436, LUT_AMPL_WIDTH),
		14901 => to_signed(32436, LUT_AMPL_WIDTH),
		14902 => to_signed(32437, LUT_AMPL_WIDTH),
		14903 => to_signed(32437, LUT_AMPL_WIDTH),
		14904 => to_signed(32438, LUT_AMPL_WIDTH),
		14905 => to_signed(32438, LUT_AMPL_WIDTH),
		14906 => to_signed(32439, LUT_AMPL_WIDTH),
		14907 => to_signed(32439, LUT_AMPL_WIDTH),
		14908 => to_signed(32439, LUT_AMPL_WIDTH),
		14909 => to_signed(32440, LUT_AMPL_WIDTH),
		14910 => to_signed(32440, LUT_AMPL_WIDTH),
		14911 => to_signed(32441, LUT_AMPL_WIDTH),
		14912 => to_signed(32441, LUT_AMPL_WIDTH),
		14913 => to_signed(32442, LUT_AMPL_WIDTH),
		14914 => to_signed(32442, LUT_AMPL_WIDTH),
		14915 => to_signed(32443, LUT_AMPL_WIDTH),
		14916 => to_signed(32443, LUT_AMPL_WIDTH),
		14917 => to_signed(32443, LUT_AMPL_WIDTH),
		14918 => to_signed(32444, LUT_AMPL_WIDTH),
		14919 => to_signed(32444, LUT_AMPL_WIDTH),
		14920 => to_signed(32445, LUT_AMPL_WIDTH),
		14921 => to_signed(32445, LUT_AMPL_WIDTH),
		14922 => to_signed(32446, LUT_AMPL_WIDTH),
		14923 => to_signed(32446, LUT_AMPL_WIDTH),
		14924 => to_signed(32447, LUT_AMPL_WIDTH),
		14925 => to_signed(32447, LUT_AMPL_WIDTH),
		14926 => to_signed(32447, LUT_AMPL_WIDTH),
		14927 => to_signed(32448, LUT_AMPL_WIDTH),
		14928 => to_signed(32448, LUT_AMPL_WIDTH),
		14929 => to_signed(32449, LUT_AMPL_WIDTH),
		14930 => to_signed(32449, LUT_AMPL_WIDTH),
		14931 => to_signed(32450, LUT_AMPL_WIDTH),
		14932 => to_signed(32450, LUT_AMPL_WIDTH),
		14933 => to_signed(32450, LUT_AMPL_WIDTH),
		14934 => to_signed(32451, LUT_AMPL_WIDTH),
		14935 => to_signed(32451, LUT_AMPL_WIDTH),
		14936 => to_signed(32452, LUT_AMPL_WIDTH),
		14937 => to_signed(32452, LUT_AMPL_WIDTH),
		14938 => to_signed(32453, LUT_AMPL_WIDTH),
		14939 => to_signed(32453, LUT_AMPL_WIDTH),
		14940 => to_signed(32453, LUT_AMPL_WIDTH),
		14941 => to_signed(32454, LUT_AMPL_WIDTH),
		14942 => to_signed(32454, LUT_AMPL_WIDTH),
		14943 => to_signed(32455, LUT_AMPL_WIDTH),
		14944 => to_signed(32455, LUT_AMPL_WIDTH),
		14945 => to_signed(32456, LUT_AMPL_WIDTH),
		14946 => to_signed(32456, LUT_AMPL_WIDTH),
		14947 => to_signed(32457, LUT_AMPL_WIDTH),
		14948 => to_signed(32457, LUT_AMPL_WIDTH),
		14949 => to_signed(32457, LUT_AMPL_WIDTH),
		14950 => to_signed(32458, LUT_AMPL_WIDTH),
		14951 => to_signed(32458, LUT_AMPL_WIDTH),
		14952 => to_signed(32459, LUT_AMPL_WIDTH),
		14953 => to_signed(32459, LUT_AMPL_WIDTH),
		14954 => to_signed(32460, LUT_AMPL_WIDTH),
		14955 => to_signed(32460, LUT_AMPL_WIDTH),
		14956 => to_signed(32460, LUT_AMPL_WIDTH),
		14957 => to_signed(32461, LUT_AMPL_WIDTH),
		14958 => to_signed(32461, LUT_AMPL_WIDTH),
		14959 => to_signed(32462, LUT_AMPL_WIDTH),
		14960 => to_signed(32462, LUT_AMPL_WIDTH),
		14961 => to_signed(32463, LUT_AMPL_WIDTH),
		14962 => to_signed(32463, LUT_AMPL_WIDTH),
		14963 => to_signed(32463, LUT_AMPL_WIDTH),
		14964 => to_signed(32464, LUT_AMPL_WIDTH),
		14965 => to_signed(32464, LUT_AMPL_WIDTH),
		14966 => to_signed(32465, LUT_AMPL_WIDTH),
		14967 => to_signed(32465, LUT_AMPL_WIDTH),
		14968 => to_signed(32466, LUT_AMPL_WIDTH),
		14969 => to_signed(32466, LUT_AMPL_WIDTH),
		14970 => to_signed(32466, LUT_AMPL_WIDTH),
		14971 => to_signed(32467, LUT_AMPL_WIDTH),
		14972 => to_signed(32467, LUT_AMPL_WIDTH),
		14973 => to_signed(32468, LUT_AMPL_WIDTH),
		14974 => to_signed(32468, LUT_AMPL_WIDTH),
		14975 => to_signed(32468, LUT_AMPL_WIDTH),
		14976 => to_signed(32469, LUT_AMPL_WIDTH),
		14977 => to_signed(32469, LUT_AMPL_WIDTH),
		14978 => to_signed(32470, LUT_AMPL_WIDTH),
		14979 => to_signed(32470, LUT_AMPL_WIDTH),
		14980 => to_signed(32471, LUT_AMPL_WIDTH),
		14981 => to_signed(32471, LUT_AMPL_WIDTH),
		14982 => to_signed(32471, LUT_AMPL_WIDTH),
		14983 => to_signed(32472, LUT_AMPL_WIDTH),
		14984 => to_signed(32472, LUT_AMPL_WIDTH),
		14985 => to_signed(32473, LUT_AMPL_WIDTH),
		14986 => to_signed(32473, LUT_AMPL_WIDTH),
		14987 => to_signed(32474, LUT_AMPL_WIDTH),
		14988 => to_signed(32474, LUT_AMPL_WIDTH),
		14989 => to_signed(32474, LUT_AMPL_WIDTH),
		14990 => to_signed(32475, LUT_AMPL_WIDTH),
		14991 => to_signed(32475, LUT_AMPL_WIDTH),
		14992 => to_signed(32476, LUT_AMPL_WIDTH),
		14993 => to_signed(32476, LUT_AMPL_WIDTH),
		14994 => to_signed(32476, LUT_AMPL_WIDTH),
		14995 => to_signed(32477, LUT_AMPL_WIDTH),
		14996 => to_signed(32477, LUT_AMPL_WIDTH),
		14997 => to_signed(32478, LUT_AMPL_WIDTH),
		14998 => to_signed(32478, LUT_AMPL_WIDTH),
		14999 => to_signed(32479, LUT_AMPL_WIDTH),
		15000 => to_signed(32479, LUT_AMPL_WIDTH),
		15001 => to_signed(32479, LUT_AMPL_WIDTH),
		15002 => to_signed(32480, LUT_AMPL_WIDTH),
		15003 => to_signed(32480, LUT_AMPL_WIDTH),
		15004 => to_signed(32481, LUT_AMPL_WIDTH),
		15005 => to_signed(32481, LUT_AMPL_WIDTH),
		15006 => to_signed(32481, LUT_AMPL_WIDTH),
		15007 => to_signed(32482, LUT_AMPL_WIDTH),
		15008 => to_signed(32482, LUT_AMPL_WIDTH),
		15009 => to_signed(32483, LUT_AMPL_WIDTH),
		15010 => to_signed(32483, LUT_AMPL_WIDTH),
		15011 => to_signed(32484, LUT_AMPL_WIDTH),
		15012 => to_signed(32484, LUT_AMPL_WIDTH),
		15013 => to_signed(32484, LUT_AMPL_WIDTH),
		15014 => to_signed(32485, LUT_AMPL_WIDTH),
		15015 => to_signed(32485, LUT_AMPL_WIDTH),
		15016 => to_signed(32486, LUT_AMPL_WIDTH),
		15017 => to_signed(32486, LUT_AMPL_WIDTH),
		15018 => to_signed(32486, LUT_AMPL_WIDTH),
		15019 => to_signed(32487, LUT_AMPL_WIDTH),
		15020 => to_signed(32487, LUT_AMPL_WIDTH),
		15021 => to_signed(32488, LUT_AMPL_WIDTH),
		15022 => to_signed(32488, LUT_AMPL_WIDTH),
		15023 => to_signed(32488, LUT_AMPL_WIDTH),
		15024 => to_signed(32489, LUT_AMPL_WIDTH),
		15025 => to_signed(32489, LUT_AMPL_WIDTH),
		15026 => to_signed(32490, LUT_AMPL_WIDTH),
		15027 => to_signed(32490, LUT_AMPL_WIDTH),
		15028 => to_signed(32490, LUT_AMPL_WIDTH),
		15029 => to_signed(32491, LUT_AMPL_WIDTH),
		15030 => to_signed(32491, LUT_AMPL_WIDTH),
		15031 => to_signed(32492, LUT_AMPL_WIDTH),
		15032 => to_signed(32492, LUT_AMPL_WIDTH),
		15033 => to_signed(32493, LUT_AMPL_WIDTH),
		15034 => to_signed(32493, LUT_AMPL_WIDTH),
		15035 => to_signed(32493, LUT_AMPL_WIDTH),
		15036 => to_signed(32494, LUT_AMPL_WIDTH),
		15037 => to_signed(32494, LUT_AMPL_WIDTH),
		15038 => to_signed(32495, LUT_AMPL_WIDTH),
		15039 => to_signed(32495, LUT_AMPL_WIDTH),
		15040 => to_signed(32495, LUT_AMPL_WIDTH),
		15041 => to_signed(32496, LUT_AMPL_WIDTH),
		15042 => to_signed(32496, LUT_AMPL_WIDTH),
		15043 => to_signed(32497, LUT_AMPL_WIDTH),
		15044 => to_signed(32497, LUT_AMPL_WIDTH),
		15045 => to_signed(32497, LUT_AMPL_WIDTH),
		15046 => to_signed(32498, LUT_AMPL_WIDTH),
		15047 => to_signed(32498, LUT_AMPL_WIDTH),
		15048 => to_signed(32499, LUT_AMPL_WIDTH),
		15049 => to_signed(32499, LUT_AMPL_WIDTH),
		15050 => to_signed(32499, LUT_AMPL_WIDTH),
		15051 => to_signed(32500, LUT_AMPL_WIDTH),
		15052 => to_signed(32500, LUT_AMPL_WIDTH),
		15053 => to_signed(32501, LUT_AMPL_WIDTH),
		15054 => to_signed(32501, LUT_AMPL_WIDTH),
		15055 => to_signed(32501, LUT_AMPL_WIDTH),
		15056 => to_signed(32502, LUT_AMPL_WIDTH),
		15057 => to_signed(32502, LUT_AMPL_WIDTH),
		15058 => to_signed(32503, LUT_AMPL_WIDTH),
		15059 => to_signed(32503, LUT_AMPL_WIDTH),
		15060 => to_signed(32503, LUT_AMPL_WIDTH),
		15061 => to_signed(32504, LUT_AMPL_WIDTH),
		15062 => to_signed(32504, LUT_AMPL_WIDTH),
		15063 => to_signed(32505, LUT_AMPL_WIDTH),
		15064 => to_signed(32505, LUT_AMPL_WIDTH),
		15065 => to_signed(32505, LUT_AMPL_WIDTH),
		15066 => to_signed(32506, LUT_AMPL_WIDTH),
		15067 => to_signed(32506, LUT_AMPL_WIDTH),
		15068 => to_signed(32507, LUT_AMPL_WIDTH),
		15069 => to_signed(32507, LUT_AMPL_WIDTH),
		15070 => to_signed(32507, LUT_AMPL_WIDTH),
		15071 => to_signed(32508, LUT_AMPL_WIDTH),
		15072 => to_signed(32508, LUT_AMPL_WIDTH),
		15073 => to_signed(32509, LUT_AMPL_WIDTH),
		15074 => to_signed(32509, LUT_AMPL_WIDTH),
		15075 => to_signed(32509, LUT_AMPL_WIDTH),
		15076 => to_signed(32510, LUT_AMPL_WIDTH),
		15077 => to_signed(32510, LUT_AMPL_WIDTH),
		15078 => to_signed(32510, LUT_AMPL_WIDTH),
		15079 => to_signed(32511, LUT_AMPL_WIDTH),
		15080 => to_signed(32511, LUT_AMPL_WIDTH),
		15081 => to_signed(32512, LUT_AMPL_WIDTH),
		15082 => to_signed(32512, LUT_AMPL_WIDTH),
		15083 => to_signed(32512, LUT_AMPL_WIDTH),
		15084 => to_signed(32513, LUT_AMPL_WIDTH),
		15085 => to_signed(32513, LUT_AMPL_WIDTH),
		15086 => to_signed(32514, LUT_AMPL_WIDTH),
		15087 => to_signed(32514, LUT_AMPL_WIDTH),
		15088 => to_signed(32514, LUT_AMPL_WIDTH),
		15089 => to_signed(32515, LUT_AMPL_WIDTH),
		15090 => to_signed(32515, LUT_AMPL_WIDTH),
		15091 => to_signed(32516, LUT_AMPL_WIDTH),
		15092 => to_signed(32516, LUT_AMPL_WIDTH),
		15093 => to_signed(32516, LUT_AMPL_WIDTH),
		15094 => to_signed(32517, LUT_AMPL_WIDTH),
		15095 => to_signed(32517, LUT_AMPL_WIDTH),
		15096 => to_signed(32517, LUT_AMPL_WIDTH),
		15097 => to_signed(32518, LUT_AMPL_WIDTH),
		15098 => to_signed(32518, LUT_AMPL_WIDTH),
		15099 => to_signed(32519, LUT_AMPL_WIDTH),
		15100 => to_signed(32519, LUT_AMPL_WIDTH),
		15101 => to_signed(32519, LUT_AMPL_WIDTH),
		15102 => to_signed(32520, LUT_AMPL_WIDTH),
		15103 => to_signed(32520, LUT_AMPL_WIDTH),
		15104 => to_signed(32521, LUT_AMPL_WIDTH),
		15105 => to_signed(32521, LUT_AMPL_WIDTH),
		15106 => to_signed(32521, LUT_AMPL_WIDTH),
		15107 => to_signed(32522, LUT_AMPL_WIDTH),
		15108 => to_signed(32522, LUT_AMPL_WIDTH),
		15109 => to_signed(32522, LUT_AMPL_WIDTH),
		15110 => to_signed(32523, LUT_AMPL_WIDTH),
		15111 => to_signed(32523, LUT_AMPL_WIDTH),
		15112 => to_signed(32524, LUT_AMPL_WIDTH),
		15113 => to_signed(32524, LUT_AMPL_WIDTH),
		15114 => to_signed(32524, LUT_AMPL_WIDTH),
		15115 => to_signed(32525, LUT_AMPL_WIDTH),
		15116 => to_signed(32525, LUT_AMPL_WIDTH),
		15117 => to_signed(32526, LUT_AMPL_WIDTH),
		15118 => to_signed(32526, LUT_AMPL_WIDTH),
		15119 => to_signed(32526, LUT_AMPL_WIDTH),
		15120 => to_signed(32527, LUT_AMPL_WIDTH),
		15121 => to_signed(32527, LUT_AMPL_WIDTH),
		15122 => to_signed(32527, LUT_AMPL_WIDTH),
		15123 => to_signed(32528, LUT_AMPL_WIDTH),
		15124 => to_signed(32528, LUT_AMPL_WIDTH),
		15125 => to_signed(32529, LUT_AMPL_WIDTH),
		15126 => to_signed(32529, LUT_AMPL_WIDTH),
		15127 => to_signed(32529, LUT_AMPL_WIDTH),
		15128 => to_signed(32530, LUT_AMPL_WIDTH),
		15129 => to_signed(32530, LUT_AMPL_WIDTH),
		15130 => to_signed(32530, LUT_AMPL_WIDTH),
		15131 => to_signed(32531, LUT_AMPL_WIDTH),
		15132 => to_signed(32531, LUT_AMPL_WIDTH),
		15133 => to_signed(32532, LUT_AMPL_WIDTH),
		15134 => to_signed(32532, LUT_AMPL_WIDTH),
		15135 => to_signed(32532, LUT_AMPL_WIDTH),
		15136 => to_signed(32533, LUT_AMPL_WIDTH),
		15137 => to_signed(32533, LUT_AMPL_WIDTH),
		15138 => to_signed(32533, LUT_AMPL_WIDTH),
		15139 => to_signed(32534, LUT_AMPL_WIDTH),
		15140 => to_signed(32534, LUT_AMPL_WIDTH),
		15141 => to_signed(32535, LUT_AMPL_WIDTH),
		15142 => to_signed(32535, LUT_AMPL_WIDTH),
		15143 => to_signed(32535, LUT_AMPL_WIDTH),
		15144 => to_signed(32536, LUT_AMPL_WIDTH),
		15145 => to_signed(32536, LUT_AMPL_WIDTH),
		15146 => to_signed(32536, LUT_AMPL_WIDTH),
		15147 => to_signed(32537, LUT_AMPL_WIDTH),
		15148 => to_signed(32537, LUT_AMPL_WIDTH),
		15149 => to_signed(32538, LUT_AMPL_WIDTH),
		15150 => to_signed(32538, LUT_AMPL_WIDTH),
		15151 => to_signed(32538, LUT_AMPL_WIDTH),
		15152 => to_signed(32539, LUT_AMPL_WIDTH),
		15153 => to_signed(32539, LUT_AMPL_WIDTH),
		15154 => to_signed(32539, LUT_AMPL_WIDTH),
		15155 => to_signed(32540, LUT_AMPL_WIDTH),
		15156 => to_signed(32540, LUT_AMPL_WIDTH),
		15157 => to_signed(32541, LUT_AMPL_WIDTH),
		15158 => to_signed(32541, LUT_AMPL_WIDTH),
		15159 => to_signed(32541, LUT_AMPL_WIDTH),
		15160 => to_signed(32542, LUT_AMPL_WIDTH),
		15161 => to_signed(32542, LUT_AMPL_WIDTH),
		15162 => to_signed(32542, LUT_AMPL_WIDTH),
		15163 => to_signed(32543, LUT_AMPL_WIDTH),
		15164 => to_signed(32543, LUT_AMPL_WIDTH),
		15165 => to_signed(32543, LUT_AMPL_WIDTH),
		15166 => to_signed(32544, LUT_AMPL_WIDTH),
		15167 => to_signed(32544, LUT_AMPL_WIDTH),
		15168 => to_signed(32545, LUT_AMPL_WIDTH),
		15169 => to_signed(32545, LUT_AMPL_WIDTH),
		15170 => to_signed(32545, LUT_AMPL_WIDTH),
		15171 => to_signed(32546, LUT_AMPL_WIDTH),
		15172 => to_signed(32546, LUT_AMPL_WIDTH),
		15173 => to_signed(32546, LUT_AMPL_WIDTH),
		15174 => to_signed(32547, LUT_AMPL_WIDTH),
		15175 => to_signed(32547, LUT_AMPL_WIDTH),
		15176 => to_signed(32547, LUT_AMPL_WIDTH),
		15177 => to_signed(32548, LUT_AMPL_WIDTH),
		15178 => to_signed(32548, LUT_AMPL_WIDTH),
		15179 => to_signed(32549, LUT_AMPL_WIDTH),
		15180 => to_signed(32549, LUT_AMPL_WIDTH),
		15181 => to_signed(32549, LUT_AMPL_WIDTH),
		15182 => to_signed(32550, LUT_AMPL_WIDTH),
		15183 => to_signed(32550, LUT_AMPL_WIDTH),
		15184 => to_signed(32550, LUT_AMPL_WIDTH),
		15185 => to_signed(32551, LUT_AMPL_WIDTH),
		15186 => to_signed(32551, LUT_AMPL_WIDTH),
		15187 => to_signed(32551, LUT_AMPL_WIDTH),
		15188 => to_signed(32552, LUT_AMPL_WIDTH),
		15189 => to_signed(32552, LUT_AMPL_WIDTH),
		15190 => to_signed(32553, LUT_AMPL_WIDTH),
		15191 => to_signed(32553, LUT_AMPL_WIDTH),
		15192 => to_signed(32553, LUT_AMPL_WIDTH),
		15193 => to_signed(32554, LUT_AMPL_WIDTH),
		15194 => to_signed(32554, LUT_AMPL_WIDTH),
		15195 => to_signed(32554, LUT_AMPL_WIDTH),
		15196 => to_signed(32555, LUT_AMPL_WIDTH),
		15197 => to_signed(32555, LUT_AMPL_WIDTH),
		15198 => to_signed(32555, LUT_AMPL_WIDTH),
		15199 => to_signed(32556, LUT_AMPL_WIDTH),
		15200 => to_signed(32556, LUT_AMPL_WIDTH),
		15201 => to_signed(32556, LUT_AMPL_WIDTH),
		15202 => to_signed(32557, LUT_AMPL_WIDTH),
		15203 => to_signed(32557, LUT_AMPL_WIDTH),
		15204 => to_signed(32558, LUT_AMPL_WIDTH),
		15205 => to_signed(32558, LUT_AMPL_WIDTH),
		15206 => to_signed(32558, LUT_AMPL_WIDTH),
		15207 => to_signed(32559, LUT_AMPL_WIDTH),
		15208 => to_signed(32559, LUT_AMPL_WIDTH),
		15209 => to_signed(32559, LUT_AMPL_WIDTH),
		15210 => to_signed(32560, LUT_AMPL_WIDTH),
		15211 => to_signed(32560, LUT_AMPL_WIDTH),
		15212 => to_signed(32560, LUT_AMPL_WIDTH),
		15213 => to_signed(32561, LUT_AMPL_WIDTH),
		15214 => to_signed(32561, LUT_AMPL_WIDTH),
		15215 => to_signed(32561, LUT_AMPL_WIDTH),
		15216 => to_signed(32562, LUT_AMPL_WIDTH),
		15217 => to_signed(32562, LUT_AMPL_WIDTH),
		15218 => to_signed(32562, LUT_AMPL_WIDTH),
		15219 => to_signed(32563, LUT_AMPL_WIDTH),
		15220 => to_signed(32563, LUT_AMPL_WIDTH),
		15221 => to_signed(32564, LUT_AMPL_WIDTH),
		15222 => to_signed(32564, LUT_AMPL_WIDTH),
		15223 => to_signed(32564, LUT_AMPL_WIDTH),
		15224 => to_signed(32565, LUT_AMPL_WIDTH),
		15225 => to_signed(32565, LUT_AMPL_WIDTH),
		15226 => to_signed(32565, LUT_AMPL_WIDTH),
		15227 => to_signed(32566, LUT_AMPL_WIDTH),
		15228 => to_signed(32566, LUT_AMPL_WIDTH),
		15229 => to_signed(32566, LUT_AMPL_WIDTH),
		15230 => to_signed(32567, LUT_AMPL_WIDTH),
		15231 => to_signed(32567, LUT_AMPL_WIDTH),
		15232 => to_signed(32567, LUT_AMPL_WIDTH),
		15233 => to_signed(32568, LUT_AMPL_WIDTH),
		15234 => to_signed(32568, LUT_AMPL_WIDTH),
		15235 => to_signed(32568, LUT_AMPL_WIDTH),
		15236 => to_signed(32569, LUT_AMPL_WIDTH),
		15237 => to_signed(32569, LUT_AMPL_WIDTH),
		15238 => to_signed(32569, LUT_AMPL_WIDTH),
		15239 => to_signed(32570, LUT_AMPL_WIDTH),
		15240 => to_signed(32570, LUT_AMPL_WIDTH),
		15241 => to_signed(32570, LUT_AMPL_WIDTH),
		15242 => to_signed(32571, LUT_AMPL_WIDTH),
		15243 => to_signed(32571, LUT_AMPL_WIDTH),
		15244 => to_signed(32571, LUT_AMPL_WIDTH),
		15245 => to_signed(32572, LUT_AMPL_WIDTH),
		15246 => to_signed(32572, LUT_AMPL_WIDTH),
		15247 => to_signed(32573, LUT_AMPL_WIDTH),
		15248 => to_signed(32573, LUT_AMPL_WIDTH),
		15249 => to_signed(32573, LUT_AMPL_WIDTH),
		15250 => to_signed(32574, LUT_AMPL_WIDTH),
		15251 => to_signed(32574, LUT_AMPL_WIDTH),
		15252 => to_signed(32574, LUT_AMPL_WIDTH),
		15253 => to_signed(32575, LUT_AMPL_WIDTH),
		15254 => to_signed(32575, LUT_AMPL_WIDTH),
		15255 => to_signed(32575, LUT_AMPL_WIDTH),
		15256 => to_signed(32576, LUT_AMPL_WIDTH),
		15257 => to_signed(32576, LUT_AMPL_WIDTH),
		15258 => to_signed(32576, LUT_AMPL_WIDTH),
		15259 => to_signed(32577, LUT_AMPL_WIDTH),
		15260 => to_signed(32577, LUT_AMPL_WIDTH),
		15261 => to_signed(32577, LUT_AMPL_WIDTH),
		15262 => to_signed(32578, LUT_AMPL_WIDTH),
		15263 => to_signed(32578, LUT_AMPL_WIDTH),
		15264 => to_signed(32578, LUT_AMPL_WIDTH),
		15265 => to_signed(32579, LUT_AMPL_WIDTH),
		15266 => to_signed(32579, LUT_AMPL_WIDTH),
		15267 => to_signed(32579, LUT_AMPL_WIDTH),
		15268 => to_signed(32580, LUT_AMPL_WIDTH),
		15269 => to_signed(32580, LUT_AMPL_WIDTH),
		15270 => to_signed(32580, LUT_AMPL_WIDTH),
		15271 => to_signed(32581, LUT_AMPL_WIDTH),
		15272 => to_signed(32581, LUT_AMPL_WIDTH),
		15273 => to_signed(32581, LUT_AMPL_WIDTH),
		15274 => to_signed(32582, LUT_AMPL_WIDTH),
		15275 => to_signed(32582, LUT_AMPL_WIDTH),
		15276 => to_signed(32582, LUT_AMPL_WIDTH),
		15277 => to_signed(32583, LUT_AMPL_WIDTH),
		15278 => to_signed(32583, LUT_AMPL_WIDTH),
		15279 => to_signed(32583, LUT_AMPL_WIDTH),
		15280 => to_signed(32584, LUT_AMPL_WIDTH),
		15281 => to_signed(32584, LUT_AMPL_WIDTH),
		15282 => to_signed(32584, LUT_AMPL_WIDTH),
		15283 => to_signed(32585, LUT_AMPL_WIDTH),
		15284 => to_signed(32585, LUT_AMPL_WIDTH),
		15285 => to_signed(32585, LUT_AMPL_WIDTH),
		15286 => to_signed(32586, LUT_AMPL_WIDTH),
		15287 => to_signed(32586, LUT_AMPL_WIDTH),
		15288 => to_signed(32586, LUT_AMPL_WIDTH),
		15289 => to_signed(32587, LUT_AMPL_WIDTH),
		15290 => to_signed(32587, LUT_AMPL_WIDTH),
		15291 => to_signed(32587, LUT_AMPL_WIDTH),
		15292 => to_signed(32588, LUT_AMPL_WIDTH),
		15293 => to_signed(32588, LUT_AMPL_WIDTH),
		15294 => to_signed(32588, LUT_AMPL_WIDTH),
		15295 => to_signed(32589, LUT_AMPL_WIDTH),
		15296 => to_signed(32589, LUT_AMPL_WIDTH),
		15297 => to_signed(32589, LUT_AMPL_WIDTH),
		15298 => to_signed(32590, LUT_AMPL_WIDTH),
		15299 => to_signed(32590, LUT_AMPL_WIDTH),
		15300 => to_signed(32590, LUT_AMPL_WIDTH),
		15301 => to_signed(32591, LUT_AMPL_WIDTH),
		15302 => to_signed(32591, LUT_AMPL_WIDTH),
		15303 => to_signed(32591, LUT_AMPL_WIDTH),
		15304 => to_signed(32592, LUT_AMPL_WIDTH),
		15305 => to_signed(32592, LUT_AMPL_WIDTH),
		15306 => to_signed(32592, LUT_AMPL_WIDTH),
		15307 => to_signed(32592, LUT_AMPL_WIDTH),
		15308 => to_signed(32593, LUT_AMPL_WIDTH),
		15309 => to_signed(32593, LUT_AMPL_WIDTH),
		15310 => to_signed(32593, LUT_AMPL_WIDTH),
		15311 => to_signed(32594, LUT_AMPL_WIDTH),
		15312 => to_signed(32594, LUT_AMPL_WIDTH),
		15313 => to_signed(32594, LUT_AMPL_WIDTH),
		15314 => to_signed(32595, LUT_AMPL_WIDTH),
		15315 => to_signed(32595, LUT_AMPL_WIDTH),
		15316 => to_signed(32595, LUT_AMPL_WIDTH),
		15317 => to_signed(32596, LUT_AMPL_WIDTH),
		15318 => to_signed(32596, LUT_AMPL_WIDTH),
		15319 => to_signed(32596, LUT_AMPL_WIDTH),
		15320 => to_signed(32597, LUT_AMPL_WIDTH),
		15321 => to_signed(32597, LUT_AMPL_WIDTH),
		15322 => to_signed(32597, LUT_AMPL_WIDTH),
		15323 => to_signed(32598, LUT_AMPL_WIDTH),
		15324 => to_signed(32598, LUT_AMPL_WIDTH),
		15325 => to_signed(32598, LUT_AMPL_WIDTH),
		15326 => to_signed(32599, LUT_AMPL_WIDTH),
		15327 => to_signed(32599, LUT_AMPL_WIDTH),
		15328 => to_signed(32599, LUT_AMPL_WIDTH),
		15329 => to_signed(32600, LUT_AMPL_WIDTH),
		15330 => to_signed(32600, LUT_AMPL_WIDTH),
		15331 => to_signed(32600, LUT_AMPL_WIDTH),
		15332 => to_signed(32600, LUT_AMPL_WIDTH),
		15333 => to_signed(32601, LUT_AMPL_WIDTH),
		15334 => to_signed(32601, LUT_AMPL_WIDTH),
		15335 => to_signed(32601, LUT_AMPL_WIDTH),
		15336 => to_signed(32602, LUT_AMPL_WIDTH),
		15337 => to_signed(32602, LUT_AMPL_WIDTH),
		15338 => to_signed(32602, LUT_AMPL_WIDTH),
		15339 => to_signed(32603, LUT_AMPL_WIDTH),
		15340 => to_signed(32603, LUT_AMPL_WIDTH),
		15341 => to_signed(32603, LUT_AMPL_WIDTH),
		15342 => to_signed(32604, LUT_AMPL_WIDTH),
		15343 => to_signed(32604, LUT_AMPL_WIDTH),
		15344 => to_signed(32604, LUT_AMPL_WIDTH),
		15345 => to_signed(32605, LUT_AMPL_WIDTH),
		15346 => to_signed(32605, LUT_AMPL_WIDTH),
		15347 => to_signed(32605, LUT_AMPL_WIDTH),
		15348 => to_signed(32606, LUT_AMPL_WIDTH),
		15349 => to_signed(32606, LUT_AMPL_WIDTH),
		15350 => to_signed(32606, LUT_AMPL_WIDTH),
		15351 => to_signed(32606, LUT_AMPL_WIDTH),
		15352 => to_signed(32607, LUT_AMPL_WIDTH),
		15353 => to_signed(32607, LUT_AMPL_WIDTH),
		15354 => to_signed(32607, LUT_AMPL_WIDTH),
		15355 => to_signed(32608, LUT_AMPL_WIDTH),
		15356 => to_signed(32608, LUT_AMPL_WIDTH),
		15357 => to_signed(32608, LUT_AMPL_WIDTH),
		15358 => to_signed(32609, LUT_AMPL_WIDTH),
		15359 => to_signed(32609, LUT_AMPL_WIDTH),
		15360 => to_signed(32609, LUT_AMPL_WIDTH),
		15361 => to_signed(32610, LUT_AMPL_WIDTH),
		15362 => to_signed(32610, LUT_AMPL_WIDTH),
		15363 => to_signed(32610, LUT_AMPL_WIDTH),
		15364 => to_signed(32610, LUT_AMPL_WIDTH),
		15365 => to_signed(32611, LUT_AMPL_WIDTH),
		15366 => to_signed(32611, LUT_AMPL_WIDTH),
		15367 => to_signed(32611, LUT_AMPL_WIDTH),
		15368 => to_signed(32612, LUT_AMPL_WIDTH),
		15369 => to_signed(32612, LUT_AMPL_WIDTH),
		15370 => to_signed(32612, LUT_AMPL_WIDTH),
		15371 => to_signed(32613, LUT_AMPL_WIDTH),
		15372 => to_signed(32613, LUT_AMPL_WIDTH),
		15373 => to_signed(32613, LUT_AMPL_WIDTH),
		15374 => to_signed(32613, LUT_AMPL_WIDTH),
		15375 => to_signed(32614, LUT_AMPL_WIDTH),
		15376 => to_signed(32614, LUT_AMPL_WIDTH),
		15377 => to_signed(32614, LUT_AMPL_WIDTH),
		15378 => to_signed(32615, LUT_AMPL_WIDTH),
		15379 => to_signed(32615, LUT_AMPL_WIDTH),
		15380 => to_signed(32615, LUT_AMPL_WIDTH),
		15381 => to_signed(32616, LUT_AMPL_WIDTH),
		15382 => to_signed(32616, LUT_AMPL_WIDTH),
		15383 => to_signed(32616, LUT_AMPL_WIDTH),
		15384 => to_signed(32617, LUT_AMPL_WIDTH),
		15385 => to_signed(32617, LUT_AMPL_WIDTH),
		15386 => to_signed(32617, LUT_AMPL_WIDTH),
		15387 => to_signed(32617, LUT_AMPL_WIDTH),
		15388 => to_signed(32618, LUT_AMPL_WIDTH),
		15389 => to_signed(32618, LUT_AMPL_WIDTH),
		15390 => to_signed(32618, LUT_AMPL_WIDTH),
		15391 => to_signed(32619, LUT_AMPL_WIDTH),
		15392 => to_signed(32619, LUT_AMPL_WIDTH),
		15393 => to_signed(32619, LUT_AMPL_WIDTH),
		15394 => to_signed(32620, LUT_AMPL_WIDTH),
		15395 => to_signed(32620, LUT_AMPL_WIDTH),
		15396 => to_signed(32620, LUT_AMPL_WIDTH),
		15397 => to_signed(32620, LUT_AMPL_WIDTH),
		15398 => to_signed(32621, LUT_AMPL_WIDTH),
		15399 => to_signed(32621, LUT_AMPL_WIDTH),
		15400 => to_signed(32621, LUT_AMPL_WIDTH),
		15401 => to_signed(32622, LUT_AMPL_WIDTH),
		15402 => to_signed(32622, LUT_AMPL_WIDTH),
		15403 => to_signed(32622, LUT_AMPL_WIDTH),
		15404 => to_signed(32622, LUT_AMPL_WIDTH),
		15405 => to_signed(32623, LUT_AMPL_WIDTH),
		15406 => to_signed(32623, LUT_AMPL_WIDTH),
		15407 => to_signed(32623, LUT_AMPL_WIDTH),
		15408 => to_signed(32624, LUT_AMPL_WIDTH),
		15409 => to_signed(32624, LUT_AMPL_WIDTH),
		15410 => to_signed(32624, LUT_AMPL_WIDTH),
		15411 => to_signed(32625, LUT_AMPL_WIDTH),
		15412 => to_signed(32625, LUT_AMPL_WIDTH),
		15413 => to_signed(32625, LUT_AMPL_WIDTH),
		15414 => to_signed(32625, LUT_AMPL_WIDTH),
		15415 => to_signed(32626, LUT_AMPL_WIDTH),
		15416 => to_signed(32626, LUT_AMPL_WIDTH),
		15417 => to_signed(32626, LUT_AMPL_WIDTH),
		15418 => to_signed(32627, LUT_AMPL_WIDTH),
		15419 => to_signed(32627, LUT_AMPL_WIDTH),
		15420 => to_signed(32627, LUT_AMPL_WIDTH),
		15421 => to_signed(32627, LUT_AMPL_WIDTH),
		15422 => to_signed(32628, LUT_AMPL_WIDTH),
		15423 => to_signed(32628, LUT_AMPL_WIDTH),
		15424 => to_signed(32628, LUT_AMPL_WIDTH),
		15425 => to_signed(32629, LUT_AMPL_WIDTH),
		15426 => to_signed(32629, LUT_AMPL_WIDTH),
		15427 => to_signed(32629, LUT_AMPL_WIDTH),
		15428 => to_signed(32629, LUT_AMPL_WIDTH),
		15429 => to_signed(32630, LUT_AMPL_WIDTH),
		15430 => to_signed(32630, LUT_AMPL_WIDTH),
		15431 => to_signed(32630, LUT_AMPL_WIDTH),
		15432 => to_signed(32631, LUT_AMPL_WIDTH),
		15433 => to_signed(32631, LUT_AMPL_WIDTH),
		15434 => to_signed(32631, LUT_AMPL_WIDTH),
		15435 => to_signed(32631, LUT_AMPL_WIDTH),
		15436 => to_signed(32632, LUT_AMPL_WIDTH),
		15437 => to_signed(32632, LUT_AMPL_WIDTH),
		15438 => to_signed(32632, LUT_AMPL_WIDTH),
		15439 => to_signed(32633, LUT_AMPL_WIDTH),
		15440 => to_signed(32633, LUT_AMPL_WIDTH),
		15441 => to_signed(32633, LUT_AMPL_WIDTH),
		15442 => to_signed(32633, LUT_AMPL_WIDTH),
		15443 => to_signed(32634, LUT_AMPL_WIDTH),
		15444 => to_signed(32634, LUT_AMPL_WIDTH),
		15445 => to_signed(32634, LUT_AMPL_WIDTH),
		15446 => to_signed(32635, LUT_AMPL_WIDTH),
		15447 => to_signed(32635, LUT_AMPL_WIDTH),
		15448 => to_signed(32635, LUT_AMPL_WIDTH),
		15449 => to_signed(32635, LUT_AMPL_WIDTH),
		15450 => to_signed(32636, LUT_AMPL_WIDTH),
		15451 => to_signed(32636, LUT_AMPL_WIDTH),
		15452 => to_signed(32636, LUT_AMPL_WIDTH),
		15453 => to_signed(32637, LUT_AMPL_WIDTH),
		15454 => to_signed(32637, LUT_AMPL_WIDTH),
		15455 => to_signed(32637, LUT_AMPL_WIDTH),
		15456 => to_signed(32637, LUT_AMPL_WIDTH),
		15457 => to_signed(32638, LUT_AMPL_WIDTH),
		15458 => to_signed(32638, LUT_AMPL_WIDTH),
		15459 => to_signed(32638, LUT_AMPL_WIDTH),
		15460 => to_signed(32639, LUT_AMPL_WIDTH),
		15461 => to_signed(32639, LUT_AMPL_WIDTH),
		15462 => to_signed(32639, LUT_AMPL_WIDTH),
		15463 => to_signed(32639, LUT_AMPL_WIDTH),
		15464 => to_signed(32640, LUT_AMPL_WIDTH),
		15465 => to_signed(32640, LUT_AMPL_WIDTH),
		15466 => to_signed(32640, LUT_AMPL_WIDTH),
		15467 => to_signed(32640, LUT_AMPL_WIDTH),
		15468 => to_signed(32641, LUT_AMPL_WIDTH),
		15469 => to_signed(32641, LUT_AMPL_WIDTH),
		15470 => to_signed(32641, LUT_AMPL_WIDTH),
		15471 => to_signed(32642, LUT_AMPL_WIDTH),
		15472 => to_signed(32642, LUT_AMPL_WIDTH),
		15473 => to_signed(32642, LUT_AMPL_WIDTH),
		15474 => to_signed(32642, LUT_AMPL_WIDTH),
		15475 => to_signed(32643, LUT_AMPL_WIDTH),
		15476 => to_signed(32643, LUT_AMPL_WIDTH),
		15477 => to_signed(32643, LUT_AMPL_WIDTH),
		15478 => to_signed(32643, LUT_AMPL_WIDTH),
		15479 => to_signed(32644, LUT_AMPL_WIDTH),
		15480 => to_signed(32644, LUT_AMPL_WIDTH),
		15481 => to_signed(32644, LUT_AMPL_WIDTH),
		15482 => to_signed(32645, LUT_AMPL_WIDTH),
		15483 => to_signed(32645, LUT_AMPL_WIDTH),
		15484 => to_signed(32645, LUT_AMPL_WIDTH),
		15485 => to_signed(32645, LUT_AMPL_WIDTH),
		15486 => to_signed(32646, LUT_AMPL_WIDTH),
		15487 => to_signed(32646, LUT_AMPL_WIDTH),
		15488 => to_signed(32646, LUT_AMPL_WIDTH),
		15489 => to_signed(32646, LUT_AMPL_WIDTH),
		15490 => to_signed(32647, LUT_AMPL_WIDTH),
		15491 => to_signed(32647, LUT_AMPL_WIDTH),
		15492 => to_signed(32647, LUT_AMPL_WIDTH),
		15493 => to_signed(32648, LUT_AMPL_WIDTH),
		15494 => to_signed(32648, LUT_AMPL_WIDTH),
		15495 => to_signed(32648, LUT_AMPL_WIDTH),
		15496 => to_signed(32648, LUT_AMPL_WIDTH),
		15497 => to_signed(32649, LUT_AMPL_WIDTH),
		15498 => to_signed(32649, LUT_AMPL_WIDTH),
		15499 => to_signed(32649, LUT_AMPL_WIDTH),
		15500 => to_signed(32649, LUT_AMPL_WIDTH),
		15501 => to_signed(32650, LUT_AMPL_WIDTH),
		15502 => to_signed(32650, LUT_AMPL_WIDTH),
		15503 => to_signed(32650, LUT_AMPL_WIDTH),
		15504 => to_signed(32650, LUT_AMPL_WIDTH),
		15505 => to_signed(32651, LUT_AMPL_WIDTH),
		15506 => to_signed(32651, LUT_AMPL_WIDTH),
		15507 => to_signed(32651, LUT_AMPL_WIDTH),
		15508 => to_signed(32652, LUT_AMPL_WIDTH),
		15509 => to_signed(32652, LUT_AMPL_WIDTH),
		15510 => to_signed(32652, LUT_AMPL_WIDTH),
		15511 => to_signed(32652, LUT_AMPL_WIDTH),
		15512 => to_signed(32653, LUT_AMPL_WIDTH),
		15513 => to_signed(32653, LUT_AMPL_WIDTH),
		15514 => to_signed(32653, LUT_AMPL_WIDTH),
		15515 => to_signed(32653, LUT_AMPL_WIDTH),
		15516 => to_signed(32654, LUT_AMPL_WIDTH),
		15517 => to_signed(32654, LUT_AMPL_WIDTH),
		15518 => to_signed(32654, LUT_AMPL_WIDTH),
		15519 => to_signed(32654, LUT_AMPL_WIDTH),
		15520 => to_signed(32655, LUT_AMPL_WIDTH),
		15521 => to_signed(32655, LUT_AMPL_WIDTH),
		15522 => to_signed(32655, LUT_AMPL_WIDTH),
		15523 => to_signed(32655, LUT_AMPL_WIDTH),
		15524 => to_signed(32656, LUT_AMPL_WIDTH),
		15525 => to_signed(32656, LUT_AMPL_WIDTH),
		15526 => to_signed(32656, LUT_AMPL_WIDTH),
		15527 => to_signed(32656, LUT_AMPL_WIDTH),
		15528 => to_signed(32657, LUT_AMPL_WIDTH),
		15529 => to_signed(32657, LUT_AMPL_WIDTH),
		15530 => to_signed(32657, LUT_AMPL_WIDTH),
		15531 => to_signed(32657, LUT_AMPL_WIDTH),
		15532 => to_signed(32658, LUT_AMPL_WIDTH),
		15533 => to_signed(32658, LUT_AMPL_WIDTH),
		15534 => to_signed(32658, LUT_AMPL_WIDTH),
		15535 => to_signed(32659, LUT_AMPL_WIDTH),
		15536 => to_signed(32659, LUT_AMPL_WIDTH),
		15537 => to_signed(32659, LUT_AMPL_WIDTH),
		15538 => to_signed(32659, LUT_AMPL_WIDTH),
		15539 => to_signed(32660, LUT_AMPL_WIDTH),
		15540 => to_signed(32660, LUT_AMPL_WIDTH),
		15541 => to_signed(32660, LUT_AMPL_WIDTH),
		15542 => to_signed(32660, LUT_AMPL_WIDTH),
		15543 => to_signed(32661, LUT_AMPL_WIDTH),
		15544 => to_signed(32661, LUT_AMPL_WIDTH),
		15545 => to_signed(32661, LUT_AMPL_WIDTH),
		15546 => to_signed(32661, LUT_AMPL_WIDTH),
		15547 => to_signed(32662, LUT_AMPL_WIDTH),
		15548 => to_signed(32662, LUT_AMPL_WIDTH),
		15549 => to_signed(32662, LUT_AMPL_WIDTH),
		15550 => to_signed(32662, LUT_AMPL_WIDTH),
		15551 => to_signed(32663, LUT_AMPL_WIDTH),
		15552 => to_signed(32663, LUT_AMPL_WIDTH),
		15553 => to_signed(32663, LUT_AMPL_WIDTH),
		15554 => to_signed(32663, LUT_AMPL_WIDTH),
		15555 => to_signed(32664, LUT_AMPL_WIDTH),
		15556 => to_signed(32664, LUT_AMPL_WIDTH),
		15557 => to_signed(32664, LUT_AMPL_WIDTH),
		15558 => to_signed(32664, LUT_AMPL_WIDTH),
		15559 => to_signed(32665, LUT_AMPL_WIDTH),
		15560 => to_signed(32665, LUT_AMPL_WIDTH),
		15561 => to_signed(32665, LUT_AMPL_WIDTH),
		15562 => to_signed(32665, LUT_AMPL_WIDTH),
		15563 => to_signed(32666, LUT_AMPL_WIDTH),
		15564 => to_signed(32666, LUT_AMPL_WIDTH),
		15565 => to_signed(32666, LUT_AMPL_WIDTH),
		15566 => to_signed(32666, LUT_AMPL_WIDTH),
		15567 => to_signed(32667, LUT_AMPL_WIDTH),
		15568 => to_signed(32667, LUT_AMPL_WIDTH),
		15569 => to_signed(32667, LUT_AMPL_WIDTH),
		15570 => to_signed(32667, LUT_AMPL_WIDTH),
		15571 => to_signed(32668, LUT_AMPL_WIDTH),
		15572 => to_signed(32668, LUT_AMPL_WIDTH),
		15573 => to_signed(32668, LUT_AMPL_WIDTH),
		15574 => to_signed(32668, LUT_AMPL_WIDTH),
		15575 => to_signed(32668, LUT_AMPL_WIDTH),
		15576 => to_signed(32669, LUT_AMPL_WIDTH),
		15577 => to_signed(32669, LUT_AMPL_WIDTH),
		15578 => to_signed(32669, LUT_AMPL_WIDTH),
		15579 => to_signed(32669, LUT_AMPL_WIDTH),
		15580 => to_signed(32670, LUT_AMPL_WIDTH),
		15581 => to_signed(32670, LUT_AMPL_WIDTH),
		15582 => to_signed(32670, LUT_AMPL_WIDTH),
		15583 => to_signed(32670, LUT_AMPL_WIDTH),
		15584 => to_signed(32671, LUT_AMPL_WIDTH),
		15585 => to_signed(32671, LUT_AMPL_WIDTH),
		15586 => to_signed(32671, LUT_AMPL_WIDTH),
		15587 => to_signed(32671, LUT_AMPL_WIDTH),
		15588 => to_signed(32672, LUT_AMPL_WIDTH),
		15589 => to_signed(32672, LUT_AMPL_WIDTH),
		15590 => to_signed(32672, LUT_AMPL_WIDTH),
		15591 => to_signed(32672, LUT_AMPL_WIDTH),
		15592 => to_signed(32673, LUT_AMPL_WIDTH),
		15593 => to_signed(32673, LUT_AMPL_WIDTH),
		15594 => to_signed(32673, LUT_AMPL_WIDTH),
		15595 => to_signed(32673, LUT_AMPL_WIDTH),
		15596 => to_signed(32674, LUT_AMPL_WIDTH),
		15597 => to_signed(32674, LUT_AMPL_WIDTH),
		15598 => to_signed(32674, LUT_AMPL_WIDTH),
		15599 => to_signed(32674, LUT_AMPL_WIDTH),
		15600 => to_signed(32674, LUT_AMPL_WIDTH),
		15601 => to_signed(32675, LUT_AMPL_WIDTH),
		15602 => to_signed(32675, LUT_AMPL_WIDTH),
		15603 => to_signed(32675, LUT_AMPL_WIDTH),
		15604 => to_signed(32675, LUT_AMPL_WIDTH),
		15605 => to_signed(32676, LUT_AMPL_WIDTH),
		15606 => to_signed(32676, LUT_AMPL_WIDTH),
		15607 => to_signed(32676, LUT_AMPL_WIDTH),
		15608 => to_signed(32676, LUT_AMPL_WIDTH),
		15609 => to_signed(32677, LUT_AMPL_WIDTH),
		15610 => to_signed(32677, LUT_AMPL_WIDTH),
		15611 => to_signed(32677, LUT_AMPL_WIDTH),
		15612 => to_signed(32677, LUT_AMPL_WIDTH),
		15613 => to_signed(32678, LUT_AMPL_WIDTH),
		15614 => to_signed(32678, LUT_AMPL_WIDTH),
		15615 => to_signed(32678, LUT_AMPL_WIDTH),
		15616 => to_signed(32678, LUT_AMPL_WIDTH),
		15617 => to_signed(32678, LUT_AMPL_WIDTH),
		15618 => to_signed(32679, LUT_AMPL_WIDTH),
		15619 => to_signed(32679, LUT_AMPL_WIDTH),
		15620 => to_signed(32679, LUT_AMPL_WIDTH),
		15621 => to_signed(32679, LUT_AMPL_WIDTH),
		15622 => to_signed(32680, LUT_AMPL_WIDTH),
		15623 => to_signed(32680, LUT_AMPL_WIDTH),
		15624 => to_signed(32680, LUT_AMPL_WIDTH),
		15625 => to_signed(32680, LUT_AMPL_WIDTH),
		15626 => to_signed(32681, LUT_AMPL_WIDTH),
		15627 => to_signed(32681, LUT_AMPL_WIDTH),
		15628 => to_signed(32681, LUT_AMPL_WIDTH),
		15629 => to_signed(32681, LUT_AMPL_WIDTH),
		15630 => to_signed(32681, LUT_AMPL_WIDTH),
		15631 => to_signed(32682, LUT_AMPL_WIDTH),
		15632 => to_signed(32682, LUT_AMPL_WIDTH),
		15633 => to_signed(32682, LUT_AMPL_WIDTH),
		15634 => to_signed(32682, LUT_AMPL_WIDTH),
		15635 => to_signed(32683, LUT_AMPL_WIDTH),
		15636 => to_signed(32683, LUT_AMPL_WIDTH),
		15637 => to_signed(32683, LUT_AMPL_WIDTH),
		15638 => to_signed(32683, LUT_AMPL_WIDTH),
		15639 => to_signed(32683, LUT_AMPL_WIDTH),
		15640 => to_signed(32684, LUT_AMPL_WIDTH),
		15641 => to_signed(32684, LUT_AMPL_WIDTH),
		15642 => to_signed(32684, LUT_AMPL_WIDTH),
		15643 => to_signed(32684, LUT_AMPL_WIDTH),
		15644 => to_signed(32685, LUT_AMPL_WIDTH),
		15645 => to_signed(32685, LUT_AMPL_WIDTH),
		15646 => to_signed(32685, LUT_AMPL_WIDTH),
		15647 => to_signed(32685, LUT_AMPL_WIDTH),
		15648 => to_signed(32685, LUT_AMPL_WIDTH),
		15649 => to_signed(32686, LUT_AMPL_WIDTH),
		15650 => to_signed(32686, LUT_AMPL_WIDTH),
		15651 => to_signed(32686, LUT_AMPL_WIDTH),
		15652 => to_signed(32686, LUT_AMPL_WIDTH),
		15653 => to_signed(32687, LUT_AMPL_WIDTH),
		15654 => to_signed(32687, LUT_AMPL_WIDTH),
		15655 => to_signed(32687, LUT_AMPL_WIDTH),
		15656 => to_signed(32687, LUT_AMPL_WIDTH),
		15657 => to_signed(32687, LUT_AMPL_WIDTH),
		15658 => to_signed(32688, LUT_AMPL_WIDTH),
		15659 => to_signed(32688, LUT_AMPL_WIDTH),
		15660 => to_signed(32688, LUT_AMPL_WIDTH),
		15661 => to_signed(32688, LUT_AMPL_WIDTH),
		15662 => to_signed(32689, LUT_AMPL_WIDTH),
		15663 => to_signed(32689, LUT_AMPL_WIDTH),
		15664 => to_signed(32689, LUT_AMPL_WIDTH),
		15665 => to_signed(32689, LUT_AMPL_WIDTH),
		15666 => to_signed(32689, LUT_AMPL_WIDTH),
		15667 => to_signed(32690, LUT_AMPL_WIDTH),
		15668 => to_signed(32690, LUT_AMPL_WIDTH),
		15669 => to_signed(32690, LUT_AMPL_WIDTH),
		15670 => to_signed(32690, LUT_AMPL_WIDTH),
		15671 => to_signed(32690, LUT_AMPL_WIDTH),
		15672 => to_signed(32691, LUT_AMPL_WIDTH),
		15673 => to_signed(32691, LUT_AMPL_WIDTH),
		15674 => to_signed(32691, LUT_AMPL_WIDTH),
		15675 => to_signed(32691, LUT_AMPL_WIDTH),
		15676 => to_signed(32692, LUT_AMPL_WIDTH),
		15677 => to_signed(32692, LUT_AMPL_WIDTH),
		15678 => to_signed(32692, LUT_AMPL_WIDTH),
		15679 => to_signed(32692, LUT_AMPL_WIDTH),
		15680 => to_signed(32692, LUT_AMPL_WIDTH),
		15681 => to_signed(32693, LUT_AMPL_WIDTH),
		15682 => to_signed(32693, LUT_AMPL_WIDTH),
		15683 => to_signed(32693, LUT_AMPL_WIDTH),
		15684 => to_signed(32693, LUT_AMPL_WIDTH),
		15685 => to_signed(32693, LUT_AMPL_WIDTH),
		15686 => to_signed(32694, LUT_AMPL_WIDTH),
		15687 => to_signed(32694, LUT_AMPL_WIDTH),
		15688 => to_signed(32694, LUT_AMPL_WIDTH),
		15689 => to_signed(32694, LUT_AMPL_WIDTH),
		15690 => to_signed(32694, LUT_AMPL_WIDTH),
		15691 => to_signed(32695, LUT_AMPL_WIDTH),
		15692 => to_signed(32695, LUT_AMPL_WIDTH),
		15693 => to_signed(32695, LUT_AMPL_WIDTH),
		15694 => to_signed(32695, LUT_AMPL_WIDTH),
		15695 => to_signed(32696, LUT_AMPL_WIDTH),
		15696 => to_signed(32696, LUT_AMPL_WIDTH),
		15697 => to_signed(32696, LUT_AMPL_WIDTH),
		15698 => to_signed(32696, LUT_AMPL_WIDTH),
		15699 => to_signed(32696, LUT_AMPL_WIDTH),
		15700 => to_signed(32697, LUT_AMPL_WIDTH),
		15701 => to_signed(32697, LUT_AMPL_WIDTH),
		15702 => to_signed(32697, LUT_AMPL_WIDTH),
		15703 => to_signed(32697, LUT_AMPL_WIDTH),
		15704 => to_signed(32697, LUT_AMPL_WIDTH),
		15705 => to_signed(32698, LUT_AMPL_WIDTH),
		15706 => to_signed(32698, LUT_AMPL_WIDTH),
		15707 => to_signed(32698, LUT_AMPL_WIDTH),
		15708 => to_signed(32698, LUT_AMPL_WIDTH),
		15709 => to_signed(32698, LUT_AMPL_WIDTH),
		15710 => to_signed(32699, LUT_AMPL_WIDTH),
		15711 => to_signed(32699, LUT_AMPL_WIDTH),
		15712 => to_signed(32699, LUT_AMPL_WIDTH),
		15713 => to_signed(32699, LUT_AMPL_WIDTH),
		15714 => to_signed(32699, LUT_AMPL_WIDTH),
		15715 => to_signed(32700, LUT_AMPL_WIDTH),
		15716 => to_signed(32700, LUT_AMPL_WIDTH),
		15717 => to_signed(32700, LUT_AMPL_WIDTH),
		15718 => to_signed(32700, LUT_AMPL_WIDTH),
		15719 => to_signed(32700, LUT_AMPL_WIDTH),
		15720 => to_signed(32701, LUT_AMPL_WIDTH),
		15721 => to_signed(32701, LUT_AMPL_WIDTH),
		15722 => to_signed(32701, LUT_AMPL_WIDTH),
		15723 => to_signed(32701, LUT_AMPL_WIDTH),
		15724 => to_signed(32701, LUT_AMPL_WIDTH),
		15725 => to_signed(32702, LUT_AMPL_WIDTH),
		15726 => to_signed(32702, LUT_AMPL_WIDTH),
		15727 => to_signed(32702, LUT_AMPL_WIDTH),
		15728 => to_signed(32702, LUT_AMPL_WIDTH),
		15729 => to_signed(32702, LUT_AMPL_WIDTH),
		15730 => to_signed(32703, LUT_AMPL_WIDTH),
		15731 => to_signed(32703, LUT_AMPL_WIDTH),
		15732 => to_signed(32703, LUT_AMPL_WIDTH),
		15733 => to_signed(32703, LUT_AMPL_WIDTH),
		15734 => to_signed(32703, LUT_AMPL_WIDTH),
		15735 => to_signed(32704, LUT_AMPL_WIDTH),
		15736 => to_signed(32704, LUT_AMPL_WIDTH),
		15737 => to_signed(32704, LUT_AMPL_WIDTH),
		15738 => to_signed(32704, LUT_AMPL_WIDTH),
		15739 => to_signed(32704, LUT_AMPL_WIDTH),
		15740 => to_signed(32705, LUT_AMPL_WIDTH),
		15741 => to_signed(32705, LUT_AMPL_WIDTH),
		15742 => to_signed(32705, LUT_AMPL_WIDTH),
		15743 => to_signed(32705, LUT_AMPL_WIDTH),
		15744 => to_signed(32705, LUT_AMPL_WIDTH),
		15745 => to_signed(32706, LUT_AMPL_WIDTH),
		15746 => to_signed(32706, LUT_AMPL_WIDTH),
		15747 => to_signed(32706, LUT_AMPL_WIDTH),
		15748 => to_signed(32706, LUT_AMPL_WIDTH),
		15749 => to_signed(32706, LUT_AMPL_WIDTH),
		15750 => to_signed(32706, LUT_AMPL_WIDTH),
		15751 => to_signed(32707, LUT_AMPL_WIDTH),
		15752 => to_signed(32707, LUT_AMPL_WIDTH),
		15753 => to_signed(32707, LUT_AMPL_WIDTH),
		15754 => to_signed(32707, LUT_AMPL_WIDTH),
		15755 => to_signed(32707, LUT_AMPL_WIDTH),
		15756 => to_signed(32708, LUT_AMPL_WIDTH),
		15757 => to_signed(32708, LUT_AMPL_WIDTH),
		15758 => to_signed(32708, LUT_AMPL_WIDTH),
		15759 => to_signed(32708, LUT_AMPL_WIDTH),
		15760 => to_signed(32708, LUT_AMPL_WIDTH),
		15761 => to_signed(32709, LUT_AMPL_WIDTH),
		15762 => to_signed(32709, LUT_AMPL_WIDTH),
		15763 => to_signed(32709, LUT_AMPL_WIDTH),
		15764 => to_signed(32709, LUT_AMPL_WIDTH),
		15765 => to_signed(32709, LUT_AMPL_WIDTH),
		15766 => to_signed(32710, LUT_AMPL_WIDTH),
		15767 => to_signed(32710, LUT_AMPL_WIDTH),
		15768 => to_signed(32710, LUT_AMPL_WIDTH),
		15769 => to_signed(32710, LUT_AMPL_WIDTH),
		15770 => to_signed(32710, LUT_AMPL_WIDTH),
		15771 => to_signed(32710, LUT_AMPL_WIDTH),
		15772 => to_signed(32711, LUT_AMPL_WIDTH),
		15773 => to_signed(32711, LUT_AMPL_WIDTH),
		15774 => to_signed(32711, LUT_AMPL_WIDTH),
		15775 => to_signed(32711, LUT_AMPL_WIDTH),
		15776 => to_signed(32711, LUT_AMPL_WIDTH),
		15777 => to_signed(32712, LUT_AMPL_WIDTH),
		15778 => to_signed(32712, LUT_AMPL_WIDTH),
		15779 => to_signed(32712, LUT_AMPL_WIDTH),
		15780 => to_signed(32712, LUT_AMPL_WIDTH),
		15781 => to_signed(32712, LUT_AMPL_WIDTH),
		15782 => to_signed(32712, LUT_AMPL_WIDTH),
		15783 => to_signed(32713, LUT_AMPL_WIDTH),
		15784 => to_signed(32713, LUT_AMPL_WIDTH),
		15785 => to_signed(32713, LUT_AMPL_WIDTH),
		15786 => to_signed(32713, LUT_AMPL_WIDTH),
		15787 => to_signed(32713, LUT_AMPL_WIDTH),
		15788 => to_signed(32714, LUT_AMPL_WIDTH),
		15789 => to_signed(32714, LUT_AMPL_WIDTH),
		15790 => to_signed(32714, LUT_AMPL_WIDTH),
		15791 => to_signed(32714, LUT_AMPL_WIDTH),
		15792 => to_signed(32714, LUT_AMPL_WIDTH),
		15793 => to_signed(32714, LUT_AMPL_WIDTH),
		15794 => to_signed(32715, LUT_AMPL_WIDTH),
		15795 => to_signed(32715, LUT_AMPL_WIDTH),
		15796 => to_signed(32715, LUT_AMPL_WIDTH),
		15797 => to_signed(32715, LUT_AMPL_WIDTH),
		15798 => to_signed(32715, LUT_AMPL_WIDTH),
		15799 => to_signed(32715, LUT_AMPL_WIDTH),
		15800 => to_signed(32716, LUT_AMPL_WIDTH),
		15801 => to_signed(32716, LUT_AMPL_WIDTH),
		15802 => to_signed(32716, LUT_AMPL_WIDTH),
		15803 => to_signed(32716, LUT_AMPL_WIDTH),
		15804 => to_signed(32716, LUT_AMPL_WIDTH),
		15805 => to_signed(32717, LUT_AMPL_WIDTH),
		15806 => to_signed(32717, LUT_AMPL_WIDTH),
		15807 => to_signed(32717, LUT_AMPL_WIDTH),
		15808 => to_signed(32717, LUT_AMPL_WIDTH),
		15809 => to_signed(32717, LUT_AMPL_WIDTH),
		15810 => to_signed(32717, LUT_AMPL_WIDTH),
		15811 => to_signed(32718, LUT_AMPL_WIDTH),
		15812 => to_signed(32718, LUT_AMPL_WIDTH),
		15813 => to_signed(32718, LUT_AMPL_WIDTH),
		15814 => to_signed(32718, LUT_AMPL_WIDTH),
		15815 => to_signed(32718, LUT_AMPL_WIDTH),
		15816 => to_signed(32718, LUT_AMPL_WIDTH),
		15817 => to_signed(32719, LUT_AMPL_WIDTH),
		15818 => to_signed(32719, LUT_AMPL_WIDTH),
		15819 => to_signed(32719, LUT_AMPL_WIDTH),
		15820 => to_signed(32719, LUT_AMPL_WIDTH),
		15821 => to_signed(32719, LUT_AMPL_WIDTH),
		15822 => to_signed(32719, LUT_AMPL_WIDTH),
		15823 => to_signed(32720, LUT_AMPL_WIDTH),
		15824 => to_signed(32720, LUT_AMPL_WIDTH),
		15825 => to_signed(32720, LUT_AMPL_WIDTH),
		15826 => to_signed(32720, LUT_AMPL_WIDTH),
		15827 => to_signed(32720, LUT_AMPL_WIDTH),
		15828 => to_signed(32720, LUT_AMPL_WIDTH),
		15829 => to_signed(32721, LUT_AMPL_WIDTH),
		15830 => to_signed(32721, LUT_AMPL_WIDTH),
		15831 => to_signed(32721, LUT_AMPL_WIDTH),
		15832 => to_signed(32721, LUT_AMPL_WIDTH),
		15833 => to_signed(32721, LUT_AMPL_WIDTH),
		15834 => to_signed(32721, LUT_AMPL_WIDTH),
		15835 => to_signed(32722, LUT_AMPL_WIDTH),
		15836 => to_signed(32722, LUT_AMPL_WIDTH),
		15837 => to_signed(32722, LUT_AMPL_WIDTH),
		15838 => to_signed(32722, LUT_AMPL_WIDTH),
		15839 => to_signed(32722, LUT_AMPL_WIDTH),
		15840 => to_signed(32722, LUT_AMPL_WIDTH),
		15841 => to_signed(32723, LUT_AMPL_WIDTH),
		15842 => to_signed(32723, LUT_AMPL_WIDTH),
		15843 => to_signed(32723, LUT_AMPL_WIDTH),
		15844 => to_signed(32723, LUT_AMPL_WIDTH),
		15845 => to_signed(32723, LUT_AMPL_WIDTH),
		15846 => to_signed(32723, LUT_AMPL_WIDTH),
		15847 => to_signed(32724, LUT_AMPL_WIDTH),
		15848 => to_signed(32724, LUT_AMPL_WIDTH),
		15849 => to_signed(32724, LUT_AMPL_WIDTH),
		15850 => to_signed(32724, LUT_AMPL_WIDTH),
		15851 => to_signed(32724, LUT_AMPL_WIDTH),
		15852 => to_signed(32724, LUT_AMPL_WIDTH),
		15853 => to_signed(32725, LUT_AMPL_WIDTH),
		15854 => to_signed(32725, LUT_AMPL_WIDTH),
		15855 => to_signed(32725, LUT_AMPL_WIDTH),
		15856 => to_signed(32725, LUT_AMPL_WIDTH),
		15857 => to_signed(32725, LUT_AMPL_WIDTH),
		15858 => to_signed(32725, LUT_AMPL_WIDTH),
		15859 => to_signed(32726, LUT_AMPL_WIDTH),
		15860 => to_signed(32726, LUT_AMPL_WIDTH),
		15861 => to_signed(32726, LUT_AMPL_WIDTH),
		15862 => to_signed(32726, LUT_AMPL_WIDTH),
		15863 => to_signed(32726, LUT_AMPL_WIDTH),
		15864 => to_signed(32726, LUT_AMPL_WIDTH),
		15865 => to_signed(32726, LUT_AMPL_WIDTH),
		15866 => to_signed(32727, LUT_AMPL_WIDTH),
		15867 => to_signed(32727, LUT_AMPL_WIDTH),
		15868 => to_signed(32727, LUT_AMPL_WIDTH),
		15869 => to_signed(32727, LUT_AMPL_WIDTH),
		15870 => to_signed(32727, LUT_AMPL_WIDTH),
		15871 => to_signed(32727, LUT_AMPL_WIDTH),
		15872 => to_signed(32728, LUT_AMPL_WIDTH),
		15873 => to_signed(32728, LUT_AMPL_WIDTH),
		15874 => to_signed(32728, LUT_AMPL_WIDTH),
		15875 => to_signed(32728, LUT_AMPL_WIDTH),
		15876 => to_signed(32728, LUT_AMPL_WIDTH),
		15877 => to_signed(32728, LUT_AMPL_WIDTH),
		15878 => to_signed(32728, LUT_AMPL_WIDTH),
		15879 => to_signed(32729, LUT_AMPL_WIDTH),
		15880 => to_signed(32729, LUT_AMPL_WIDTH),
		15881 => to_signed(32729, LUT_AMPL_WIDTH),
		15882 => to_signed(32729, LUT_AMPL_WIDTH),
		15883 => to_signed(32729, LUT_AMPL_WIDTH),
		15884 => to_signed(32729, LUT_AMPL_WIDTH),
		15885 => to_signed(32730, LUT_AMPL_WIDTH),
		15886 => to_signed(32730, LUT_AMPL_WIDTH),
		15887 => to_signed(32730, LUT_AMPL_WIDTH),
		15888 => to_signed(32730, LUT_AMPL_WIDTH),
		15889 => to_signed(32730, LUT_AMPL_WIDTH),
		15890 => to_signed(32730, LUT_AMPL_WIDTH),
		15891 => to_signed(32730, LUT_AMPL_WIDTH),
		15892 => to_signed(32731, LUT_AMPL_WIDTH),
		15893 => to_signed(32731, LUT_AMPL_WIDTH),
		15894 => to_signed(32731, LUT_AMPL_WIDTH),
		15895 => to_signed(32731, LUT_AMPL_WIDTH),
		15896 => to_signed(32731, LUT_AMPL_WIDTH),
		15897 => to_signed(32731, LUT_AMPL_WIDTH),
		15898 => to_signed(32731, LUT_AMPL_WIDTH),
		15899 => to_signed(32732, LUT_AMPL_WIDTH),
		15900 => to_signed(32732, LUT_AMPL_WIDTH),
		15901 => to_signed(32732, LUT_AMPL_WIDTH),
		15902 => to_signed(32732, LUT_AMPL_WIDTH),
		15903 => to_signed(32732, LUT_AMPL_WIDTH),
		15904 => to_signed(32732, LUT_AMPL_WIDTH),
		15905 => to_signed(32732, LUT_AMPL_WIDTH),
		15906 => to_signed(32733, LUT_AMPL_WIDTH),
		15907 => to_signed(32733, LUT_AMPL_WIDTH),
		15908 => to_signed(32733, LUT_AMPL_WIDTH),
		15909 => to_signed(32733, LUT_AMPL_WIDTH),
		15910 => to_signed(32733, LUT_AMPL_WIDTH),
		15911 => to_signed(32733, LUT_AMPL_WIDTH),
		15912 => to_signed(32733, LUT_AMPL_WIDTH),
		15913 => to_signed(32734, LUT_AMPL_WIDTH),
		15914 => to_signed(32734, LUT_AMPL_WIDTH),
		15915 => to_signed(32734, LUT_AMPL_WIDTH),
		15916 => to_signed(32734, LUT_AMPL_WIDTH),
		15917 => to_signed(32734, LUT_AMPL_WIDTH),
		15918 => to_signed(32734, LUT_AMPL_WIDTH),
		15919 => to_signed(32734, LUT_AMPL_WIDTH),
		15920 => to_signed(32735, LUT_AMPL_WIDTH),
		15921 => to_signed(32735, LUT_AMPL_WIDTH),
		15922 => to_signed(32735, LUT_AMPL_WIDTH),
		15923 => to_signed(32735, LUT_AMPL_WIDTH),
		15924 => to_signed(32735, LUT_AMPL_WIDTH),
		15925 => to_signed(32735, LUT_AMPL_WIDTH),
		15926 => to_signed(32735, LUT_AMPL_WIDTH),
		15927 => to_signed(32736, LUT_AMPL_WIDTH),
		15928 => to_signed(32736, LUT_AMPL_WIDTH),
		15929 => to_signed(32736, LUT_AMPL_WIDTH),
		15930 => to_signed(32736, LUT_AMPL_WIDTH),
		15931 => to_signed(32736, LUT_AMPL_WIDTH),
		15932 => to_signed(32736, LUT_AMPL_WIDTH),
		15933 => to_signed(32736, LUT_AMPL_WIDTH),
		15934 => to_signed(32737, LUT_AMPL_WIDTH),
		15935 => to_signed(32737, LUT_AMPL_WIDTH),
		15936 => to_signed(32737, LUT_AMPL_WIDTH),
		15937 => to_signed(32737, LUT_AMPL_WIDTH),
		15938 => to_signed(32737, LUT_AMPL_WIDTH),
		15939 => to_signed(32737, LUT_AMPL_WIDTH),
		15940 => to_signed(32737, LUT_AMPL_WIDTH),
		15941 => to_signed(32737, LUT_AMPL_WIDTH),
		15942 => to_signed(32738, LUT_AMPL_WIDTH),
		15943 => to_signed(32738, LUT_AMPL_WIDTH),
		15944 => to_signed(32738, LUT_AMPL_WIDTH),
		15945 => to_signed(32738, LUT_AMPL_WIDTH),
		15946 => to_signed(32738, LUT_AMPL_WIDTH),
		15947 => to_signed(32738, LUT_AMPL_WIDTH),
		15948 => to_signed(32738, LUT_AMPL_WIDTH),
		15949 => to_signed(32739, LUT_AMPL_WIDTH),
		15950 => to_signed(32739, LUT_AMPL_WIDTH),
		15951 => to_signed(32739, LUT_AMPL_WIDTH),
		15952 => to_signed(32739, LUT_AMPL_WIDTH),
		15953 => to_signed(32739, LUT_AMPL_WIDTH),
		15954 => to_signed(32739, LUT_AMPL_WIDTH),
		15955 => to_signed(32739, LUT_AMPL_WIDTH),
		15956 => to_signed(32739, LUT_AMPL_WIDTH),
		15957 => to_signed(32740, LUT_AMPL_WIDTH),
		15958 => to_signed(32740, LUT_AMPL_WIDTH),
		15959 => to_signed(32740, LUT_AMPL_WIDTH),
		15960 => to_signed(32740, LUT_AMPL_WIDTH),
		15961 => to_signed(32740, LUT_AMPL_WIDTH),
		15962 => to_signed(32740, LUT_AMPL_WIDTH),
		15963 => to_signed(32740, LUT_AMPL_WIDTH),
		15964 => to_signed(32740, LUT_AMPL_WIDTH),
		15965 => to_signed(32741, LUT_AMPL_WIDTH),
		15966 => to_signed(32741, LUT_AMPL_WIDTH),
		15967 => to_signed(32741, LUT_AMPL_WIDTH),
		15968 => to_signed(32741, LUT_AMPL_WIDTH),
		15969 => to_signed(32741, LUT_AMPL_WIDTH),
		15970 => to_signed(32741, LUT_AMPL_WIDTH),
		15971 => to_signed(32741, LUT_AMPL_WIDTH),
		15972 => to_signed(32741, LUT_AMPL_WIDTH),
		15973 => to_signed(32742, LUT_AMPL_WIDTH),
		15974 => to_signed(32742, LUT_AMPL_WIDTH),
		15975 => to_signed(32742, LUT_AMPL_WIDTH),
		15976 => to_signed(32742, LUT_AMPL_WIDTH),
		15977 => to_signed(32742, LUT_AMPL_WIDTH),
		15978 => to_signed(32742, LUT_AMPL_WIDTH),
		15979 => to_signed(32742, LUT_AMPL_WIDTH),
		15980 => to_signed(32742, LUT_AMPL_WIDTH),
		15981 => to_signed(32743, LUT_AMPL_WIDTH),
		15982 => to_signed(32743, LUT_AMPL_WIDTH),
		15983 => to_signed(32743, LUT_AMPL_WIDTH),
		15984 => to_signed(32743, LUT_AMPL_WIDTH),
		15985 => to_signed(32743, LUT_AMPL_WIDTH),
		15986 => to_signed(32743, LUT_AMPL_WIDTH),
		15987 => to_signed(32743, LUT_AMPL_WIDTH),
		15988 => to_signed(32743, LUT_AMPL_WIDTH),
		15989 => to_signed(32744, LUT_AMPL_WIDTH),
		15990 => to_signed(32744, LUT_AMPL_WIDTH),
		15991 => to_signed(32744, LUT_AMPL_WIDTH),
		15992 => to_signed(32744, LUT_AMPL_WIDTH),
		15993 => to_signed(32744, LUT_AMPL_WIDTH),
		15994 => to_signed(32744, LUT_AMPL_WIDTH),
		15995 => to_signed(32744, LUT_AMPL_WIDTH),
		15996 => to_signed(32744, LUT_AMPL_WIDTH),
		15997 => to_signed(32744, LUT_AMPL_WIDTH),
		15998 => to_signed(32745, LUT_AMPL_WIDTH),
		15999 => to_signed(32745, LUT_AMPL_WIDTH),
		16000 => to_signed(32745, LUT_AMPL_WIDTH),
		16001 => to_signed(32745, LUT_AMPL_WIDTH),
		16002 => to_signed(32745, LUT_AMPL_WIDTH),
		16003 => to_signed(32745, LUT_AMPL_WIDTH),
		16004 => to_signed(32745, LUT_AMPL_WIDTH),
		16005 => to_signed(32745, LUT_AMPL_WIDTH),
		16006 => to_signed(32745, LUT_AMPL_WIDTH),
		16007 => to_signed(32746, LUT_AMPL_WIDTH),
		16008 => to_signed(32746, LUT_AMPL_WIDTH),
		16009 => to_signed(32746, LUT_AMPL_WIDTH),
		16010 => to_signed(32746, LUT_AMPL_WIDTH),
		16011 => to_signed(32746, LUT_AMPL_WIDTH),
		16012 => to_signed(32746, LUT_AMPL_WIDTH),
		16013 => to_signed(32746, LUT_AMPL_WIDTH),
		16014 => to_signed(32746, LUT_AMPL_WIDTH),
		16015 => to_signed(32746, LUT_AMPL_WIDTH),
		16016 => to_signed(32747, LUT_AMPL_WIDTH),
		16017 => to_signed(32747, LUT_AMPL_WIDTH),
		16018 => to_signed(32747, LUT_AMPL_WIDTH),
		16019 => to_signed(32747, LUT_AMPL_WIDTH),
		16020 => to_signed(32747, LUT_AMPL_WIDTH),
		16021 => to_signed(32747, LUT_AMPL_WIDTH),
		16022 => to_signed(32747, LUT_AMPL_WIDTH),
		16023 => to_signed(32747, LUT_AMPL_WIDTH),
		16024 => to_signed(32747, LUT_AMPL_WIDTH),
		16025 => to_signed(32748, LUT_AMPL_WIDTH),
		16026 => to_signed(32748, LUT_AMPL_WIDTH),
		16027 => to_signed(32748, LUT_AMPL_WIDTH),
		16028 => to_signed(32748, LUT_AMPL_WIDTH),
		16029 => to_signed(32748, LUT_AMPL_WIDTH),
		16030 => to_signed(32748, LUT_AMPL_WIDTH),
		16031 => to_signed(32748, LUT_AMPL_WIDTH),
		16032 => to_signed(32748, LUT_AMPL_WIDTH),
		16033 => to_signed(32748, LUT_AMPL_WIDTH),
		16034 => to_signed(32749, LUT_AMPL_WIDTH),
		16035 => to_signed(32749, LUT_AMPL_WIDTH),
		16036 => to_signed(32749, LUT_AMPL_WIDTH),
		16037 => to_signed(32749, LUT_AMPL_WIDTH),
		16038 => to_signed(32749, LUT_AMPL_WIDTH),
		16039 => to_signed(32749, LUT_AMPL_WIDTH),
		16040 => to_signed(32749, LUT_AMPL_WIDTH),
		16041 => to_signed(32749, LUT_AMPL_WIDTH),
		16042 => to_signed(32749, LUT_AMPL_WIDTH),
		16043 => to_signed(32749, LUT_AMPL_WIDTH),
		16044 => to_signed(32750, LUT_AMPL_WIDTH),
		16045 => to_signed(32750, LUT_AMPL_WIDTH),
		16046 => to_signed(32750, LUT_AMPL_WIDTH),
		16047 => to_signed(32750, LUT_AMPL_WIDTH),
		16048 => to_signed(32750, LUT_AMPL_WIDTH),
		16049 => to_signed(32750, LUT_AMPL_WIDTH),
		16050 => to_signed(32750, LUT_AMPL_WIDTH),
		16051 => to_signed(32750, LUT_AMPL_WIDTH),
		16052 => to_signed(32750, LUT_AMPL_WIDTH),
		16053 => to_signed(32751, LUT_AMPL_WIDTH),
		16054 => to_signed(32751, LUT_AMPL_WIDTH),
		16055 => to_signed(32751, LUT_AMPL_WIDTH),
		16056 => to_signed(32751, LUT_AMPL_WIDTH),
		16057 => to_signed(32751, LUT_AMPL_WIDTH),
		16058 => to_signed(32751, LUT_AMPL_WIDTH),
		16059 => to_signed(32751, LUT_AMPL_WIDTH),
		16060 => to_signed(32751, LUT_AMPL_WIDTH),
		16061 => to_signed(32751, LUT_AMPL_WIDTH),
		16062 => to_signed(32751, LUT_AMPL_WIDTH),
		16063 => to_signed(32751, LUT_AMPL_WIDTH),
		16064 => to_signed(32752, LUT_AMPL_WIDTH),
		16065 => to_signed(32752, LUT_AMPL_WIDTH),
		16066 => to_signed(32752, LUT_AMPL_WIDTH),
		16067 => to_signed(32752, LUT_AMPL_WIDTH),
		16068 => to_signed(32752, LUT_AMPL_WIDTH),
		16069 => to_signed(32752, LUT_AMPL_WIDTH),
		16070 => to_signed(32752, LUT_AMPL_WIDTH),
		16071 => to_signed(32752, LUT_AMPL_WIDTH),
		16072 => to_signed(32752, LUT_AMPL_WIDTH),
		16073 => to_signed(32752, LUT_AMPL_WIDTH),
		16074 => to_signed(32753, LUT_AMPL_WIDTH),
		16075 => to_signed(32753, LUT_AMPL_WIDTH),
		16076 => to_signed(32753, LUT_AMPL_WIDTH),
		16077 => to_signed(32753, LUT_AMPL_WIDTH),
		16078 => to_signed(32753, LUT_AMPL_WIDTH),
		16079 => to_signed(32753, LUT_AMPL_WIDTH),
		16080 => to_signed(32753, LUT_AMPL_WIDTH),
		16081 => to_signed(32753, LUT_AMPL_WIDTH),
		16082 => to_signed(32753, LUT_AMPL_WIDTH),
		16083 => to_signed(32753, LUT_AMPL_WIDTH),
		16084 => to_signed(32753, LUT_AMPL_WIDTH),
		16085 => to_signed(32754, LUT_AMPL_WIDTH),
		16086 => to_signed(32754, LUT_AMPL_WIDTH),
		16087 => to_signed(32754, LUT_AMPL_WIDTH),
		16088 => to_signed(32754, LUT_AMPL_WIDTH),
		16089 => to_signed(32754, LUT_AMPL_WIDTH),
		16090 => to_signed(32754, LUT_AMPL_WIDTH),
		16091 => to_signed(32754, LUT_AMPL_WIDTH),
		16092 => to_signed(32754, LUT_AMPL_WIDTH),
		16093 => to_signed(32754, LUT_AMPL_WIDTH),
		16094 => to_signed(32754, LUT_AMPL_WIDTH),
		16095 => to_signed(32754, LUT_AMPL_WIDTH),
		16096 => to_signed(32755, LUT_AMPL_WIDTH),
		16097 => to_signed(32755, LUT_AMPL_WIDTH),
		16098 => to_signed(32755, LUT_AMPL_WIDTH),
		16099 => to_signed(32755, LUT_AMPL_WIDTH),
		16100 => to_signed(32755, LUT_AMPL_WIDTH),
		16101 => to_signed(32755, LUT_AMPL_WIDTH),
		16102 => to_signed(32755, LUT_AMPL_WIDTH),
		16103 => to_signed(32755, LUT_AMPL_WIDTH),
		16104 => to_signed(32755, LUT_AMPL_WIDTH),
		16105 => to_signed(32755, LUT_AMPL_WIDTH),
		16106 => to_signed(32755, LUT_AMPL_WIDTH),
		16107 => to_signed(32755, LUT_AMPL_WIDTH),
		16108 => to_signed(32756, LUT_AMPL_WIDTH),
		16109 => to_signed(32756, LUT_AMPL_WIDTH),
		16110 => to_signed(32756, LUT_AMPL_WIDTH),
		16111 => to_signed(32756, LUT_AMPL_WIDTH),
		16112 => to_signed(32756, LUT_AMPL_WIDTH),
		16113 => to_signed(32756, LUT_AMPL_WIDTH),
		16114 => to_signed(32756, LUT_AMPL_WIDTH),
		16115 => to_signed(32756, LUT_AMPL_WIDTH),
		16116 => to_signed(32756, LUT_AMPL_WIDTH),
		16117 => to_signed(32756, LUT_AMPL_WIDTH),
		16118 => to_signed(32756, LUT_AMPL_WIDTH),
		16119 => to_signed(32756, LUT_AMPL_WIDTH),
		16120 => to_signed(32757, LUT_AMPL_WIDTH),
		16121 => to_signed(32757, LUT_AMPL_WIDTH),
		16122 => to_signed(32757, LUT_AMPL_WIDTH),
		16123 => to_signed(32757, LUT_AMPL_WIDTH),
		16124 => to_signed(32757, LUT_AMPL_WIDTH),
		16125 => to_signed(32757, LUT_AMPL_WIDTH),
		16126 => to_signed(32757, LUT_AMPL_WIDTH),
		16127 => to_signed(32757, LUT_AMPL_WIDTH),
		16128 => to_signed(32757, LUT_AMPL_WIDTH),
		16129 => to_signed(32757, LUT_AMPL_WIDTH),
		16130 => to_signed(32757, LUT_AMPL_WIDTH),
		16131 => to_signed(32757, LUT_AMPL_WIDTH),
		16132 => to_signed(32757, LUT_AMPL_WIDTH),
		16133 => to_signed(32758, LUT_AMPL_WIDTH),
		16134 => to_signed(32758, LUT_AMPL_WIDTH),
		16135 => to_signed(32758, LUT_AMPL_WIDTH),
		16136 => to_signed(32758, LUT_AMPL_WIDTH),
		16137 => to_signed(32758, LUT_AMPL_WIDTH),
		16138 => to_signed(32758, LUT_AMPL_WIDTH),
		16139 => to_signed(32758, LUT_AMPL_WIDTH),
		16140 => to_signed(32758, LUT_AMPL_WIDTH),
		16141 => to_signed(32758, LUT_AMPL_WIDTH),
		16142 => to_signed(32758, LUT_AMPL_WIDTH),
		16143 => to_signed(32758, LUT_AMPL_WIDTH),
		16144 => to_signed(32758, LUT_AMPL_WIDTH),
		16145 => to_signed(32758, LUT_AMPL_WIDTH),
		16146 => to_signed(32758, LUT_AMPL_WIDTH),
		16147 => to_signed(32759, LUT_AMPL_WIDTH),
		16148 => to_signed(32759, LUT_AMPL_WIDTH),
		16149 => to_signed(32759, LUT_AMPL_WIDTH),
		16150 => to_signed(32759, LUT_AMPL_WIDTH),
		16151 => to_signed(32759, LUT_AMPL_WIDTH),
		16152 => to_signed(32759, LUT_AMPL_WIDTH),
		16153 => to_signed(32759, LUT_AMPL_WIDTH),
		16154 => to_signed(32759, LUT_AMPL_WIDTH),
		16155 => to_signed(32759, LUT_AMPL_WIDTH),
		16156 => to_signed(32759, LUT_AMPL_WIDTH),
		16157 => to_signed(32759, LUT_AMPL_WIDTH),
		16158 => to_signed(32759, LUT_AMPL_WIDTH),
		16159 => to_signed(32759, LUT_AMPL_WIDTH),
		16160 => to_signed(32759, LUT_AMPL_WIDTH),
		16161 => to_signed(32760, LUT_AMPL_WIDTH),
		16162 => to_signed(32760, LUT_AMPL_WIDTH),
		16163 => to_signed(32760, LUT_AMPL_WIDTH),
		16164 => to_signed(32760, LUT_AMPL_WIDTH),
		16165 => to_signed(32760, LUT_AMPL_WIDTH),
		16166 => to_signed(32760, LUT_AMPL_WIDTH),
		16167 => to_signed(32760, LUT_AMPL_WIDTH),
		16168 => to_signed(32760, LUT_AMPL_WIDTH),
		16169 => to_signed(32760, LUT_AMPL_WIDTH),
		16170 => to_signed(32760, LUT_AMPL_WIDTH),
		16171 => to_signed(32760, LUT_AMPL_WIDTH),
		16172 => to_signed(32760, LUT_AMPL_WIDTH),
		16173 => to_signed(32760, LUT_AMPL_WIDTH),
		16174 => to_signed(32760, LUT_AMPL_WIDTH),
		16175 => to_signed(32760, LUT_AMPL_WIDTH),
		16176 => to_signed(32760, LUT_AMPL_WIDTH),
		16177 => to_signed(32761, LUT_AMPL_WIDTH),
		16178 => to_signed(32761, LUT_AMPL_WIDTH),
		16179 => to_signed(32761, LUT_AMPL_WIDTH),
		16180 => to_signed(32761, LUT_AMPL_WIDTH),
		16181 => to_signed(32761, LUT_AMPL_WIDTH),
		16182 => to_signed(32761, LUT_AMPL_WIDTH),
		16183 => to_signed(32761, LUT_AMPL_WIDTH),
		16184 => to_signed(32761, LUT_AMPL_WIDTH),
		16185 => to_signed(32761, LUT_AMPL_WIDTH),
		16186 => to_signed(32761, LUT_AMPL_WIDTH),
		16187 => to_signed(32761, LUT_AMPL_WIDTH),
		16188 => to_signed(32761, LUT_AMPL_WIDTH),
		16189 => to_signed(32761, LUT_AMPL_WIDTH),
		16190 => to_signed(32761, LUT_AMPL_WIDTH),
		16191 => to_signed(32761, LUT_AMPL_WIDTH),
		16192 => to_signed(32761, LUT_AMPL_WIDTH),
		16193 => to_signed(32762, LUT_AMPL_WIDTH),
		16194 => to_signed(32762, LUT_AMPL_WIDTH),
		16195 => to_signed(32762, LUT_AMPL_WIDTH),
		16196 => to_signed(32762, LUT_AMPL_WIDTH),
		16197 => to_signed(32762, LUT_AMPL_WIDTH),
		16198 => to_signed(32762, LUT_AMPL_WIDTH),
		16199 => to_signed(32762, LUT_AMPL_WIDTH),
		16200 => to_signed(32762, LUT_AMPL_WIDTH),
		16201 => to_signed(32762, LUT_AMPL_WIDTH),
		16202 => to_signed(32762, LUT_AMPL_WIDTH),
		16203 => to_signed(32762, LUT_AMPL_WIDTH),
		16204 => to_signed(32762, LUT_AMPL_WIDTH),
		16205 => to_signed(32762, LUT_AMPL_WIDTH),
		16206 => to_signed(32762, LUT_AMPL_WIDTH),
		16207 => to_signed(32762, LUT_AMPL_WIDTH),
		16208 => to_signed(32762, LUT_AMPL_WIDTH),
		16209 => to_signed(32762, LUT_AMPL_WIDTH),
		16210 => to_signed(32762, LUT_AMPL_WIDTH),
		16211 => to_signed(32762, LUT_AMPL_WIDTH),
		16212 => to_signed(32763, LUT_AMPL_WIDTH),
		16213 => to_signed(32763, LUT_AMPL_WIDTH),
		16214 => to_signed(32763, LUT_AMPL_WIDTH),
		16215 => to_signed(32763, LUT_AMPL_WIDTH),
		16216 => to_signed(32763, LUT_AMPL_WIDTH),
		16217 => to_signed(32763, LUT_AMPL_WIDTH),
		16218 => to_signed(32763, LUT_AMPL_WIDTH),
		16219 => to_signed(32763, LUT_AMPL_WIDTH),
		16220 => to_signed(32763, LUT_AMPL_WIDTH),
		16221 => to_signed(32763, LUT_AMPL_WIDTH),
		16222 => to_signed(32763, LUT_AMPL_WIDTH),
		16223 => to_signed(32763, LUT_AMPL_WIDTH),
		16224 => to_signed(32763, LUT_AMPL_WIDTH),
		16225 => to_signed(32763, LUT_AMPL_WIDTH),
		16226 => to_signed(32763, LUT_AMPL_WIDTH),
		16227 => to_signed(32763, LUT_AMPL_WIDTH),
		16228 => to_signed(32763, LUT_AMPL_WIDTH),
		16229 => to_signed(32763, LUT_AMPL_WIDTH),
		16230 => to_signed(32763, LUT_AMPL_WIDTH),
		16231 => to_signed(32763, LUT_AMPL_WIDTH),
		16232 => to_signed(32764, LUT_AMPL_WIDTH),
		16233 => to_signed(32764, LUT_AMPL_WIDTH),
		16234 => to_signed(32764, LUT_AMPL_WIDTH),
		16235 => to_signed(32764, LUT_AMPL_WIDTH),
		16236 => to_signed(32764, LUT_AMPL_WIDTH),
		16237 => to_signed(32764, LUT_AMPL_WIDTH),
		16238 => to_signed(32764, LUT_AMPL_WIDTH),
		16239 => to_signed(32764, LUT_AMPL_WIDTH),
		16240 => to_signed(32764, LUT_AMPL_WIDTH),
		16241 => to_signed(32764, LUT_AMPL_WIDTH),
		16242 => to_signed(32764, LUT_AMPL_WIDTH),
		16243 => to_signed(32764, LUT_AMPL_WIDTH),
		16244 => to_signed(32764, LUT_AMPL_WIDTH),
		16245 => to_signed(32764, LUT_AMPL_WIDTH),
		16246 => to_signed(32764, LUT_AMPL_WIDTH),
		16247 => to_signed(32764, LUT_AMPL_WIDTH),
		16248 => to_signed(32764, LUT_AMPL_WIDTH),
		16249 => to_signed(32764, LUT_AMPL_WIDTH),
		16250 => to_signed(32764, LUT_AMPL_WIDTH),
		16251 => to_signed(32764, LUT_AMPL_WIDTH),
		16252 => to_signed(32764, LUT_AMPL_WIDTH),
		16253 => to_signed(32764, LUT_AMPL_WIDTH),
		16254 => to_signed(32764, LUT_AMPL_WIDTH),
		16255 => to_signed(32764, LUT_AMPL_WIDTH),
		16256 => to_signed(32765, LUT_AMPL_WIDTH),
		16257 => to_signed(32765, LUT_AMPL_WIDTH),
		16258 => to_signed(32765, LUT_AMPL_WIDTH),
		16259 => to_signed(32765, LUT_AMPL_WIDTH),
		16260 => to_signed(32765, LUT_AMPL_WIDTH),
		16261 => to_signed(32765, LUT_AMPL_WIDTH),
		16262 => to_signed(32765, LUT_AMPL_WIDTH),
		16263 => to_signed(32765, LUT_AMPL_WIDTH),
		16264 => to_signed(32765, LUT_AMPL_WIDTH),
		16265 => to_signed(32765, LUT_AMPL_WIDTH),
		16266 => to_signed(32765, LUT_AMPL_WIDTH),
		16267 => to_signed(32765, LUT_AMPL_WIDTH),
		16268 => to_signed(32765, LUT_AMPL_WIDTH),
		16269 => to_signed(32765, LUT_AMPL_WIDTH),
		16270 => to_signed(32765, LUT_AMPL_WIDTH),
		16271 => to_signed(32765, LUT_AMPL_WIDTH),
		16272 => to_signed(32765, LUT_AMPL_WIDTH),
		16273 => to_signed(32765, LUT_AMPL_WIDTH),
		16274 => to_signed(32765, LUT_AMPL_WIDTH),
		16275 => to_signed(32765, LUT_AMPL_WIDTH),
		16276 => to_signed(32765, LUT_AMPL_WIDTH),
		16277 => to_signed(32765, LUT_AMPL_WIDTH),
		16278 => to_signed(32765, LUT_AMPL_WIDTH),
		16279 => to_signed(32765, LUT_AMPL_WIDTH),
		16280 => to_signed(32765, LUT_AMPL_WIDTH),
		16281 => to_signed(32765, LUT_AMPL_WIDTH),
		16282 => to_signed(32765, LUT_AMPL_WIDTH),
		16283 => to_signed(32765, LUT_AMPL_WIDTH),
		16284 => to_signed(32765, LUT_AMPL_WIDTH),
		16285 => to_signed(32766, LUT_AMPL_WIDTH),
		16286 => to_signed(32766, LUT_AMPL_WIDTH),
		16287 => to_signed(32766, LUT_AMPL_WIDTH),
		16288 => to_signed(32766, LUT_AMPL_WIDTH),
		16289 => to_signed(32766, LUT_AMPL_WIDTH),
		16290 => to_signed(32766, LUT_AMPL_WIDTH),
		16291 => to_signed(32766, LUT_AMPL_WIDTH),
		16292 => to_signed(32766, LUT_AMPL_WIDTH),
		16293 => to_signed(32766, LUT_AMPL_WIDTH),
		16294 => to_signed(32766, LUT_AMPL_WIDTH),
		16295 => to_signed(32766, LUT_AMPL_WIDTH),
		16296 => to_signed(32766, LUT_AMPL_WIDTH),
		16297 => to_signed(32766, LUT_AMPL_WIDTH),
		16298 => to_signed(32766, LUT_AMPL_WIDTH),
		16299 => to_signed(32766, LUT_AMPL_WIDTH),
		16300 => to_signed(32766, LUT_AMPL_WIDTH),
		16301 => to_signed(32766, LUT_AMPL_WIDTH),
		16302 => to_signed(32766, LUT_AMPL_WIDTH),
		16303 => to_signed(32766, LUT_AMPL_WIDTH),
		16304 => to_signed(32766, LUT_AMPL_WIDTH),
		16305 => to_signed(32766, LUT_AMPL_WIDTH),
		16306 => to_signed(32766, LUT_AMPL_WIDTH),
		16307 => to_signed(32766, LUT_AMPL_WIDTH),
		16308 => to_signed(32766, LUT_AMPL_WIDTH),
		16309 => to_signed(32766, LUT_AMPL_WIDTH),
		16310 => to_signed(32766, LUT_AMPL_WIDTH),
		16311 => to_signed(32766, LUT_AMPL_WIDTH),
		16312 => to_signed(32766, LUT_AMPL_WIDTH),
		16313 => to_signed(32766, LUT_AMPL_WIDTH),
		16314 => to_signed(32766, LUT_AMPL_WIDTH),
		16315 => to_signed(32766, LUT_AMPL_WIDTH),
		16316 => to_signed(32766, LUT_AMPL_WIDTH),
		16317 => to_signed(32766, LUT_AMPL_WIDTH),
		16318 => to_signed(32766, LUT_AMPL_WIDTH),
		16319 => to_signed(32766, LUT_AMPL_WIDTH),
		16320 => to_signed(32766, LUT_AMPL_WIDTH),
		16321 => to_signed(32766, LUT_AMPL_WIDTH),
		16322 => to_signed(32766, LUT_AMPL_WIDTH),
		16323 => to_signed(32766, LUT_AMPL_WIDTH),
		16324 => to_signed(32766, LUT_AMPL_WIDTH),
		16325 => to_signed(32766, LUT_AMPL_WIDTH),
		16326 => to_signed(32766, LUT_AMPL_WIDTH),
		16327 => to_signed(32767, LUT_AMPL_WIDTH),
		16328 => to_signed(32767, LUT_AMPL_WIDTH),
		16329 => to_signed(32767, LUT_AMPL_WIDTH),
		16330 => to_signed(32767, LUT_AMPL_WIDTH),
		16331 => to_signed(32767, LUT_AMPL_WIDTH),
		16332 => to_signed(32767, LUT_AMPL_WIDTH),
		16333 => to_signed(32767, LUT_AMPL_WIDTH),
		16334 => to_signed(32767, LUT_AMPL_WIDTH),
		16335 => to_signed(32767, LUT_AMPL_WIDTH),
		16336 => to_signed(32767, LUT_AMPL_WIDTH),
		16337 => to_signed(32767, LUT_AMPL_WIDTH),
		16338 => to_signed(32767, LUT_AMPL_WIDTH),
		16339 => to_signed(32767, LUT_AMPL_WIDTH),
		16340 => to_signed(32767, LUT_AMPL_WIDTH),
		16341 => to_signed(32767, LUT_AMPL_WIDTH),
		16342 => to_signed(32767, LUT_AMPL_WIDTH),
		16343 => to_signed(32767, LUT_AMPL_WIDTH),
		16344 => to_signed(32767, LUT_AMPL_WIDTH),
		16345 => to_signed(32767, LUT_AMPL_WIDTH),
		16346 => to_signed(32767, LUT_AMPL_WIDTH),
		16347 => to_signed(32767, LUT_AMPL_WIDTH),
		16348 => to_signed(32767, LUT_AMPL_WIDTH),
		16349 => to_signed(32767, LUT_AMPL_WIDTH),
		16350 => to_signed(32767, LUT_AMPL_WIDTH),
		16351 => to_signed(32767, LUT_AMPL_WIDTH),
		16352 => to_signed(32767, LUT_AMPL_WIDTH),
		16353 => to_signed(32767, LUT_AMPL_WIDTH),
		16354 => to_signed(32767, LUT_AMPL_WIDTH),
		16355 => to_signed(32767, LUT_AMPL_WIDTH),
		16356 => to_signed(32767, LUT_AMPL_WIDTH),
		16357 => to_signed(32767, LUT_AMPL_WIDTH),
		16358 => to_signed(32767, LUT_AMPL_WIDTH),
		16359 => to_signed(32767, LUT_AMPL_WIDTH),
		16360 => to_signed(32767, LUT_AMPL_WIDTH),
		16361 => to_signed(32767, LUT_AMPL_WIDTH),
		16362 => to_signed(32767, LUT_AMPL_WIDTH),
		16363 => to_signed(32767, LUT_AMPL_WIDTH),
		16364 => to_signed(32767, LUT_AMPL_WIDTH),
		16365 => to_signed(32767, LUT_AMPL_WIDTH),
		16366 => to_signed(32767, LUT_AMPL_WIDTH),
		16367 => to_signed(32767, LUT_AMPL_WIDTH),
		16368 => to_signed(32767, LUT_AMPL_WIDTH),
		16369 => to_signed(32767, LUT_AMPL_WIDTH),
		16370 => to_signed(32767, LUT_AMPL_WIDTH),
		16371 => to_signed(32767, LUT_AMPL_WIDTH),
		16372 => to_signed(32767, LUT_AMPL_WIDTH),
		16373 => to_signed(32767, LUT_AMPL_WIDTH),
		16374 => to_signed(32767, LUT_AMPL_WIDTH),
		16375 => to_signed(32767, LUT_AMPL_WIDTH),
		16376 => to_signed(32767, LUT_AMPL_WIDTH),
		16377 => to_signed(32767, LUT_AMPL_WIDTH),
		16378 => to_signed(32767, LUT_AMPL_WIDTH),
		16379 => to_signed(32767, LUT_AMPL_WIDTH),
		16380 => to_signed(32767, LUT_AMPL_WIDTH),
		16381 => to_signed(32767, LUT_AMPL_WIDTH),
		16382 => to_signed(32767, LUT_AMPL_WIDTH),
		16383 => to_signed(32767, LUT_AMPL_WIDTH),
		16384 => to_signed(32767, LUT_AMPL_WIDTH),
		16385 => to_signed(32767, LUT_AMPL_WIDTH),
		16386 => to_signed(32767, LUT_AMPL_WIDTH),
		16387 => to_signed(32767, LUT_AMPL_WIDTH),
		16388 => to_signed(32767, LUT_AMPL_WIDTH),
		16389 => to_signed(32767, LUT_AMPL_WIDTH),
		16390 => to_signed(32767, LUT_AMPL_WIDTH),
		16391 => to_signed(32767, LUT_AMPL_WIDTH),
		16392 => to_signed(32767, LUT_AMPL_WIDTH),
		16393 => to_signed(32767, LUT_AMPL_WIDTH),
		16394 => to_signed(32767, LUT_AMPL_WIDTH),
		16395 => to_signed(32767, LUT_AMPL_WIDTH),
		16396 => to_signed(32767, LUT_AMPL_WIDTH),
		16397 => to_signed(32767, LUT_AMPL_WIDTH),
		16398 => to_signed(32767, LUT_AMPL_WIDTH),
		16399 => to_signed(32767, LUT_AMPL_WIDTH),
		16400 => to_signed(32767, LUT_AMPL_WIDTH),
		16401 => to_signed(32767, LUT_AMPL_WIDTH),
		16402 => to_signed(32767, LUT_AMPL_WIDTH),
		16403 => to_signed(32767, LUT_AMPL_WIDTH),
		16404 => to_signed(32767, LUT_AMPL_WIDTH),
		16405 => to_signed(32767, LUT_AMPL_WIDTH),
		16406 => to_signed(32767, LUT_AMPL_WIDTH),
		16407 => to_signed(32767, LUT_AMPL_WIDTH),
		16408 => to_signed(32767, LUT_AMPL_WIDTH),
		16409 => to_signed(32767, LUT_AMPL_WIDTH),
		16410 => to_signed(32767, LUT_AMPL_WIDTH),
		16411 => to_signed(32767, LUT_AMPL_WIDTH),
		16412 => to_signed(32767, LUT_AMPL_WIDTH),
		16413 => to_signed(32767, LUT_AMPL_WIDTH),
		16414 => to_signed(32767, LUT_AMPL_WIDTH),
		16415 => to_signed(32767, LUT_AMPL_WIDTH),
		16416 => to_signed(32767, LUT_AMPL_WIDTH),
		16417 => to_signed(32767, LUT_AMPL_WIDTH),
		16418 => to_signed(32767, LUT_AMPL_WIDTH),
		16419 => to_signed(32767, LUT_AMPL_WIDTH),
		16420 => to_signed(32767, LUT_AMPL_WIDTH),
		16421 => to_signed(32767, LUT_AMPL_WIDTH),
		16422 => to_signed(32767, LUT_AMPL_WIDTH),
		16423 => to_signed(32767, LUT_AMPL_WIDTH),
		16424 => to_signed(32767, LUT_AMPL_WIDTH),
		16425 => to_signed(32767, LUT_AMPL_WIDTH),
		16426 => to_signed(32767, LUT_AMPL_WIDTH),
		16427 => to_signed(32767, LUT_AMPL_WIDTH),
		16428 => to_signed(32767, LUT_AMPL_WIDTH),
		16429 => to_signed(32767, LUT_AMPL_WIDTH),
		16430 => to_signed(32767, LUT_AMPL_WIDTH),
		16431 => to_signed(32767, LUT_AMPL_WIDTH),
		16432 => to_signed(32767, LUT_AMPL_WIDTH),
		16433 => to_signed(32767, LUT_AMPL_WIDTH),
		16434 => to_signed(32767, LUT_AMPL_WIDTH),
		16435 => to_signed(32767, LUT_AMPL_WIDTH),
		16436 => to_signed(32767, LUT_AMPL_WIDTH),
		16437 => to_signed(32767, LUT_AMPL_WIDTH),
		16438 => to_signed(32767, LUT_AMPL_WIDTH),
		16439 => to_signed(32767, LUT_AMPL_WIDTH),
		16440 => to_signed(32767, LUT_AMPL_WIDTH),
		16441 => to_signed(32767, LUT_AMPL_WIDTH),
		16442 => to_signed(32766, LUT_AMPL_WIDTH),
		16443 => to_signed(32766, LUT_AMPL_WIDTH),
		16444 => to_signed(32766, LUT_AMPL_WIDTH),
		16445 => to_signed(32766, LUT_AMPL_WIDTH),
		16446 => to_signed(32766, LUT_AMPL_WIDTH),
		16447 => to_signed(32766, LUT_AMPL_WIDTH),
		16448 => to_signed(32766, LUT_AMPL_WIDTH),
		16449 => to_signed(32766, LUT_AMPL_WIDTH),
		16450 => to_signed(32766, LUT_AMPL_WIDTH),
		16451 => to_signed(32766, LUT_AMPL_WIDTH),
		16452 => to_signed(32766, LUT_AMPL_WIDTH),
		16453 => to_signed(32766, LUT_AMPL_WIDTH),
		16454 => to_signed(32766, LUT_AMPL_WIDTH),
		16455 => to_signed(32766, LUT_AMPL_WIDTH),
		16456 => to_signed(32766, LUT_AMPL_WIDTH),
		16457 => to_signed(32766, LUT_AMPL_WIDTH),
		16458 => to_signed(32766, LUT_AMPL_WIDTH),
		16459 => to_signed(32766, LUT_AMPL_WIDTH),
		16460 => to_signed(32766, LUT_AMPL_WIDTH),
		16461 => to_signed(32766, LUT_AMPL_WIDTH),
		16462 => to_signed(32766, LUT_AMPL_WIDTH),
		16463 => to_signed(32766, LUT_AMPL_WIDTH),
		16464 => to_signed(32766, LUT_AMPL_WIDTH),
		16465 => to_signed(32766, LUT_AMPL_WIDTH),
		16466 => to_signed(32766, LUT_AMPL_WIDTH),
		16467 => to_signed(32766, LUT_AMPL_WIDTH),
		16468 => to_signed(32766, LUT_AMPL_WIDTH),
		16469 => to_signed(32766, LUT_AMPL_WIDTH),
		16470 => to_signed(32766, LUT_AMPL_WIDTH),
		16471 => to_signed(32766, LUT_AMPL_WIDTH),
		16472 => to_signed(32766, LUT_AMPL_WIDTH),
		16473 => to_signed(32766, LUT_AMPL_WIDTH),
		16474 => to_signed(32766, LUT_AMPL_WIDTH),
		16475 => to_signed(32766, LUT_AMPL_WIDTH),
		16476 => to_signed(32766, LUT_AMPL_WIDTH),
		16477 => to_signed(32766, LUT_AMPL_WIDTH),
		16478 => to_signed(32766, LUT_AMPL_WIDTH),
		16479 => to_signed(32766, LUT_AMPL_WIDTH),
		16480 => to_signed(32766, LUT_AMPL_WIDTH),
		16481 => to_signed(32766, LUT_AMPL_WIDTH),
		16482 => to_signed(32766, LUT_AMPL_WIDTH),
		16483 => to_signed(32766, LUT_AMPL_WIDTH),
		16484 => to_signed(32765, LUT_AMPL_WIDTH),
		16485 => to_signed(32765, LUT_AMPL_WIDTH),
		16486 => to_signed(32765, LUT_AMPL_WIDTH),
		16487 => to_signed(32765, LUT_AMPL_WIDTH),
		16488 => to_signed(32765, LUT_AMPL_WIDTH),
		16489 => to_signed(32765, LUT_AMPL_WIDTH),
		16490 => to_signed(32765, LUT_AMPL_WIDTH),
		16491 => to_signed(32765, LUT_AMPL_WIDTH),
		16492 => to_signed(32765, LUT_AMPL_WIDTH),
		16493 => to_signed(32765, LUT_AMPL_WIDTH),
		16494 => to_signed(32765, LUT_AMPL_WIDTH),
		16495 => to_signed(32765, LUT_AMPL_WIDTH),
		16496 => to_signed(32765, LUT_AMPL_WIDTH),
		16497 => to_signed(32765, LUT_AMPL_WIDTH),
		16498 => to_signed(32765, LUT_AMPL_WIDTH),
		16499 => to_signed(32765, LUT_AMPL_WIDTH),
		16500 => to_signed(32765, LUT_AMPL_WIDTH),
		16501 => to_signed(32765, LUT_AMPL_WIDTH),
		16502 => to_signed(32765, LUT_AMPL_WIDTH),
		16503 => to_signed(32765, LUT_AMPL_WIDTH),
		16504 => to_signed(32765, LUT_AMPL_WIDTH),
		16505 => to_signed(32765, LUT_AMPL_WIDTH),
		16506 => to_signed(32765, LUT_AMPL_WIDTH),
		16507 => to_signed(32765, LUT_AMPL_WIDTH),
		16508 => to_signed(32765, LUT_AMPL_WIDTH),
		16509 => to_signed(32765, LUT_AMPL_WIDTH),
		16510 => to_signed(32765, LUT_AMPL_WIDTH),
		16511 => to_signed(32765, LUT_AMPL_WIDTH),
		16512 => to_signed(32765, LUT_AMPL_WIDTH),
		16513 => to_signed(32764, LUT_AMPL_WIDTH),
		16514 => to_signed(32764, LUT_AMPL_WIDTH),
		16515 => to_signed(32764, LUT_AMPL_WIDTH),
		16516 => to_signed(32764, LUT_AMPL_WIDTH),
		16517 => to_signed(32764, LUT_AMPL_WIDTH),
		16518 => to_signed(32764, LUT_AMPL_WIDTH),
		16519 => to_signed(32764, LUT_AMPL_WIDTH),
		16520 => to_signed(32764, LUT_AMPL_WIDTH),
		16521 => to_signed(32764, LUT_AMPL_WIDTH),
		16522 => to_signed(32764, LUT_AMPL_WIDTH),
		16523 => to_signed(32764, LUT_AMPL_WIDTH),
		16524 => to_signed(32764, LUT_AMPL_WIDTH),
		16525 => to_signed(32764, LUT_AMPL_WIDTH),
		16526 => to_signed(32764, LUT_AMPL_WIDTH),
		16527 => to_signed(32764, LUT_AMPL_WIDTH),
		16528 => to_signed(32764, LUT_AMPL_WIDTH),
		16529 => to_signed(32764, LUT_AMPL_WIDTH),
		16530 => to_signed(32764, LUT_AMPL_WIDTH),
		16531 => to_signed(32764, LUT_AMPL_WIDTH),
		16532 => to_signed(32764, LUT_AMPL_WIDTH),
		16533 => to_signed(32764, LUT_AMPL_WIDTH),
		16534 => to_signed(32764, LUT_AMPL_WIDTH),
		16535 => to_signed(32764, LUT_AMPL_WIDTH),
		16536 => to_signed(32764, LUT_AMPL_WIDTH),
		16537 => to_signed(32763, LUT_AMPL_WIDTH),
		16538 => to_signed(32763, LUT_AMPL_WIDTH),
		16539 => to_signed(32763, LUT_AMPL_WIDTH),
		16540 => to_signed(32763, LUT_AMPL_WIDTH),
		16541 => to_signed(32763, LUT_AMPL_WIDTH),
		16542 => to_signed(32763, LUT_AMPL_WIDTH),
		16543 => to_signed(32763, LUT_AMPL_WIDTH),
		16544 => to_signed(32763, LUT_AMPL_WIDTH),
		16545 => to_signed(32763, LUT_AMPL_WIDTH),
		16546 => to_signed(32763, LUT_AMPL_WIDTH),
		16547 => to_signed(32763, LUT_AMPL_WIDTH),
		16548 => to_signed(32763, LUT_AMPL_WIDTH),
		16549 => to_signed(32763, LUT_AMPL_WIDTH),
		16550 => to_signed(32763, LUT_AMPL_WIDTH),
		16551 => to_signed(32763, LUT_AMPL_WIDTH),
		16552 => to_signed(32763, LUT_AMPL_WIDTH),
		16553 => to_signed(32763, LUT_AMPL_WIDTH),
		16554 => to_signed(32763, LUT_AMPL_WIDTH),
		16555 => to_signed(32763, LUT_AMPL_WIDTH),
		16556 => to_signed(32763, LUT_AMPL_WIDTH),
		16557 => to_signed(32762, LUT_AMPL_WIDTH),
		16558 => to_signed(32762, LUT_AMPL_WIDTH),
		16559 => to_signed(32762, LUT_AMPL_WIDTH),
		16560 => to_signed(32762, LUT_AMPL_WIDTH),
		16561 => to_signed(32762, LUT_AMPL_WIDTH),
		16562 => to_signed(32762, LUT_AMPL_WIDTH),
		16563 => to_signed(32762, LUT_AMPL_WIDTH),
		16564 => to_signed(32762, LUT_AMPL_WIDTH),
		16565 => to_signed(32762, LUT_AMPL_WIDTH),
		16566 => to_signed(32762, LUT_AMPL_WIDTH),
		16567 => to_signed(32762, LUT_AMPL_WIDTH),
		16568 => to_signed(32762, LUT_AMPL_WIDTH),
		16569 => to_signed(32762, LUT_AMPL_WIDTH),
		16570 => to_signed(32762, LUT_AMPL_WIDTH),
		16571 => to_signed(32762, LUT_AMPL_WIDTH),
		16572 => to_signed(32762, LUT_AMPL_WIDTH),
		16573 => to_signed(32762, LUT_AMPL_WIDTH),
		16574 => to_signed(32762, LUT_AMPL_WIDTH),
		16575 => to_signed(32762, LUT_AMPL_WIDTH),
		16576 => to_signed(32761, LUT_AMPL_WIDTH),
		16577 => to_signed(32761, LUT_AMPL_WIDTH),
		16578 => to_signed(32761, LUT_AMPL_WIDTH),
		16579 => to_signed(32761, LUT_AMPL_WIDTH),
		16580 => to_signed(32761, LUT_AMPL_WIDTH),
		16581 => to_signed(32761, LUT_AMPL_WIDTH),
		16582 => to_signed(32761, LUT_AMPL_WIDTH),
		16583 => to_signed(32761, LUT_AMPL_WIDTH),
		16584 => to_signed(32761, LUT_AMPL_WIDTH),
		16585 => to_signed(32761, LUT_AMPL_WIDTH),
		16586 => to_signed(32761, LUT_AMPL_WIDTH),
		16587 => to_signed(32761, LUT_AMPL_WIDTH),
		16588 => to_signed(32761, LUT_AMPL_WIDTH),
		16589 => to_signed(32761, LUT_AMPL_WIDTH),
		16590 => to_signed(32761, LUT_AMPL_WIDTH),
		16591 => to_signed(32761, LUT_AMPL_WIDTH),
		16592 => to_signed(32760, LUT_AMPL_WIDTH),
		16593 => to_signed(32760, LUT_AMPL_WIDTH),
		16594 => to_signed(32760, LUT_AMPL_WIDTH),
		16595 => to_signed(32760, LUT_AMPL_WIDTH),
		16596 => to_signed(32760, LUT_AMPL_WIDTH),
		16597 => to_signed(32760, LUT_AMPL_WIDTH),
		16598 => to_signed(32760, LUT_AMPL_WIDTH),
		16599 => to_signed(32760, LUT_AMPL_WIDTH),
		16600 => to_signed(32760, LUT_AMPL_WIDTH),
		16601 => to_signed(32760, LUT_AMPL_WIDTH),
		16602 => to_signed(32760, LUT_AMPL_WIDTH),
		16603 => to_signed(32760, LUT_AMPL_WIDTH),
		16604 => to_signed(32760, LUT_AMPL_WIDTH),
		16605 => to_signed(32760, LUT_AMPL_WIDTH),
		16606 => to_signed(32760, LUT_AMPL_WIDTH),
		16607 => to_signed(32760, LUT_AMPL_WIDTH),
		16608 => to_signed(32759, LUT_AMPL_WIDTH),
		16609 => to_signed(32759, LUT_AMPL_WIDTH),
		16610 => to_signed(32759, LUT_AMPL_WIDTH),
		16611 => to_signed(32759, LUT_AMPL_WIDTH),
		16612 => to_signed(32759, LUT_AMPL_WIDTH),
		16613 => to_signed(32759, LUT_AMPL_WIDTH),
		16614 => to_signed(32759, LUT_AMPL_WIDTH),
		16615 => to_signed(32759, LUT_AMPL_WIDTH),
		16616 => to_signed(32759, LUT_AMPL_WIDTH),
		16617 => to_signed(32759, LUT_AMPL_WIDTH),
		16618 => to_signed(32759, LUT_AMPL_WIDTH),
		16619 => to_signed(32759, LUT_AMPL_WIDTH),
		16620 => to_signed(32759, LUT_AMPL_WIDTH),
		16621 => to_signed(32759, LUT_AMPL_WIDTH),
		16622 => to_signed(32758, LUT_AMPL_WIDTH),
		16623 => to_signed(32758, LUT_AMPL_WIDTH),
		16624 => to_signed(32758, LUT_AMPL_WIDTH),
		16625 => to_signed(32758, LUT_AMPL_WIDTH),
		16626 => to_signed(32758, LUT_AMPL_WIDTH),
		16627 => to_signed(32758, LUT_AMPL_WIDTH),
		16628 => to_signed(32758, LUT_AMPL_WIDTH),
		16629 => to_signed(32758, LUT_AMPL_WIDTH),
		16630 => to_signed(32758, LUT_AMPL_WIDTH),
		16631 => to_signed(32758, LUT_AMPL_WIDTH),
		16632 => to_signed(32758, LUT_AMPL_WIDTH),
		16633 => to_signed(32758, LUT_AMPL_WIDTH),
		16634 => to_signed(32758, LUT_AMPL_WIDTH),
		16635 => to_signed(32758, LUT_AMPL_WIDTH),
		16636 => to_signed(32757, LUT_AMPL_WIDTH),
		16637 => to_signed(32757, LUT_AMPL_WIDTH),
		16638 => to_signed(32757, LUT_AMPL_WIDTH),
		16639 => to_signed(32757, LUT_AMPL_WIDTH),
		16640 => to_signed(32757, LUT_AMPL_WIDTH),
		16641 => to_signed(32757, LUT_AMPL_WIDTH),
		16642 => to_signed(32757, LUT_AMPL_WIDTH),
		16643 => to_signed(32757, LUT_AMPL_WIDTH),
		16644 => to_signed(32757, LUT_AMPL_WIDTH),
		16645 => to_signed(32757, LUT_AMPL_WIDTH),
		16646 => to_signed(32757, LUT_AMPL_WIDTH),
		16647 => to_signed(32757, LUT_AMPL_WIDTH),
		16648 => to_signed(32757, LUT_AMPL_WIDTH),
		16649 => to_signed(32756, LUT_AMPL_WIDTH),
		16650 => to_signed(32756, LUT_AMPL_WIDTH),
		16651 => to_signed(32756, LUT_AMPL_WIDTH),
		16652 => to_signed(32756, LUT_AMPL_WIDTH),
		16653 => to_signed(32756, LUT_AMPL_WIDTH),
		16654 => to_signed(32756, LUT_AMPL_WIDTH),
		16655 => to_signed(32756, LUT_AMPL_WIDTH),
		16656 => to_signed(32756, LUT_AMPL_WIDTH),
		16657 => to_signed(32756, LUT_AMPL_WIDTH),
		16658 => to_signed(32756, LUT_AMPL_WIDTH),
		16659 => to_signed(32756, LUT_AMPL_WIDTH),
		16660 => to_signed(32756, LUT_AMPL_WIDTH),
		16661 => to_signed(32755, LUT_AMPL_WIDTH),
		16662 => to_signed(32755, LUT_AMPL_WIDTH),
		16663 => to_signed(32755, LUT_AMPL_WIDTH),
		16664 => to_signed(32755, LUT_AMPL_WIDTH),
		16665 => to_signed(32755, LUT_AMPL_WIDTH),
		16666 => to_signed(32755, LUT_AMPL_WIDTH),
		16667 => to_signed(32755, LUT_AMPL_WIDTH),
		16668 => to_signed(32755, LUT_AMPL_WIDTH),
		16669 => to_signed(32755, LUT_AMPL_WIDTH),
		16670 => to_signed(32755, LUT_AMPL_WIDTH),
		16671 => to_signed(32755, LUT_AMPL_WIDTH),
		16672 => to_signed(32755, LUT_AMPL_WIDTH),
		16673 => to_signed(32754, LUT_AMPL_WIDTH),
		16674 => to_signed(32754, LUT_AMPL_WIDTH),
		16675 => to_signed(32754, LUT_AMPL_WIDTH),
		16676 => to_signed(32754, LUT_AMPL_WIDTH),
		16677 => to_signed(32754, LUT_AMPL_WIDTH),
		16678 => to_signed(32754, LUT_AMPL_WIDTH),
		16679 => to_signed(32754, LUT_AMPL_WIDTH),
		16680 => to_signed(32754, LUT_AMPL_WIDTH),
		16681 => to_signed(32754, LUT_AMPL_WIDTH),
		16682 => to_signed(32754, LUT_AMPL_WIDTH),
		16683 => to_signed(32754, LUT_AMPL_WIDTH),
		16684 => to_signed(32753, LUT_AMPL_WIDTH),
		16685 => to_signed(32753, LUT_AMPL_WIDTH),
		16686 => to_signed(32753, LUT_AMPL_WIDTH),
		16687 => to_signed(32753, LUT_AMPL_WIDTH),
		16688 => to_signed(32753, LUT_AMPL_WIDTH),
		16689 => to_signed(32753, LUT_AMPL_WIDTH),
		16690 => to_signed(32753, LUT_AMPL_WIDTH),
		16691 => to_signed(32753, LUT_AMPL_WIDTH),
		16692 => to_signed(32753, LUT_AMPL_WIDTH),
		16693 => to_signed(32753, LUT_AMPL_WIDTH),
		16694 => to_signed(32753, LUT_AMPL_WIDTH),
		16695 => to_signed(32752, LUT_AMPL_WIDTH),
		16696 => to_signed(32752, LUT_AMPL_WIDTH),
		16697 => to_signed(32752, LUT_AMPL_WIDTH),
		16698 => to_signed(32752, LUT_AMPL_WIDTH),
		16699 => to_signed(32752, LUT_AMPL_WIDTH),
		16700 => to_signed(32752, LUT_AMPL_WIDTH),
		16701 => to_signed(32752, LUT_AMPL_WIDTH),
		16702 => to_signed(32752, LUT_AMPL_WIDTH),
		16703 => to_signed(32752, LUT_AMPL_WIDTH),
		16704 => to_signed(32752, LUT_AMPL_WIDTH),
		16705 => to_signed(32751, LUT_AMPL_WIDTH),
		16706 => to_signed(32751, LUT_AMPL_WIDTH),
		16707 => to_signed(32751, LUT_AMPL_WIDTH),
		16708 => to_signed(32751, LUT_AMPL_WIDTH),
		16709 => to_signed(32751, LUT_AMPL_WIDTH),
		16710 => to_signed(32751, LUT_AMPL_WIDTH),
		16711 => to_signed(32751, LUT_AMPL_WIDTH),
		16712 => to_signed(32751, LUT_AMPL_WIDTH),
		16713 => to_signed(32751, LUT_AMPL_WIDTH),
		16714 => to_signed(32751, LUT_AMPL_WIDTH),
		16715 => to_signed(32751, LUT_AMPL_WIDTH),
		16716 => to_signed(32750, LUT_AMPL_WIDTH),
		16717 => to_signed(32750, LUT_AMPL_WIDTH),
		16718 => to_signed(32750, LUT_AMPL_WIDTH),
		16719 => to_signed(32750, LUT_AMPL_WIDTH),
		16720 => to_signed(32750, LUT_AMPL_WIDTH),
		16721 => to_signed(32750, LUT_AMPL_WIDTH),
		16722 => to_signed(32750, LUT_AMPL_WIDTH),
		16723 => to_signed(32750, LUT_AMPL_WIDTH),
		16724 => to_signed(32750, LUT_AMPL_WIDTH),
		16725 => to_signed(32749, LUT_AMPL_WIDTH),
		16726 => to_signed(32749, LUT_AMPL_WIDTH),
		16727 => to_signed(32749, LUT_AMPL_WIDTH),
		16728 => to_signed(32749, LUT_AMPL_WIDTH),
		16729 => to_signed(32749, LUT_AMPL_WIDTH),
		16730 => to_signed(32749, LUT_AMPL_WIDTH),
		16731 => to_signed(32749, LUT_AMPL_WIDTH),
		16732 => to_signed(32749, LUT_AMPL_WIDTH),
		16733 => to_signed(32749, LUT_AMPL_WIDTH),
		16734 => to_signed(32749, LUT_AMPL_WIDTH),
		16735 => to_signed(32748, LUT_AMPL_WIDTH),
		16736 => to_signed(32748, LUT_AMPL_WIDTH),
		16737 => to_signed(32748, LUT_AMPL_WIDTH),
		16738 => to_signed(32748, LUT_AMPL_WIDTH),
		16739 => to_signed(32748, LUT_AMPL_WIDTH),
		16740 => to_signed(32748, LUT_AMPL_WIDTH),
		16741 => to_signed(32748, LUT_AMPL_WIDTH),
		16742 => to_signed(32748, LUT_AMPL_WIDTH),
		16743 => to_signed(32748, LUT_AMPL_WIDTH),
		16744 => to_signed(32747, LUT_AMPL_WIDTH),
		16745 => to_signed(32747, LUT_AMPL_WIDTH),
		16746 => to_signed(32747, LUT_AMPL_WIDTH),
		16747 => to_signed(32747, LUT_AMPL_WIDTH),
		16748 => to_signed(32747, LUT_AMPL_WIDTH),
		16749 => to_signed(32747, LUT_AMPL_WIDTH),
		16750 => to_signed(32747, LUT_AMPL_WIDTH),
		16751 => to_signed(32747, LUT_AMPL_WIDTH),
		16752 => to_signed(32747, LUT_AMPL_WIDTH),
		16753 => to_signed(32746, LUT_AMPL_WIDTH),
		16754 => to_signed(32746, LUT_AMPL_WIDTH),
		16755 => to_signed(32746, LUT_AMPL_WIDTH),
		16756 => to_signed(32746, LUT_AMPL_WIDTH),
		16757 => to_signed(32746, LUT_AMPL_WIDTH),
		16758 => to_signed(32746, LUT_AMPL_WIDTH),
		16759 => to_signed(32746, LUT_AMPL_WIDTH),
		16760 => to_signed(32746, LUT_AMPL_WIDTH),
		16761 => to_signed(32746, LUT_AMPL_WIDTH),
		16762 => to_signed(32745, LUT_AMPL_WIDTH),
		16763 => to_signed(32745, LUT_AMPL_WIDTH),
		16764 => to_signed(32745, LUT_AMPL_WIDTH),
		16765 => to_signed(32745, LUT_AMPL_WIDTH),
		16766 => to_signed(32745, LUT_AMPL_WIDTH),
		16767 => to_signed(32745, LUT_AMPL_WIDTH),
		16768 => to_signed(32745, LUT_AMPL_WIDTH),
		16769 => to_signed(32745, LUT_AMPL_WIDTH),
		16770 => to_signed(32745, LUT_AMPL_WIDTH),
		16771 => to_signed(32744, LUT_AMPL_WIDTH),
		16772 => to_signed(32744, LUT_AMPL_WIDTH),
		16773 => to_signed(32744, LUT_AMPL_WIDTH),
		16774 => to_signed(32744, LUT_AMPL_WIDTH),
		16775 => to_signed(32744, LUT_AMPL_WIDTH),
		16776 => to_signed(32744, LUT_AMPL_WIDTH),
		16777 => to_signed(32744, LUT_AMPL_WIDTH),
		16778 => to_signed(32744, LUT_AMPL_WIDTH),
		16779 => to_signed(32744, LUT_AMPL_WIDTH),
		16780 => to_signed(32743, LUT_AMPL_WIDTH),
		16781 => to_signed(32743, LUT_AMPL_WIDTH),
		16782 => to_signed(32743, LUT_AMPL_WIDTH),
		16783 => to_signed(32743, LUT_AMPL_WIDTH),
		16784 => to_signed(32743, LUT_AMPL_WIDTH),
		16785 => to_signed(32743, LUT_AMPL_WIDTH),
		16786 => to_signed(32743, LUT_AMPL_WIDTH),
		16787 => to_signed(32743, LUT_AMPL_WIDTH),
		16788 => to_signed(32742, LUT_AMPL_WIDTH),
		16789 => to_signed(32742, LUT_AMPL_WIDTH),
		16790 => to_signed(32742, LUT_AMPL_WIDTH),
		16791 => to_signed(32742, LUT_AMPL_WIDTH),
		16792 => to_signed(32742, LUT_AMPL_WIDTH),
		16793 => to_signed(32742, LUT_AMPL_WIDTH),
		16794 => to_signed(32742, LUT_AMPL_WIDTH),
		16795 => to_signed(32742, LUT_AMPL_WIDTH),
		16796 => to_signed(32741, LUT_AMPL_WIDTH),
		16797 => to_signed(32741, LUT_AMPL_WIDTH),
		16798 => to_signed(32741, LUT_AMPL_WIDTH),
		16799 => to_signed(32741, LUT_AMPL_WIDTH),
		16800 => to_signed(32741, LUT_AMPL_WIDTH),
		16801 => to_signed(32741, LUT_AMPL_WIDTH),
		16802 => to_signed(32741, LUT_AMPL_WIDTH),
		16803 => to_signed(32741, LUT_AMPL_WIDTH),
		16804 => to_signed(32740, LUT_AMPL_WIDTH),
		16805 => to_signed(32740, LUT_AMPL_WIDTH),
		16806 => to_signed(32740, LUT_AMPL_WIDTH),
		16807 => to_signed(32740, LUT_AMPL_WIDTH),
		16808 => to_signed(32740, LUT_AMPL_WIDTH),
		16809 => to_signed(32740, LUT_AMPL_WIDTH),
		16810 => to_signed(32740, LUT_AMPL_WIDTH),
		16811 => to_signed(32740, LUT_AMPL_WIDTH),
		16812 => to_signed(32739, LUT_AMPL_WIDTH),
		16813 => to_signed(32739, LUT_AMPL_WIDTH),
		16814 => to_signed(32739, LUT_AMPL_WIDTH),
		16815 => to_signed(32739, LUT_AMPL_WIDTH),
		16816 => to_signed(32739, LUT_AMPL_WIDTH),
		16817 => to_signed(32739, LUT_AMPL_WIDTH),
		16818 => to_signed(32739, LUT_AMPL_WIDTH),
		16819 => to_signed(32739, LUT_AMPL_WIDTH),
		16820 => to_signed(32738, LUT_AMPL_WIDTH),
		16821 => to_signed(32738, LUT_AMPL_WIDTH),
		16822 => to_signed(32738, LUT_AMPL_WIDTH),
		16823 => to_signed(32738, LUT_AMPL_WIDTH),
		16824 => to_signed(32738, LUT_AMPL_WIDTH),
		16825 => to_signed(32738, LUT_AMPL_WIDTH),
		16826 => to_signed(32738, LUT_AMPL_WIDTH),
		16827 => to_signed(32737, LUT_AMPL_WIDTH),
		16828 => to_signed(32737, LUT_AMPL_WIDTH),
		16829 => to_signed(32737, LUT_AMPL_WIDTH),
		16830 => to_signed(32737, LUT_AMPL_WIDTH),
		16831 => to_signed(32737, LUT_AMPL_WIDTH),
		16832 => to_signed(32737, LUT_AMPL_WIDTH),
		16833 => to_signed(32737, LUT_AMPL_WIDTH),
		16834 => to_signed(32737, LUT_AMPL_WIDTH),
		16835 => to_signed(32736, LUT_AMPL_WIDTH),
		16836 => to_signed(32736, LUT_AMPL_WIDTH),
		16837 => to_signed(32736, LUT_AMPL_WIDTH),
		16838 => to_signed(32736, LUT_AMPL_WIDTH),
		16839 => to_signed(32736, LUT_AMPL_WIDTH),
		16840 => to_signed(32736, LUT_AMPL_WIDTH),
		16841 => to_signed(32736, LUT_AMPL_WIDTH),
		16842 => to_signed(32735, LUT_AMPL_WIDTH),
		16843 => to_signed(32735, LUT_AMPL_WIDTH),
		16844 => to_signed(32735, LUT_AMPL_WIDTH),
		16845 => to_signed(32735, LUT_AMPL_WIDTH),
		16846 => to_signed(32735, LUT_AMPL_WIDTH),
		16847 => to_signed(32735, LUT_AMPL_WIDTH),
		16848 => to_signed(32735, LUT_AMPL_WIDTH),
		16849 => to_signed(32734, LUT_AMPL_WIDTH),
		16850 => to_signed(32734, LUT_AMPL_WIDTH),
		16851 => to_signed(32734, LUT_AMPL_WIDTH),
		16852 => to_signed(32734, LUT_AMPL_WIDTH),
		16853 => to_signed(32734, LUT_AMPL_WIDTH),
		16854 => to_signed(32734, LUT_AMPL_WIDTH),
		16855 => to_signed(32734, LUT_AMPL_WIDTH),
		16856 => to_signed(32733, LUT_AMPL_WIDTH),
		16857 => to_signed(32733, LUT_AMPL_WIDTH),
		16858 => to_signed(32733, LUT_AMPL_WIDTH),
		16859 => to_signed(32733, LUT_AMPL_WIDTH),
		16860 => to_signed(32733, LUT_AMPL_WIDTH),
		16861 => to_signed(32733, LUT_AMPL_WIDTH),
		16862 => to_signed(32733, LUT_AMPL_WIDTH),
		16863 => to_signed(32732, LUT_AMPL_WIDTH),
		16864 => to_signed(32732, LUT_AMPL_WIDTH),
		16865 => to_signed(32732, LUT_AMPL_WIDTH),
		16866 => to_signed(32732, LUT_AMPL_WIDTH),
		16867 => to_signed(32732, LUT_AMPL_WIDTH),
		16868 => to_signed(32732, LUT_AMPL_WIDTH),
		16869 => to_signed(32732, LUT_AMPL_WIDTH),
		16870 => to_signed(32731, LUT_AMPL_WIDTH),
		16871 => to_signed(32731, LUT_AMPL_WIDTH),
		16872 => to_signed(32731, LUT_AMPL_WIDTH),
		16873 => to_signed(32731, LUT_AMPL_WIDTH),
		16874 => to_signed(32731, LUT_AMPL_WIDTH),
		16875 => to_signed(32731, LUT_AMPL_WIDTH),
		16876 => to_signed(32731, LUT_AMPL_WIDTH),
		16877 => to_signed(32730, LUT_AMPL_WIDTH),
		16878 => to_signed(32730, LUT_AMPL_WIDTH),
		16879 => to_signed(32730, LUT_AMPL_WIDTH),
		16880 => to_signed(32730, LUT_AMPL_WIDTH),
		16881 => to_signed(32730, LUT_AMPL_WIDTH),
		16882 => to_signed(32730, LUT_AMPL_WIDTH),
		16883 => to_signed(32730, LUT_AMPL_WIDTH),
		16884 => to_signed(32729, LUT_AMPL_WIDTH),
		16885 => to_signed(32729, LUT_AMPL_WIDTH),
		16886 => to_signed(32729, LUT_AMPL_WIDTH),
		16887 => to_signed(32729, LUT_AMPL_WIDTH),
		16888 => to_signed(32729, LUT_AMPL_WIDTH),
		16889 => to_signed(32729, LUT_AMPL_WIDTH),
		16890 => to_signed(32728, LUT_AMPL_WIDTH),
		16891 => to_signed(32728, LUT_AMPL_WIDTH),
		16892 => to_signed(32728, LUT_AMPL_WIDTH),
		16893 => to_signed(32728, LUT_AMPL_WIDTH),
		16894 => to_signed(32728, LUT_AMPL_WIDTH),
		16895 => to_signed(32728, LUT_AMPL_WIDTH),
		16896 => to_signed(32728, LUT_AMPL_WIDTH),
		16897 => to_signed(32727, LUT_AMPL_WIDTH),
		16898 => to_signed(32727, LUT_AMPL_WIDTH),
		16899 => to_signed(32727, LUT_AMPL_WIDTH),
		16900 => to_signed(32727, LUT_AMPL_WIDTH),
		16901 => to_signed(32727, LUT_AMPL_WIDTH),
		16902 => to_signed(32727, LUT_AMPL_WIDTH),
		16903 => to_signed(32726, LUT_AMPL_WIDTH),
		16904 => to_signed(32726, LUT_AMPL_WIDTH),
		16905 => to_signed(32726, LUT_AMPL_WIDTH),
		16906 => to_signed(32726, LUT_AMPL_WIDTH),
		16907 => to_signed(32726, LUT_AMPL_WIDTH),
		16908 => to_signed(32726, LUT_AMPL_WIDTH),
		16909 => to_signed(32726, LUT_AMPL_WIDTH),
		16910 => to_signed(32725, LUT_AMPL_WIDTH),
		16911 => to_signed(32725, LUT_AMPL_WIDTH),
		16912 => to_signed(32725, LUT_AMPL_WIDTH),
		16913 => to_signed(32725, LUT_AMPL_WIDTH),
		16914 => to_signed(32725, LUT_AMPL_WIDTH),
		16915 => to_signed(32725, LUT_AMPL_WIDTH),
		16916 => to_signed(32724, LUT_AMPL_WIDTH),
		16917 => to_signed(32724, LUT_AMPL_WIDTH),
		16918 => to_signed(32724, LUT_AMPL_WIDTH),
		16919 => to_signed(32724, LUT_AMPL_WIDTH),
		16920 => to_signed(32724, LUT_AMPL_WIDTH),
		16921 => to_signed(32724, LUT_AMPL_WIDTH),
		16922 => to_signed(32723, LUT_AMPL_WIDTH),
		16923 => to_signed(32723, LUT_AMPL_WIDTH),
		16924 => to_signed(32723, LUT_AMPL_WIDTH),
		16925 => to_signed(32723, LUT_AMPL_WIDTH),
		16926 => to_signed(32723, LUT_AMPL_WIDTH),
		16927 => to_signed(32723, LUT_AMPL_WIDTH),
		16928 => to_signed(32722, LUT_AMPL_WIDTH),
		16929 => to_signed(32722, LUT_AMPL_WIDTH),
		16930 => to_signed(32722, LUT_AMPL_WIDTH),
		16931 => to_signed(32722, LUT_AMPL_WIDTH),
		16932 => to_signed(32722, LUT_AMPL_WIDTH),
		16933 => to_signed(32722, LUT_AMPL_WIDTH),
		16934 => to_signed(32721, LUT_AMPL_WIDTH),
		16935 => to_signed(32721, LUT_AMPL_WIDTH),
		16936 => to_signed(32721, LUT_AMPL_WIDTH),
		16937 => to_signed(32721, LUT_AMPL_WIDTH),
		16938 => to_signed(32721, LUT_AMPL_WIDTH),
		16939 => to_signed(32721, LUT_AMPL_WIDTH),
		16940 => to_signed(32720, LUT_AMPL_WIDTH),
		16941 => to_signed(32720, LUT_AMPL_WIDTH),
		16942 => to_signed(32720, LUT_AMPL_WIDTH),
		16943 => to_signed(32720, LUT_AMPL_WIDTH),
		16944 => to_signed(32720, LUT_AMPL_WIDTH),
		16945 => to_signed(32720, LUT_AMPL_WIDTH),
		16946 => to_signed(32719, LUT_AMPL_WIDTH),
		16947 => to_signed(32719, LUT_AMPL_WIDTH),
		16948 => to_signed(32719, LUT_AMPL_WIDTH),
		16949 => to_signed(32719, LUT_AMPL_WIDTH),
		16950 => to_signed(32719, LUT_AMPL_WIDTH),
		16951 => to_signed(32719, LUT_AMPL_WIDTH),
		16952 => to_signed(32718, LUT_AMPL_WIDTH),
		16953 => to_signed(32718, LUT_AMPL_WIDTH),
		16954 => to_signed(32718, LUT_AMPL_WIDTH),
		16955 => to_signed(32718, LUT_AMPL_WIDTH),
		16956 => to_signed(32718, LUT_AMPL_WIDTH),
		16957 => to_signed(32718, LUT_AMPL_WIDTH),
		16958 => to_signed(32717, LUT_AMPL_WIDTH),
		16959 => to_signed(32717, LUT_AMPL_WIDTH),
		16960 => to_signed(32717, LUT_AMPL_WIDTH),
		16961 => to_signed(32717, LUT_AMPL_WIDTH),
		16962 => to_signed(32717, LUT_AMPL_WIDTH),
		16963 => to_signed(32717, LUT_AMPL_WIDTH),
		16964 => to_signed(32716, LUT_AMPL_WIDTH),
		16965 => to_signed(32716, LUT_AMPL_WIDTH),
		16966 => to_signed(32716, LUT_AMPL_WIDTH),
		16967 => to_signed(32716, LUT_AMPL_WIDTH),
		16968 => to_signed(32716, LUT_AMPL_WIDTH),
		16969 => to_signed(32715, LUT_AMPL_WIDTH),
		16970 => to_signed(32715, LUT_AMPL_WIDTH),
		16971 => to_signed(32715, LUT_AMPL_WIDTH),
		16972 => to_signed(32715, LUT_AMPL_WIDTH),
		16973 => to_signed(32715, LUT_AMPL_WIDTH),
		16974 => to_signed(32715, LUT_AMPL_WIDTH),
		16975 => to_signed(32714, LUT_AMPL_WIDTH),
		16976 => to_signed(32714, LUT_AMPL_WIDTH),
		16977 => to_signed(32714, LUT_AMPL_WIDTH),
		16978 => to_signed(32714, LUT_AMPL_WIDTH),
		16979 => to_signed(32714, LUT_AMPL_WIDTH),
		16980 => to_signed(32714, LUT_AMPL_WIDTH),
		16981 => to_signed(32713, LUT_AMPL_WIDTH),
		16982 => to_signed(32713, LUT_AMPL_WIDTH),
		16983 => to_signed(32713, LUT_AMPL_WIDTH),
		16984 => to_signed(32713, LUT_AMPL_WIDTH),
		16985 => to_signed(32713, LUT_AMPL_WIDTH),
		16986 => to_signed(32712, LUT_AMPL_WIDTH),
		16987 => to_signed(32712, LUT_AMPL_WIDTH),
		16988 => to_signed(32712, LUT_AMPL_WIDTH),
		16989 => to_signed(32712, LUT_AMPL_WIDTH),
		16990 => to_signed(32712, LUT_AMPL_WIDTH),
		16991 => to_signed(32712, LUT_AMPL_WIDTH),
		16992 => to_signed(32711, LUT_AMPL_WIDTH),
		16993 => to_signed(32711, LUT_AMPL_WIDTH),
		16994 => to_signed(32711, LUT_AMPL_WIDTH),
		16995 => to_signed(32711, LUT_AMPL_WIDTH),
		16996 => to_signed(32711, LUT_AMPL_WIDTH),
		16997 => to_signed(32710, LUT_AMPL_WIDTH),
		16998 => to_signed(32710, LUT_AMPL_WIDTH),
		16999 => to_signed(32710, LUT_AMPL_WIDTH),
		17000 => to_signed(32710, LUT_AMPL_WIDTH),
		17001 => to_signed(32710, LUT_AMPL_WIDTH),
		17002 => to_signed(32710, LUT_AMPL_WIDTH),
		17003 => to_signed(32709, LUT_AMPL_WIDTH),
		17004 => to_signed(32709, LUT_AMPL_WIDTH),
		17005 => to_signed(32709, LUT_AMPL_WIDTH),
		17006 => to_signed(32709, LUT_AMPL_WIDTH),
		17007 => to_signed(32709, LUT_AMPL_WIDTH),
		17008 => to_signed(32708, LUT_AMPL_WIDTH),
		17009 => to_signed(32708, LUT_AMPL_WIDTH),
		17010 => to_signed(32708, LUT_AMPL_WIDTH),
		17011 => to_signed(32708, LUT_AMPL_WIDTH),
		17012 => to_signed(32708, LUT_AMPL_WIDTH),
		17013 => to_signed(32707, LUT_AMPL_WIDTH),
		17014 => to_signed(32707, LUT_AMPL_WIDTH),
		17015 => to_signed(32707, LUT_AMPL_WIDTH),
		17016 => to_signed(32707, LUT_AMPL_WIDTH),
		17017 => to_signed(32707, LUT_AMPL_WIDTH),
		17018 => to_signed(32706, LUT_AMPL_WIDTH),
		17019 => to_signed(32706, LUT_AMPL_WIDTH),
		17020 => to_signed(32706, LUT_AMPL_WIDTH),
		17021 => to_signed(32706, LUT_AMPL_WIDTH),
		17022 => to_signed(32706, LUT_AMPL_WIDTH),
		17023 => to_signed(32706, LUT_AMPL_WIDTH),
		17024 => to_signed(32705, LUT_AMPL_WIDTH),
		17025 => to_signed(32705, LUT_AMPL_WIDTH),
		17026 => to_signed(32705, LUT_AMPL_WIDTH),
		17027 => to_signed(32705, LUT_AMPL_WIDTH),
		17028 => to_signed(32705, LUT_AMPL_WIDTH),
		17029 => to_signed(32704, LUT_AMPL_WIDTH),
		17030 => to_signed(32704, LUT_AMPL_WIDTH),
		17031 => to_signed(32704, LUT_AMPL_WIDTH),
		17032 => to_signed(32704, LUT_AMPL_WIDTH),
		17033 => to_signed(32704, LUT_AMPL_WIDTH),
		17034 => to_signed(32703, LUT_AMPL_WIDTH),
		17035 => to_signed(32703, LUT_AMPL_WIDTH),
		17036 => to_signed(32703, LUT_AMPL_WIDTH),
		17037 => to_signed(32703, LUT_AMPL_WIDTH),
		17038 => to_signed(32703, LUT_AMPL_WIDTH),
		17039 => to_signed(32702, LUT_AMPL_WIDTH),
		17040 => to_signed(32702, LUT_AMPL_WIDTH),
		17041 => to_signed(32702, LUT_AMPL_WIDTH),
		17042 => to_signed(32702, LUT_AMPL_WIDTH),
		17043 => to_signed(32702, LUT_AMPL_WIDTH),
		17044 => to_signed(32701, LUT_AMPL_WIDTH),
		17045 => to_signed(32701, LUT_AMPL_WIDTH),
		17046 => to_signed(32701, LUT_AMPL_WIDTH),
		17047 => to_signed(32701, LUT_AMPL_WIDTH),
		17048 => to_signed(32701, LUT_AMPL_WIDTH),
		17049 => to_signed(32700, LUT_AMPL_WIDTH),
		17050 => to_signed(32700, LUT_AMPL_WIDTH),
		17051 => to_signed(32700, LUT_AMPL_WIDTH),
		17052 => to_signed(32700, LUT_AMPL_WIDTH),
		17053 => to_signed(32700, LUT_AMPL_WIDTH),
		17054 => to_signed(32699, LUT_AMPL_WIDTH),
		17055 => to_signed(32699, LUT_AMPL_WIDTH),
		17056 => to_signed(32699, LUT_AMPL_WIDTH),
		17057 => to_signed(32699, LUT_AMPL_WIDTH),
		17058 => to_signed(32699, LUT_AMPL_WIDTH),
		17059 => to_signed(32698, LUT_AMPL_WIDTH),
		17060 => to_signed(32698, LUT_AMPL_WIDTH),
		17061 => to_signed(32698, LUT_AMPL_WIDTH),
		17062 => to_signed(32698, LUT_AMPL_WIDTH),
		17063 => to_signed(32698, LUT_AMPL_WIDTH),
		17064 => to_signed(32697, LUT_AMPL_WIDTH),
		17065 => to_signed(32697, LUT_AMPL_WIDTH),
		17066 => to_signed(32697, LUT_AMPL_WIDTH),
		17067 => to_signed(32697, LUT_AMPL_WIDTH),
		17068 => to_signed(32697, LUT_AMPL_WIDTH),
		17069 => to_signed(32696, LUT_AMPL_WIDTH),
		17070 => to_signed(32696, LUT_AMPL_WIDTH),
		17071 => to_signed(32696, LUT_AMPL_WIDTH),
		17072 => to_signed(32696, LUT_AMPL_WIDTH),
		17073 => to_signed(32696, LUT_AMPL_WIDTH),
		17074 => to_signed(32695, LUT_AMPL_WIDTH),
		17075 => to_signed(32695, LUT_AMPL_WIDTH),
		17076 => to_signed(32695, LUT_AMPL_WIDTH),
		17077 => to_signed(32695, LUT_AMPL_WIDTH),
		17078 => to_signed(32694, LUT_AMPL_WIDTH),
		17079 => to_signed(32694, LUT_AMPL_WIDTH),
		17080 => to_signed(32694, LUT_AMPL_WIDTH),
		17081 => to_signed(32694, LUT_AMPL_WIDTH),
		17082 => to_signed(32694, LUT_AMPL_WIDTH),
		17083 => to_signed(32693, LUT_AMPL_WIDTH),
		17084 => to_signed(32693, LUT_AMPL_WIDTH),
		17085 => to_signed(32693, LUT_AMPL_WIDTH),
		17086 => to_signed(32693, LUT_AMPL_WIDTH),
		17087 => to_signed(32693, LUT_AMPL_WIDTH),
		17088 => to_signed(32692, LUT_AMPL_WIDTH),
		17089 => to_signed(32692, LUT_AMPL_WIDTH),
		17090 => to_signed(32692, LUT_AMPL_WIDTH),
		17091 => to_signed(32692, LUT_AMPL_WIDTH),
		17092 => to_signed(32692, LUT_AMPL_WIDTH),
		17093 => to_signed(32691, LUT_AMPL_WIDTH),
		17094 => to_signed(32691, LUT_AMPL_WIDTH),
		17095 => to_signed(32691, LUT_AMPL_WIDTH),
		17096 => to_signed(32691, LUT_AMPL_WIDTH),
		17097 => to_signed(32690, LUT_AMPL_WIDTH),
		17098 => to_signed(32690, LUT_AMPL_WIDTH),
		17099 => to_signed(32690, LUT_AMPL_WIDTH),
		17100 => to_signed(32690, LUT_AMPL_WIDTH),
		17101 => to_signed(32690, LUT_AMPL_WIDTH),
		17102 => to_signed(32689, LUT_AMPL_WIDTH),
		17103 => to_signed(32689, LUT_AMPL_WIDTH),
		17104 => to_signed(32689, LUT_AMPL_WIDTH),
		17105 => to_signed(32689, LUT_AMPL_WIDTH),
		17106 => to_signed(32689, LUT_AMPL_WIDTH),
		17107 => to_signed(32688, LUT_AMPL_WIDTH),
		17108 => to_signed(32688, LUT_AMPL_WIDTH),
		17109 => to_signed(32688, LUT_AMPL_WIDTH),
		17110 => to_signed(32688, LUT_AMPL_WIDTH),
		17111 => to_signed(32687, LUT_AMPL_WIDTH),
		17112 => to_signed(32687, LUT_AMPL_WIDTH),
		17113 => to_signed(32687, LUT_AMPL_WIDTH),
		17114 => to_signed(32687, LUT_AMPL_WIDTH),
		17115 => to_signed(32687, LUT_AMPL_WIDTH),
		17116 => to_signed(32686, LUT_AMPL_WIDTH),
		17117 => to_signed(32686, LUT_AMPL_WIDTH),
		17118 => to_signed(32686, LUT_AMPL_WIDTH),
		17119 => to_signed(32686, LUT_AMPL_WIDTH),
		17120 => to_signed(32685, LUT_AMPL_WIDTH),
		17121 => to_signed(32685, LUT_AMPL_WIDTH),
		17122 => to_signed(32685, LUT_AMPL_WIDTH),
		17123 => to_signed(32685, LUT_AMPL_WIDTH),
		17124 => to_signed(32685, LUT_AMPL_WIDTH),
		17125 => to_signed(32684, LUT_AMPL_WIDTH),
		17126 => to_signed(32684, LUT_AMPL_WIDTH),
		17127 => to_signed(32684, LUT_AMPL_WIDTH),
		17128 => to_signed(32684, LUT_AMPL_WIDTH),
		17129 => to_signed(32683, LUT_AMPL_WIDTH),
		17130 => to_signed(32683, LUT_AMPL_WIDTH),
		17131 => to_signed(32683, LUT_AMPL_WIDTH),
		17132 => to_signed(32683, LUT_AMPL_WIDTH),
		17133 => to_signed(32683, LUT_AMPL_WIDTH),
		17134 => to_signed(32682, LUT_AMPL_WIDTH),
		17135 => to_signed(32682, LUT_AMPL_WIDTH),
		17136 => to_signed(32682, LUT_AMPL_WIDTH),
		17137 => to_signed(32682, LUT_AMPL_WIDTH),
		17138 => to_signed(32681, LUT_AMPL_WIDTH),
		17139 => to_signed(32681, LUT_AMPL_WIDTH),
		17140 => to_signed(32681, LUT_AMPL_WIDTH),
		17141 => to_signed(32681, LUT_AMPL_WIDTH),
		17142 => to_signed(32681, LUT_AMPL_WIDTH),
		17143 => to_signed(32680, LUT_AMPL_WIDTH),
		17144 => to_signed(32680, LUT_AMPL_WIDTH),
		17145 => to_signed(32680, LUT_AMPL_WIDTH),
		17146 => to_signed(32680, LUT_AMPL_WIDTH),
		17147 => to_signed(32679, LUT_AMPL_WIDTH),
		17148 => to_signed(32679, LUT_AMPL_WIDTH),
		17149 => to_signed(32679, LUT_AMPL_WIDTH),
		17150 => to_signed(32679, LUT_AMPL_WIDTH),
		17151 => to_signed(32678, LUT_AMPL_WIDTH),
		17152 => to_signed(32678, LUT_AMPL_WIDTH),
		17153 => to_signed(32678, LUT_AMPL_WIDTH),
		17154 => to_signed(32678, LUT_AMPL_WIDTH),
		17155 => to_signed(32678, LUT_AMPL_WIDTH),
		17156 => to_signed(32677, LUT_AMPL_WIDTH),
		17157 => to_signed(32677, LUT_AMPL_WIDTH),
		17158 => to_signed(32677, LUT_AMPL_WIDTH),
		17159 => to_signed(32677, LUT_AMPL_WIDTH),
		17160 => to_signed(32676, LUT_AMPL_WIDTH),
		17161 => to_signed(32676, LUT_AMPL_WIDTH),
		17162 => to_signed(32676, LUT_AMPL_WIDTH),
		17163 => to_signed(32676, LUT_AMPL_WIDTH),
		17164 => to_signed(32675, LUT_AMPL_WIDTH),
		17165 => to_signed(32675, LUT_AMPL_WIDTH),
		17166 => to_signed(32675, LUT_AMPL_WIDTH),
		17167 => to_signed(32675, LUT_AMPL_WIDTH),
		17168 => to_signed(32674, LUT_AMPL_WIDTH),
		17169 => to_signed(32674, LUT_AMPL_WIDTH),
		17170 => to_signed(32674, LUT_AMPL_WIDTH),
		17171 => to_signed(32674, LUT_AMPL_WIDTH),
		17172 => to_signed(32674, LUT_AMPL_WIDTH),
		17173 => to_signed(32673, LUT_AMPL_WIDTH),
		17174 => to_signed(32673, LUT_AMPL_WIDTH),
		17175 => to_signed(32673, LUT_AMPL_WIDTH),
		17176 => to_signed(32673, LUT_AMPL_WIDTH),
		17177 => to_signed(32672, LUT_AMPL_WIDTH),
		17178 => to_signed(32672, LUT_AMPL_WIDTH),
		17179 => to_signed(32672, LUT_AMPL_WIDTH),
		17180 => to_signed(32672, LUT_AMPL_WIDTH),
		17181 => to_signed(32671, LUT_AMPL_WIDTH),
		17182 => to_signed(32671, LUT_AMPL_WIDTH),
		17183 => to_signed(32671, LUT_AMPL_WIDTH),
		17184 => to_signed(32671, LUT_AMPL_WIDTH),
		17185 => to_signed(32670, LUT_AMPL_WIDTH),
		17186 => to_signed(32670, LUT_AMPL_WIDTH),
		17187 => to_signed(32670, LUT_AMPL_WIDTH),
		17188 => to_signed(32670, LUT_AMPL_WIDTH),
		17189 => to_signed(32669, LUT_AMPL_WIDTH),
		17190 => to_signed(32669, LUT_AMPL_WIDTH),
		17191 => to_signed(32669, LUT_AMPL_WIDTH),
		17192 => to_signed(32669, LUT_AMPL_WIDTH),
		17193 => to_signed(32668, LUT_AMPL_WIDTH),
		17194 => to_signed(32668, LUT_AMPL_WIDTH),
		17195 => to_signed(32668, LUT_AMPL_WIDTH),
		17196 => to_signed(32668, LUT_AMPL_WIDTH),
		17197 => to_signed(32668, LUT_AMPL_WIDTH),
		17198 => to_signed(32667, LUT_AMPL_WIDTH),
		17199 => to_signed(32667, LUT_AMPL_WIDTH),
		17200 => to_signed(32667, LUT_AMPL_WIDTH),
		17201 => to_signed(32667, LUT_AMPL_WIDTH),
		17202 => to_signed(32666, LUT_AMPL_WIDTH),
		17203 => to_signed(32666, LUT_AMPL_WIDTH),
		17204 => to_signed(32666, LUT_AMPL_WIDTH),
		17205 => to_signed(32666, LUT_AMPL_WIDTH),
		17206 => to_signed(32665, LUT_AMPL_WIDTH),
		17207 => to_signed(32665, LUT_AMPL_WIDTH),
		17208 => to_signed(32665, LUT_AMPL_WIDTH),
		17209 => to_signed(32665, LUT_AMPL_WIDTH),
		17210 => to_signed(32664, LUT_AMPL_WIDTH),
		17211 => to_signed(32664, LUT_AMPL_WIDTH),
		17212 => to_signed(32664, LUT_AMPL_WIDTH),
		17213 => to_signed(32664, LUT_AMPL_WIDTH),
		17214 => to_signed(32663, LUT_AMPL_WIDTH),
		17215 => to_signed(32663, LUT_AMPL_WIDTH),
		17216 => to_signed(32663, LUT_AMPL_WIDTH),
		17217 => to_signed(32663, LUT_AMPL_WIDTH),
		17218 => to_signed(32662, LUT_AMPL_WIDTH),
		17219 => to_signed(32662, LUT_AMPL_WIDTH),
		17220 => to_signed(32662, LUT_AMPL_WIDTH),
		17221 => to_signed(32662, LUT_AMPL_WIDTH),
		17222 => to_signed(32661, LUT_AMPL_WIDTH),
		17223 => to_signed(32661, LUT_AMPL_WIDTH),
		17224 => to_signed(32661, LUT_AMPL_WIDTH),
		17225 => to_signed(32661, LUT_AMPL_WIDTH),
		17226 => to_signed(32660, LUT_AMPL_WIDTH),
		17227 => to_signed(32660, LUT_AMPL_WIDTH),
		17228 => to_signed(32660, LUT_AMPL_WIDTH),
		17229 => to_signed(32660, LUT_AMPL_WIDTH),
		17230 => to_signed(32659, LUT_AMPL_WIDTH),
		17231 => to_signed(32659, LUT_AMPL_WIDTH),
		17232 => to_signed(32659, LUT_AMPL_WIDTH),
		17233 => to_signed(32659, LUT_AMPL_WIDTH),
		17234 => to_signed(32658, LUT_AMPL_WIDTH),
		17235 => to_signed(32658, LUT_AMPL_WIDTH),
		17236 => to_signed(32658, LUT_AMPL_WIDTH),
		17237 => to_signed(32657, LUT_AMPL_WIDTH),
		17238 => to_signed(32657, LUT_AMPL_WIDTH),
		17239 => to_signed(32657, LUT_AMPL_WIDTH),
		17240 => to_signed(32657, LUT_AMPL_WIDTH),
		17241 => to_signed(32656, LUT_AMPL_WIDTH),
		17242 => to_signed(32656, LUT_AMPL_WIDTH),
		17243 => to_signed(32656, LUT_AMPL_WIDTH),
		17244 => to_signed(32656, LUT_AMPL_WIDTH),
		17245 => to_signed(32655, LUT_AMPL_WIDTH),
		17246 => to_signed(32655, LUT_AMPL_WIDTH),
		17247 => to_signed(32655, LUT_AMPL_WIDTH),
		17248 => to_signed(32655, LUT_AMPL_WIDTH),
		17249 => to_signed(32654, LUT_AMPL_WIDTH),
		17250 => to_signed(32654, LUT_AMPL_WIDTH),
		17251 => to_signed(32654, LUT_AMPL_WIDTH),
		17252 => to_signed(32654, LUT_AMPL_WIDTH),
		17253 => to_signed(32653, LUT_AMPL_WIDTH),
		17254 => to_signed(32653, LUT_AMPL_WIDTH),
		17255 => to_signed(32653, LUT_AMPL_WIDTH),
		17256 => to_signed(32653, LUT_AMPL_WIDTH),
		17257 => to_signed(32652, LUT_AMPL_WIDTH),
		17258 => to_signed(32652, LUT_AMPL_WIDTH),
		17259 => to_signed(32652, LUT_AMPL_WIDTH),
		17260 => to_signed(32652, LUT_AMPL_WIDTH),
		17261 => to_signed(32651, LUT_AMPL_WIDTH),
		17262 => to_signed(32651, LUT_AMPL_WIDTH),
		17263 => to_signed(32651, LUT_AMPL_WIDTH),
		17264 => to_signed(32650, LUT_AMPL_WIDTH),
		17265 => to_signed(32650, LUT_AMPL_WIDTH),
		17266 => to_signed(32650, LUT_AMPL_WIDTH),
		17267 => to_signed(32650, LUT_AMPL_WIDTH),
		17268 => to_signed(32649, LUT_AMPL_WIDTH),
		17269 => to_signed(32649, LUT_AMPL_WIDTH),
		17270 => to_signed(32649, LUT_AMPL_WIDTH),
		17271 => to_signed(32649, LUT_AMPL_WIDTH),
		17272 => to_signed(32648, LUT_AMPL_WIDTH),
		17273 => to_signed(32648, LUT_AMPL_WIDTH),
		17274 => to_signed(32648, LUT_AMPL_WIDTH),
		17275 => to_signed(32648, LUT_AMPL_WIDTH),
		17276 => to_signed(32647, LUT_AMPL_WIDTH),
		17277 => to_signed(32647, LUT_AMPL_WIDTH),
		17278 => to_signed(32647, LUT_AMPL_WIDTH),
		17279 => to_signed(32646, LUT_AMPL_WIDTH),
		17280 => to_signed(32646, LUT_AMPL_WIDTH),
		17281 => to_signed(32646, LUT_AMPL_WIDTH),
		17282 => to_signed(32646, LUT_AMPL_WIDTH),
		17283 => to_signed(32645, LUT_AMPL_WIDTH),
		17284 => to_signed(32645, LUT_AMPL_WIDTH),
		17285 => to_signed(32645, LUT_AMPL_WIDTH),
		17286 => to_signed(32645, LUT_AMPL_WIDTH),
		17287 => to_signed(32644, LUT_AMPL_WIDTH),
		17288 => to_signed(32644, LUT_AMPL_WIDTH),
		17289 => to_signed(32644, LUT_AMPL_WIDTH),
		17290 => to_signed(32643, LUT_AMPL_WIDTH),
		17291 => to_signed(32643, LUT_AMPL_WIDTH),
		17292 => to_signed(32643, LUT_AMPL_WIDTH),
		17293 => to_signed(32643, LUT_AMPL_WIDTH),
		17294 => to_signed(32642, LUT_AMPL_WIDTH),
		17295 => to_signed(32642, LUT_AMPL_WIDTH),
		17296 => to_signed(32642, LUT_AMPL_WIDTH),
		17297 => to_signed(32642, LUT_AMPL_WIDTH),
		17298 => to_signed(32641, LUT_AMPL_WIDTH),
		17299 => to_signed(32641, LUT_AMPL_WIDTH),
		17300 => to_signed(32641, LUT_AMPL_WIDTH),
		17301 => to_signed(32640, LUT_AMPL_WIDTH),
		17302 => to_signed(32640, LUT_AMPL_WIDTH),
		17303 => to_signed(32640, LUT_AMPL_WIDTH),
		17304 => to_signed(32640, LUT_AMPL_WIDTH),
		17305 => to_signed(32639, LUT_AMPL_WIDTH),
		17306 => to_signed(32639, LUT_AMPL_WIDTH),
		17307 => to_signed(32639, LUT_AMPL_WIDTH),
		17308 => to_signed(32639, LUT_AMPL_WIDTH),
		17309 => to_signed(32638, LUT_AMPL_WIDTH),
		17310 => to_signed(32638, LUT_AMPL_WIDTH),
		17311 => to_signed(32638, LUT_AMPL_WIDTH),
		17312 => to_signed(32637, LUT_AMPL_WIDTH),
		17313 => to_signed(32637, LUT_AMPL_WIDTH),
		17314 => to_signed(32637, LUT_AMPL_WIDTH),
		17315 => to_signed(32637, LUT_AMPL_WIDTH),
		17316 => to_signed(32636, LUT_AMPL_WIDTH),
		17317 => to_signed(32636, LUT_AMPL_WIDTH),
		17318 => to_signed(32636, LUT_AMPL_WIDTH),
		17319 => to_signed(32635, LUT_AMPL_WIDTH),
		17320 => to_signed(32635, LUT_AMPL_WIDTH),
		17321 => to_signed(32635, LUT_AMPL_WIDTH),
		17322 => to_signed(32635, LUT_AMPL_WIDTH),
		17323 => to_signed(32634, LUT_AMPL_WIDTH),
		17324 => to_signed(32634, LUT_AMPL_WIDTH),
		17325 => to_signed(32634, LUT_AMPL_WIDTH),
		17326 => to_signed(32633, LUT_AMPL_WIDTH),
		17327 => to_signed(32633, LUT_AMPL_WIDTH),
		17328 => to_signed(32633, LUT_AMPL_WIDTH),
		17329 => to_signed(32633, LUT_AMPL_WIDTH),
		17330 => to_signed(32632, LUT_AMPL_WIDTH),
		17331 => to_signed(32632, LUT_AMPL_WIDTH),
		17332 => to_signed(32632, LUT_AMPL_WIDTH),
		17333 => to_signed(32631, LUT_AMPL_WIDTH),
		17334 => to_signed(32631, LUT_AMPL_WIDTH),
		17335 => to_signed(32631, LUT_AMPL_WIDTH),
		17336 => to_signed(32631, LUT_AMPL_WIDTH),
		17337 => to_signed(32630, LUT_AMPL_WIDTH),
		17338 => to_signed(32630, LUT_AMPL_WIDTH),
		17339 => to_signed(32630, LUT_AMPL_WIDTH),
		17340 => to_signed(32629, LUT_AMPL_WIDTH),
		17341 => to_signed(32629, LUT_AMPL_WIDTH),
		17342 => to_signed(32629, LUT_AMPL_WIDTH),
		17343 => to_signed(32629, LUT_AMPL_WIDTH),
		17344 => to_signed(32628, LUT_AMPL_WIDTH),
		17345 => to_signed(32628, LUT_AMPL_WIDTH),
		17346 => to_signed(32628, LUT_AMPL_WIDTH),
		17347 => to_signed(32627, LUT_AMPL_WIDTH),
		17348 => to_signed(32627, LUT_AMPL_WIDTH),
		17349 => to_signed(32627, LUT_AMPL_WIDTH),
		17350 => to_signed(32627, LUT_AMPL_WIDTH),
		17351 => to_signed(32626, LUT_AMPL_WIDTH),
		17352 => to_signed(32626, LUT_AMPL_WIDTH),
		17353 => to_signed(32626, LUT_AMPL_WIDTH),
		17354 => to_signed(32625, LUT_AMPL_WIDTH),
		17355 => to_signed(32625, LUT_AMPL_WIDTH),
		17356 => to_signed(32625, LUT_AMPL_WIDTH),
		17357 => to_signed(32625, LUT_AMPL_WIDTH),
		17358 => to_signed(32624, LUT_AMPL_WIDTH),
		17359 => to_signed(32624, LUT_AMPL_WIDTH),
		17360 => to_signed(32624, LUT_AMPL_WIDTH),
		17361 => to_signed(32623, LUT_AMPL_WIDTH),
		17362 => to_signed(32623, LUT_AMPL_WIDTH),
		17363 => to_signed(32623, LUT_AMPL_WIDTH),
		17364 => to_signed(32622, LUT_AMPL_WIDTH),
		17365 => to_signed(32622, LUT_AMPL_WIDTH),
		17366 => to_signed(32622, LUT_AMPL_WIDTH),
		17367 => to_signed(32622, LUT_AMPL_WIDTH),
		17368 => to_signed(32621, LUT_AMPL_WIDTH),
		17369 => to_signed(32621, LUT_AMPL_WIDTH),
		17370 => to_signed(32621, LUT_AMPL_WIDTH),
		17371 => to_signed(32620, LUT_AMPL_WIDTH),
		17372 => to_signed(32620, LUT_AMPL_WIDTH),
		17373 => to_signed(32620, LUT_AMPL_WIDTH),
		17374 => to_signed(32620, LUT_AMPL_WIDTH),
		17375 => to_signed(32619, LUT_AMPL_WIDTH),
		17376 => to_signed(32619, LUT_AMPL_WIDTH),
		17377 => to_signed(32619, LUT_AMPL_WIDTH),
		17378 => to_signed(32618, LUT_AMPL_WIDTH),
		17379 => to_signed(32618, LUT_AMPL_WIDTH),
		17380 => to_signed(32618, LUT_AMPL_WIDTH),
		17381 => to_signed(32617, LUT_AMPL_WIDTH),
		17382 => to_signed(32617, LUT_AMPL_WIDTH),
		17383 => to_signed(32617, LUT_AMPL_WIDTH),
		17384 => to_signed(32617, LUT_AMPL_WIDTH),
		17385 => to_signed(32616, LUT_AMPL_WIDTH),
		17386 => to_signed(32616, LUT_AMPL_WIDTH),
		17387 => to_signed(32616, LUT_AMPL_WIDTH),
		17388 => to_signed(32615, LUT_AMPL_WIDTH),
		17389 => to_signed(32615, LUT_AMPL_WIDTH),
		17390 => to_signed(32615, LUT_AMPL_WIDTH),
		17391 => to_signed(32614, LUT_AMPL_WIDTH),
		17392 => to_signed(32614, LUT_AMPL_WIDTH),
		17393 => to_signed(32614, LUT_AMPL_WIDTH),
		17394 => to_signed(32613, LUT_AMPL_WIDTH),
		17395 => to_signed(32613, LUT_AMPL_WIDTH),
		17396 => to_signed(32613, LUT_AMPL_WIDTH),
		17397 => to_signed(32613, LUT_AMPL_WIDTH),
		17398 => to_signed(32612, LUT_AMPL_WIDTH),
		17399 => to_signed(32612, LUT_AMPL_WIDTH),
		17400 => to_signed(32612, LUT_AMPL_WIDTH),
		17401 => to_signed(32611, LUT_AMPL_WIDTH),
		17402 => to_signed(32611, LUT_AMPL_WIDTH),
		17403 => to_signed(32611, LUT_AMPL_WIDTH),
		17404 => to_signed(32610, LUT_AMPL_WIDTH),
		17405 => to_signed(32610, LUT_AMPL_WIDTH),
		17406 => to_signed(32610, LUT_AMPL_WIDTH),
		17407 => to_signed(32610, LUT_AMPL_WIDTH),
		17408 => to_signed(32609, LUT_AMPL_WIDTH),
		17409 => to_signed(32609, LUT_AMPL_WIDTH),
		17410 => to_signed(32609, LUT_AMPL_WIDTH),
		17411 => to_signed(32608, LUT_AMPL_WIDTH),
		17412 => to_signed(32608, LUT_AMPL_WIDTH),
		17413 => to_signed(32608, LUT_AMPL_WIDTH),
		17414 => to_signed(32607, LUT_AMPL_WIDTH),
		17415 => to_signed(32607, LUT_AMPL_WIDTH),
		17416 => to_signed(32607, LUT_AMPL_WIDTH),
		17417 => to_signed(32606, LUT_AMPL_WIDTH),
		17418 => to_signed(32606, LUT_AMPL_WIDTH),
		17419 => to_signed(32606, LUT_AMPL_WIDTH),
		17420 => to_signed(32606, LUT_AMPL_WIDTH),
		17421 => to_signed(32605, LUT_AMPL_WIDTH),
		17422 => to_signed(32605, LUT_AMPL_WIDTH),
		17423 => to_signed(32605, LUT_AMPL_WIDTH),
		17424 => to_signed(32604, LUT_AMPL_WIDTH),
		17425 => to_signed(32604, LUT_AMPL_WIDTH),
		17426 => to_signed(32604, LUT_AMPL_WIDTH),
		17427 => to_signed(32603, LUT_AMPL_WIDTH),
		17428 => to_signed(32603, LUT_AMPL_WIDTH),
		17429 => to_signed(32603, LUT_AMPL_WIDTH),
		17430 => to_signed(32602, LUT_AMPL_WIDTH),
		17431 => to_signed(32602, LUT_AMPL_WIDTH),
		17432 => to_signed(32602, LUT_AMPL_WIDTH),
		17433 => to_signed(32601, LUT_AMPL_WIDTH),
		17434 => to_signed(32601, LUT_AMPL_WIDTH),
		17435 => to_signed(32601, LUT_AMPL_WIDTH),
		17436 => to_signed(32600, LUT_AMPL_WIDTH),
		17437 => to_signed(32600, LUT_AMPL_WIDTH),
		17438 => to_signed(32600, LUT_AMPL_WIDTH),
		17439 => to_signed(32600, LUT_AMPL_WIDTH),
		17440 => to_signed(32599, LUT_AMPL_WIDTH),
		17441 => to_signed(32599, LUT_AMPL_WIDTH),
		17442 => to_signed(32599, LUT_AMPL_WIDTH),
		17443 => to_signed(32598, LUT_AMPL_WIDTH),
		17444 => to_signed(32598, LUT_AMPL_WIDTH),
		17445 => to_signed(32598, LUT_AMPL_WIDTH),
		17446 => to_signed(32597, LUT_AMPL_WIDTH),
		17447 => to_signed(32597, LUT_AMPL_WIDTH),
		17448 => to_signed(32597, LUT_AMPL_WIDTH),
		17449 => to_signed(32596, LUT_AMPL_WIDTH),
		17450 => to_signed(32596, LUT_AMPL_WIDTH),
		17451 => to_signed(32596, LUT_AMPL_WIDTH),
		17452 => to_signed(32595, LUT_AMPL_WIDTH),
		17453 => to_signed(32595, LUT_AMPL_WIDTH),
		17454 => to_signed(32595, LUT_AMPL_WIDTH),
		17455 => to_signed(32594, LUT_AMPL_WIDTH),
		17456 => to_signed(32594, LUT_AMPL_WIDTH),
		17457 => to_signed(32594, LUT_AMPL_WIDTH),
		17458 => to_signed(32593, LUT_AMPL_WIDTH),
		17459 => to_signed(32593, LUT_AMPL_WIDTH),
		17460 => to_signed(32593, LUT_AMPL_WIDTH),
		17461 => to_signed(32592, LUT_AMPL_WIDTH),
		17462 => to_signed(32592, LUT_AMPL_WIDTH),
		17463 => to_signed(32592, LUT_AMPL_WIDTH),
		17464 => to_signed(32592, LUT_AMPL_WIDTH),
		17465 => to_signed(32591, LUT_AMPL_WIDTH),
		17466 => to_signed(32591, LUT_AMPL_WIDTH),
		17467 => to_signed(32591, LUT_AMPL_WIDTH),
		17468 => to_signed(32590, LUT_AMPL_WIDTH),
		17469 => to_signed(32590, LUT_AMPL_WIDTH),
		17470 => to_signed(32590, LUT_AMPL_WIDTH),
		17471 => to_signed(32589, LUT_AMPL_WIDTH),
		17472 => to_signed(32589, LUT_AMPL_WIDTH),
		17473 => to_signed(32589, LUT_AMPL_WIDTH),
		17474 => to_signed(32588, LUT_AMPL_WIDTH),
		17475 => to_signed(32588, LUT_AMPL_WIDTH),
		17476 => to_signed(32588, LUT_AMPL_WIDTH),
		17477 => to_signed(32587, LUT_AMPL_WIDTH),
		17478 => to_signed(32587, LUT_AMPL_WIDTH),
		17479 => to_signed(32587, LUT_AMPL_WIDTH),
		17480 => to_signed(32586, LUT_AMPL_WIDTH),
		17481 => to_signed(32586, LUT_AMPL_WIDTH),
		17482 => to_signed(32586, LUT_AMPL_WIDTH),
		17483 => to_signed(32585, LUT_AMPL_WIDTH),
		17484 => to_signed(32585, LUT_AMPL_WIDTH),
		17485 => to_signed(32585, LUT_AMPL_WIDTH),
		17486 => to_signed(32584, LUT_AMPL_WIDTH),
		17487 => to_signed(32584, LUT_AMPL_WIDTH),
		17488 => to_signed(32584, LUT_AMPL_WIDTH),
		17489 => to_signed(32583, LUT_AMPL_WIDTH),
		17490 => to_signed(32583, LUT_AMPL_WIDTH),
		17491 => to_signed(32583, LUT_AMPL_WIDTH),
		17492 => to_signed(32582, LUT_AMPL_WIDTH),
		17493 => to_signed(32582, LUT_AMPL_WIDTH),
		17494 => to_signed(32582, LUT_AMPL_WIDTH),
		17495 => to_signed(32581, LUT_AMPL_WIDTH),
		17496 => to_signed(32581, LUT_AMPL_WIDTH),
		17497 => to_signed(32581, LUT_AMPL_WIDTH),
		17498 => to_signed(32580, LUT_AMPL_WIDTH),
		17499 => to_signed(32580, LUT_AMPL_WIDTH),
		17500 => to_signed(32580, LUT_AMPL_WIDTH),
		17501 => to_signed(32579, LUT_AMPL_WIDTH),
		17502 => to_signed(32579, LUT_AMPL_WIDTH),
		17503 => to_signed(32579, LUT_AMPL_WIDTH),
		17504 => to_signed(32578, LUT_AMPL_WIDTH),
		17505 => to_signed(32578, LUT_AMPL_WIDTH),
		17506 => to_signed(32578, LUT_AMPL_WIDTH),
		17507 => to_signed(32577, LUT_AMPL_WIDTH),
		17508 => to_signed(32577, LUT_AMPL_WIDTH),
		17509 => to_signed(32577, LUT_AMPL_WIDTH),
		17510 => to_signed(32576, LUT_AMPL_WIDTH),
		17511 => to_signed(32576, LUT_AMPL_WIDTH),
		17512 => to_signed(32576, LUT_AMPL_WIDTH),
		17513 => to_signed(32575, LUT_AMPL_WIDTH),
		17514 => to_signed(32575, LUT_AMPL_WIDTH),
		17515 => to_signed(32575, LUT_AMPL_WIDTH),
		17516 => to_signed(32574, LUT_AMPL_WIDTH),
		17517 => to_signed(32574, LUT_AMPL_WIDTH),
		17518 => to_signed(32574, LUT_AMPL_WIDTH),
		17519 => to_signed(32573, LUT_AMPL_WIDTH),
		17520 => to_signed(32573, LUT_AMPL_WIDTH),
		17521 => to_signed(32573, LUT_AMPL_WIDTH),
		17522 => to_signed(32572, LUT_AMPL_WIDTH),
		17523 => to_signed(32572, LUT_AMPL_WIDTH),
		17524 => to_signed(32571, LUT_AMPL_WIDTH),
		17525 => to_signed(32571, LUT_AMPL_WIDTH),
		17526 => to_signed(32571, LUT_AMPL_WIDTH),
		17527 => to_signed(32570, LUT_AMPL_WIDTH),
		17528 => to_signed(32570, LUT_AMPL_WIDTH),
		17529 => to_signed(32570, LUT_AMPL_WIDTH),
		17530 => to_signed(32569, LUT_AMPL_WIDTH),
		17531 => to_signed(32569, LUT_AMPL_WIDTH),
		17532 => to_signed(32569, LUT_AMPL_WIDTH),
		17533 => to_signed(32568, LUT_AMPL_WIDTH),
		17534 => to_signed(32568, LUT_AMPL_WIDTH),
		17535 => to_signed(32568, LUT_AMPL_WIDTH),
		17536 => to_signed(32567, LUT_AMPL_WIDTH),
		17537 => to_signed(32567, LUT_AMPL_WIDTH),
		17538 => to_signed(32567, LUT_AMPL_WIDTH),
		17539 => to_signed(32566, LUT_AMPL_WIDTH),
		17540 => to_signed(32566, LUT_AMPL_WIDTH),
		17541 => to_signed(32566, LUT_AMPL_WIDTH),
		17542 => to_signed(32565, LUT_AMPL_WIDTH),
		17543 => to_signed(32565, LUT_AMPL_WIDTH),
		17544 => to_signed(32565, LUT_AMPL_WIDTH),
		17545 => to_signed(32564, LUT_AMPL_WIDTH),
		17546 => to_signed(32564, LUT_AMPL_WIDTH),
		17547 => to_signed(32564, LUT_AMPL_WIDTH),
		17548 => to_signed(32563, LUT_AMPL_WIDTH),
		17549 => to_signed(32563, LUT_AMPL_WIDTH),
		17550 => to_signed(32562, LUT_AMPL_WIDTH),
		17551 => to_signed(32562, LUT_AMPL_WIDTH),
		17552 => to_signed(32562, LUT_AMPL_WIDTH),
		17553 => to_signed(32561, LUT_AMPL_WIDTH),
		17554 => to_signed(32561, LUT_AMPL_WIDTH),
		17555 => to_signed(32561, LUT_AMPL_WIDTH),
		17556 => to_signed(32560, LUT_AMPL_WIDTH),
		17557 => to_signed(32560, LUT_AMPL_WIDTH),
		17558 => to_signed(32560, LUT_AMPL_WIDTH),
		17559 => to_signed(32559, LUT_AMPL_WIDTH),
		17560 => to_signed(32559, LUT_AMPL_WIDTH),
		17561 => to_signed(32559, LUT_AMPL_WIDTH),
		17562 => to_signed(32558, LUT_AMPL_WIDTH),
		17563 => to_signed(32558, LUT_AMPL_WIDTH),
		17564 => to_signed(32558, LUT_AMPL_WIDTH),
		17565 => to_signed(32557, LUT_AMPL_WIDTH),
		17566 => to_signed(32557, LUT_AMPL_WIDTH),
		17567 => to_signed(32556, LUT_AMPL_WIDTH),
		17568 => to_signed(32556, LUT_AMPL_WIDTH),
		17569 => to_signed(32556, LUT_AMPL_WIDTH),
		17570 => to_signed(32555, LUT_AMPL_WIDTH),
		17571 => to_signed(32555, LUT_AMPL_WIDTH),
		17572 => to_signed(32555, LUT_AMPL_WIDTH),
		17573 => to_signed(32554, LUT_AMPL_WIDTH),
		17574 => to_signed(32554, LUT_AMPL_WIDTH),
		17575 => to_signed(32554, LUT_AMPL_WIDTH),
		17576 => to_signed(32553, LUT_AMPL_WIDTH),
		17577 => to_signed(32553, LUT_AMPL_WIDTH),
		17578 => to_signed(32553, LUT_AMPL_WIDTH),
		17579 => to_signed(32552, LUT_AMPL_WIDTH),
		17580 => to_signed(32552, LUT_AMPL_WIDTH),
		17581 => to_signed(32551, LUT_AMPL_WIDTH),
		17582 => to_signed(32551, LUT_AMPL_WIDTH),
		17583 => to_signed(32551, LUT_AMPL_WIDTH),
		17584 => to_signed(32550, LUT_AMPL_WIDTH),
		17585 => to_signed(32550, LUT_AMPL_WIDTH),
		17586 => to_signed(32550, LUT_AMPL_WIDTH),
		17587 => to_signed(32549, LUT_AMPL_WIDTH),
		17588 => to_signed(32549, LUT_AMPL_WIDTH),
		17589 => to_signed(32549, LUT_AMPL_WIDTH),
		17590 => to_signed(32548, LUT_AMPL_WIDTH),
		17591 => to_signed(32548, LUT_AMPL_WIDTH),
		17592 => to_signed(32547, LUT_AMPL_WIDTH),
		17593 => to_signed(32547, LUT_AMPL_WIDTH),
		17594 => to_signed(32547, LUT_AMPL_WIDTH),
		17595 => to_signed(32546, LUT_AMPL_WIDTH),
		17596 => to_signed(32546, LUT_AMPL_WIDTH),
		17597 => to_signed(32546, LUT_AMPL_WIDTH),
		17598 => to_signed(32545, LUT_AMPL_WIDTH),
		17599 => to_signed(32545, LUT_AMPL_WIDTH),
		17600 => to_signed(32545, LUT_AMPL_WIDTH),
		17601 => to_signed(32544, LUT_AMPL_WIDTH),
		17602 => to_signed(32544, LUT_AMPL_WIDTH),
		17603 => to_signed(32543, LUT_AMPL_WIDTH),
		17604 => to_signed(32543, LUT_AMPL_WIDTH),
		17605 => to_signed(32543, LUT_AMPL_WIDTH),
		17606 => to_signed(32542, LUT_AMPL_WIDTH),
		17607 => to_signed(32542, LUT_AMPL_WIDTH),
		17608 => to_signed(32542, LUT_AMPL_WIDTH),
		17609 => to_signed(32541, LUT_AMPL_WIDTH),
		17610 => to_signed(32541, LUT_AMPL_WIDTH),
		17611 => to_signed(32541, LUT_AMPL_WIDTH),
		17612 => to_signed(32540, LUT_AMPL_WIDTH),
		17613 => to_signed(32540, LUT_AMPL_WIDTH),
		17614 => to_signed(32539, LUT_AMPL_WIDTH),
		17615 => to_signed(32539, LUT_AMPL_WIDTH),
		17616 => to_signed(32539, LUT_AMPL_WIDTH),
		17617 => to_signed(32538, LUT_AMPL_WIDTH),
		17618 => to_signed(32538, LUT_AMPL_WIDTH),
		17619 => to_signed(32538, LUT_AMPL_WIDTH),
		17620 => to_signed(32537, LUT_AMPL_WIDTH),
		17621 => to_signed(32537, LUT_AMPL_WIDTH),
		17622 => to_signed(32536, LUT_AMPL_WIDTH),
		17623 => to_signed(32536, LUT_AMPL_WIDTH),
		17624 => to_signed(32536, LUT_AMPL_WIDTH),
		17625 => to_signed(32535, LUT_AMPL_WIDTH),
		17626 => to_signed(32535, LUT_AMPL_WIDTH),
		17627 => to_signed(32535, LUT_AMPL_WIDTH),
		17628 => to_signed(32534, LUT_AMPL_WIDTH),
		17629 => to_signed(32534, LUT_AMPL_WIDTH),
		17630 => to_signed(32533, LUT_AMPL_WIDTH),
		17631 => to_signed(32533, LUT_AMPL_WIDTH),
		17632 => to_signed(32533, LUT_AMPL_WIDTH),
		17633 => to_signed(32532, LUT_AMPL_WIDTH),
		17634 => to_signed(32532, LUT_AMPL_WIDTH),
		17635 => to_signed(32532, LUT_AMPL_WIDTH),
		17636 => to_signed(32531, LUT_AMPL_WIDTH),
		17637 => to_signed(32531, LUT_AMPL_WIDTH),
		17638 => to_signed(32530, LUT_AMPL_WIDTH),
		17639 => to_signed(32530, LUT_AMPL_WIDTH),
		17640 => to_signed(32530, LUT_AMPL_WIDTH),
		17641 => to_signed(32529, LUT_AMPL_WIDTH),
		17642 => to_signed(32529, LUT_AMPL_WIDTH),
		17643 => to_signed(32529, LUT_AMPL_WIDTH),
		17644 => to_signed(32528, LUT_AMPL_WIDTH),
		17645 => to_signed(32528, LUT_AMPL_WIDTH),
		17646 => to_signed(32527, LUT_AMPL_WIDTH),
		17647 => to_signed(32527, LUT_AMPL_WIDTH),
		17648 => to_signed(32527, LUT_AMPL_WIDTH),
		17649 => to_signed(32526, LUT_AMPL_WIDTH),
		17650 => to_signed(32526, LUT_AMPL_WIDTH),
		17651 => to_signed(32526, LUT_AMPL_WIDTH),
		17652 => to_signed(32525, LUT_AMPL_WIDTH),
		17653 => to_signed(32525, LUT_AMPL_WIDTH),
		17654 => to_signed(32524, LUT_AMPL_WIDTH),
		17655 => to_signed(32524, LUT_AMPL_WIDTH),
		17656 => to_signed(32524, LUT_AMPL_WIDTH),
		17657 => to_signed(32523, LUT_AMPL_WIDTH),
		17658 => to_signed(32523, LUT_AMPL_WIDTH),
		17659 => to_signed(32522, LUT_AMPL_WIDTH),
		17660 => to_signed(32522, LUT_AMPL_WIDTH),
		17661 => to_signed(32522, LUT_AMPL_WIDTH),
		17662 => to_signed(32521, LUT_AMPL_WIDTH),
		17663 => to_signed(32521, LUT_AMPL_WIDTH),
		17664 => to_signed(32521, LUT_AMPL_WIDTH),
		17665 => to_signed(32520, LUT_AMPL_WIDTH),
		17666 => to_signed(32520, LUT_AMPL_WIDTH),
		17667 => to_signed(32519, LUT_AMPL_WIDTH),
		17668 => to_signed(32519, LUT_AMPL_WIDTH),
		17669 => to_signed(32519, LUT_AMPL_WIDTH),
		17670 => to_signed(32518, LUT_AMPL_WIDTH),
		17671 => to_signed(32518, LUT_AMPL_WIDTH),
		17672 => to_signed(32517, LUT_AMPL_WIDTH),
		17673 => to_signed(32517, LUT_AMPL_WIDTH),
		17674 => to_signed(32517, LUT_AMPL_WIDTH),
		17675 => to_signed(32516, LUT_AMPL_WIDTH),
		17676 => to_signed(32516, LUT_AMPL_WIDTH),
		17677 => to_signed(32516, LUT_AMPL_WIDTH),
		17678 => to_signed(32515, LUT_AMPL_WIDTH),
		17679 => to_signed(32515, LUT_AMPL_WIDTH),
		17680 => to_signed(32514, LUT_AMPL_WIDTH),
		17681 => to_signed(32514, LUT_AMPL_WIDTH),
		17682 => to_signed(32514, LUT_AMPL_WIDTH),
		17683 => to_signed(32513, LUT_AMPL_WIDTH),
		17684 => to_signed(32513, LUT_AMPL_WIDTH),
		17685 => to_signed(32512, LUT_AMPL_WIDTH),
		17686 => to_signed(32512, LUT_AMPL_WIDTH),
		17687 => to_signed(32512, LUT_AMPL_WIDTH),
		17688 => to_signed(32511, LUT_AMPL_WIDTH),
		17689 => to_signed(32511, LUT_AMPL_WIDTH),
		17690 => to_signed(32510, LUT_AMPL_WIDTH),
		17691 => to_signed(32510, LUT_AMPL_WIDTH),
		17692 => to_signed(32510, LUT_AMPL_WIDTH),
		17693 => to_signed(32509, LUT_AMPL_WIDTH),
		17694 => to_signed(32509, LUT_AMPL_WIDTH),
		17695 => to_signed(32509, LUT_AMPL_WIDTH),
		17696 => to_signed(32508, LUT_AMPL_WIDTH),
		17697 => to_signed(32508, LUT_AMPL_WIDTH),
		17698 => to_signed(32507, LUT_AMPL_WIDTH),
		17699 => to_signed(32507, LUT_AMPL_WIDTH),
		17700 => to_signed(32507, LUT_AMPL_WIDTH),
		17701 => to_signed(32506, LUT_AMPL_WIDTH),
		17702 => to_signed(32506, LUT_AMPL_WIDTH),
		17703 => to_signed(32505, LUT_AMPL_WIDTH),
		17704 => to_signed(32505, LUT_AMPL_WIDTH),
		17705 => to_signed(32505, LUT_AMPL_WIDTH),
		17706 => to_signed(32504, LUT_AMPL_WIDTH),
		17707 => to_signed(32504, LUT_AMPL_WIDTH),
		17708 => to_signed(32503, LUT_AMPL_WIDTH),
		17709 => to_signed(32503, LUT_AMPL_WIDTH),
		17710 => to_signed(32503, LUT_AMPL_WIDTH),
		17711 => to_signed(32502, LUT_AMPL_WIDTH),
		17712 => to_signed(32502, LUT_AMPL_WIDTH),
		17713 => to_signed(32501, LUT_AMPL_WIDTH),
		17714 => to_signed(32501, LUT_AMPL_WIDTH),
		17715 => to_signed(32501, LUT_AMPL_WIDTH),
		17716 => to_signed(32500, LUT_AMPL_WIDTH),
		17717 => to_signed(32500, LUT_AMPL_WIDTH),
		17718 => to_signed(32499, LUT_AMPL_WIDTH),
		17719 => to_signed(32499, LUT_AMPL_WIDTH),
		17720 => to_signed(32499, LUT_AMPL_WIDTH),
		17721 => to_signed(32498, LUT_AMPL_WIDTH),
		17722 => to_signed(32498, LUT_AMPL_WIDTH),
		17723 => to_signed(32497, LUT_AMPL_WIDTH),
		17724 => to_signed(32497, LUT_AMPL_WIDTH),
		17725 => to_signed(32497, LUT_AMPL_WIDTH),
		17726 => to_signed(32496, LUT_AMPL_WIDTH),
		17727 => to_signed(32496, LUT_AMPL_WIDTH),
		17728 => to_signed(32495, LUT_AMPL_WIDTH),
		17729 => to_signed(32495, LUT_AMPL_WIDTH),
		17730 => to_signed(32495, LUT_AMPL_WIDTH),
		17731 => to_signed(32494, LUT_AMPL_WIDTH),
		17732 => to_signed(32494, LUT_AMPL_WIDTH),
		17733 => to_signed(32493, LUT_AMPL_WIDTH),
		17734 => to_signed(32493, LUT_AMPL_WIDTH),
		17735 => to_signed(32493, LUT_AMPL_WIDTH),
		17736 => to_signed(32492, LUT_AMPL_WIDTH),
		17737 => to_signed(32492, LUT_AMPL_WIDTH),
		17738 => to_signed(32491, LUT_AMPL_WIDTH),
		17739 => to_signed(32491, LUT_AMPL_WIDTH),
		17740 => to_signed(32490, LUT_AMPL_WIDTH),
		17741 => to_signed(32490, LUT_AMPL_WIDTH),
		17742 => to_signed(32490, LUT_AMPL_WIDTH),
		17743 => to_signed(32489, LUT_AMPL_WIDTH),
		17744 => to_signed(32489, LUT_AMPL_WIDTH),
		17745 => to_signed(32488, LUT_AMPL_WIDTH),
		17746 => to_signed(32488, LUT_AMPL_WIDTH),
		17747 => to_signed(32488, LUT_AMPL_WIDTH),
		17748 => to_signed(32487, LUT_AMPL_WIDTH),
		17749 => to_signed(32487, LUT_AMPL_WIDTH),
		17750 => to_signed(32486, LUT_AMPL_WIDTH),
		17751 => to_signed(32486, LUT_AMPL_WIDTH),
		17752 => to_signed(32486, LUT_AMPL_WIDTH),
		17753 => to_signed(32485, LUT_AMPL_WIDTH),
		17754 => to_signed(32485, LUT_AMPL_WIDTH),
		17755 => to_signed(32484, LUT_AMPL_WIDTH),
		17756 => to_signed(32484, LUT_AMPL_WIDTH),
		17757 => to_signed(32484, LUT_AMPL_WIDTH),
		17758 => to_signed(32483, LUT_AMPL_WIDTH),
		17759 => to_signed(32483, LUT_AMPL_WIDTH),
		17760 => to_signed(32482, LUT_AMPL_WIDTH),
		17761 => to_signed(32482, LUT_AMPL_WIDTH),
		17762 => to_signed(32481, LUT_AMPL_WIDTH),
		17763 => to_signed(32481, LUT_AMPL_WIDTH),
		17764 => to_signed(32481, LUT_AMPL_WIDTH),
		17765 => to_signed(32480, LUT_AMPL_WIDTH),
		17766 => to_signed(32480, LUT_AMPL_WIDTH),
		17767 => to_signed(32479, LUT_AMPL_WIDTH),
		17768 => to_signed(32479, LUT_AMPL_WIDTH),
		17769 => to_signed(32479, LUT_AMPL_WIDTH),
		17770 => to_signed(32478, LUT_AMPL_WIDTH),
		17771 => to_signed(32478, LUT_AMPL_WIDTH),
		17772 => to_signed(32477, LUT_AMPL_WIDTH),
		17773 => to_signed(32477, LUT_AMPL_WIDTH),
		17774 => to_signed(32476, LUT_AMPL_WIDTH),
		17775 => to_signed(32476, LUT_AMPL_WIDTH),
		17776 => to_signed(32476, LUT_AMPL_WIDTH),
		17777 => to_signed(32475, LUT_AMPL_WIDTH),
		17778 => to_signed(32475, LUT_AMPL_WIDTH),
		17779 => to_signed(32474, LUT_AMPL_WIDTH),
		17780 => to_signed(32474, LUT_AMPL_WIDTH),
		17781 => to_signed(32474, LUT_AMPL_WIDTH),
		17782 => to_signed(32473, LUT_AMPL_WIDTH),
		17783 => to_signed(32473, LUT_AMPL_WIDTH),
		17784 => to_signed(32472, LUT_AMPL_WIDTH),
		17785 => to_signed(32472, LUT_AMPL_WIDTH),
		17786 => to_signed(32471, LUT_AMPL_WIDTH),
		17787 => to_signed(32471, LUT_AMPL_WIDTH),
		17788 => to_signed(32471, LUT_AMPL_WIDTH),
		17789 => to_signed(32470, LUT_AMPL_WIDTH),
		17790 => to_signed(32470, LUT_AMPL_WIDTH),
		17791 => to_signed(32469, LUT_AMPL_WIDTH),
		17792 => to_signed(32469, LUT_AMPL_WIDTH),
		17793 => to_signed(32468, LUT_AMPL_WIDTH),
		17794 => to_signed(32468, LUT_AMPL_WIDTH),
		17795 => to_signed(32468, LUT_AMPL_WIDTH),
		17796 => to_signed(32467, LUT_AMPL_WIDTH),
		17797 => to_signed(32467, LUT_AMPL_WIDTH),
		17798 => to_signed(32466, LUT_AMPL_WIDTH),
		17799 => to_signed(32466, LUT_AMPL_WIDTH),
		17800 => to_signed(32466, LUT_AMPL_WIDTH),
		17801 => to_signed(32465, LUT_AMPL_WIDTH),
		17802 => to_signed(32465, LUT_AMPL_WIDTH),
		17803 => to_signed(32464, LUT_AMPL_WIDTH),
		17804 => to_signed(32464, LUT_AMPL_WIDTH),
		17805 => to_signed(32463, LUT_AMPL_WIDTH),
		17806 => to_signed(32463, LUT_AMPL_WIDTH),
		17807 => to_signed(32463, LUT_AMPL_WIDTH),
		17808 => to_signed(32462, LUT_AMPL_WIDTH),
		17809 => to_signed(32462, LUT_AMPL_WIDTH),
		17810 => to_signed(32461, LUT_AMPL_WIDTH),
		17811 => to_signed(32461, LUT_AMPL_WIDTH),
		17812 => to_signed(32460, LUT_AMPL_WIDTH),
		17813 => to_signed(32460, LUT_AMPL_WIDTH),
		17814 => to_signed(32460, LUT_AMPL_WIDTH),
		17815 => to_signed(32459, LUT_AMPL_WIDTH),
		17816 => to_signed(32459, LUT_AMPL_WIDTH),
		17817 => to_signed(32458, LUT_AMPL_WIDTH),
		17818 => to_signed(32458, LUT_AMPL_WIDTH),
		17819 => to_signed(32457, LUT_AMPL_WIDTH),
		17820 => to_signed(32457, LUT_AMPL_WIDTH),
		17821 => to_signed(32457, LUT_AMPL_WIDTH),
		17822 => to_signed(32456, LUT_AMPL_WIDTH),
		17823 => to_signed(32456, LUT_AMPL_WIDTH),
		17824 => to_signed(32455, LUT_AMPL_WIDTH),
		17825 => to_signed(32455, LUT_AMPL_WIDTH),
		17826 => to_signed(32454, LUT_AMPL_WIDTH),
		17827 => to_signed(32454, LUT_AMPL_WIDTH),
		17828 => to_signed(32453, LUT_AMPL_WIDTH),
		17829 => to_signed(32453, LUT_AMPL_WIDTH),
		17830 => to_signed(32453, LUT_AMPL_WIDTH),
		17831 => to_signed(32452, LUT_AMPL_WIDTH),
		17832 => to_signed(32452, LUT_AMPL_WIDTH),
		17833 => to_signed(32451, LUT_AMPL_WIDTH),
		17834 => to_signed(32451, LUT_AMPL_WIDTH),
		17835 => to_signed(32450, LUT_AMPL_WIDTH),
		17836 => to_signed(32450, LUT_AMPL_WIDTH),
		17837 => to_signed(32450, LUT_AMPL_WIDTH),
		17838 => to_signed(32449, LUT_AMPL_WIDTH),
		17839 => to_signed(32449, LUT_AMPL_WIDTH),
		17840 => to_signed(32448, LUT_AMPL_WIDTH),
		17841 => to_signed(32448, LUT_AMPL_WIDTH),
		17842 => to_signed(32447, LUT_AMPL_WIDTH),
		17843 => to_signed(32447, LUT_AMPL_WIDTH),
		17844 => to_signed(32447, LUT_AMPL_WIDTH),
		17845 => to_signed(32446, LUT_AMPL_WIDTH),
		17846 => to_signed(32446, LUT_AMPL_WIDTH),
		17847 => to_signed(32445, LUT_AMPL_WIDTH),
		17848 => to_signed(32445, LUT_AMPL_WIDTH),
		17849 => to_signed(32444, LUT_AMPL_WIDTH),
		17850 => to_signed(32444, LUT_AMPL_WIDTH),
		17851 => to_signed(32443, LUT_AMPL_WIDTH),
		17852 => to_signed(32443, LUT_AMPL_WIDTH),
		17853 => to_signed(32443, LUT_AMPL_WIDTH),
		17854 => to_signed(32442, LUT_AMPL_WIDTH),
		17855 => to_signed(32442, LUT_AMPL_WIDTH),
		17856 => to_signed(32441, LUT_AMPL_WIDTH),
		17857 => to_signed(32441, LUT_AMPL_WIDTH),
		17858 => to_signed(32440, LUT_AMPL_WIDTH),
		17859 => to_signed(32440, LUT_AMPL_WIDTH),
		17860 => to_signed(32439, LUT_AMPL_WIDTH),
		17861 => to_signed(32439, LUT_AMPL_WIDTH),
		17862 => to_signed(32439, LUT_AMPL_WIDTH),
		17863 => to_signed(32438, LUT_AMPL_WIDTH),
		17864 => to_signed(32438, LUT_AMPL_WIDTH),
		17865 => to_signed(32437, LUT_AMPL_WIDTH),
		17866 => to_signed(32437, LUT_AMPL_WIDTH),
		17867 => to_signed(32436, LUT_AMPL_WIDTH),
		17868 => to_signed(32436, LUT_AMPL_WIDTH),
		17869 => to_signed(32435, LUT_AMPL_WIDTH),
		17870 => to_signed(32435, LUT_AMPL_WIDTH),
		17871 => to_signed(32435, LUT_AMPL_WIDTH),
		17872 => to_signed(32434, LUT_AMPL_WIDTH),
		17873 => to_signed(32434, LUT_AMPL_WIDTH),
		17874 => to_signed(32433, LUT_AMPL_WIDTH),
		17875 => to_signed(32433, LUT_AMPL_WIDTH),
		17876 => to_signed(32432, LUT_AMPL_WIDTH),
		17877 => to_signed(32432, LUT_AMPL_WIDTH),
		17878 => to_signed(32431, LUT_AMPL_WIDTH),
		17879 => to_signed(32431, LUT_AMPL_WIDTH),
		17880 => to_signed(32431, LUT_AMPL_WIDTH),
		17881 => to_signed(32430, LUT_AMPL_WIDTH),
		17882 => to_signed(32430, LUT_AMPL_WIDTH),
		17883 => to_signed(32429, LUT_AMPL_WIDTH),
		17884 => to_signed(32429, LUT_AMPL_WIDTH),
		17885 => to_signed(32428, LUT_AMPL_WIDTH),
		17886 => to_signed(32428, LUT_AMPL_WIDTH),
		17887 => to_signed(32427, LUT_AMPL_WIDTH),
		17888 => to_signed(32427, LUT_AMPL_WIDTH),
		17889 => to_signed(32426, LUT_AMPL_WIDTH),
		17890 => to_signed(32426, LUT_AMPL_WIDTH),
		17891 => to_signed(32426, LUT_AMPL_WIDTH),
		17892 => to_signed(32425, LUT_AMPL_WIDTH),
		17893 => to_signed(32425, LUT_AMPL_WIDTH),
		17894 => to_signed(32424, LUT_AMPL_WIDTH),
		17895 => to_signed(32424, LUT_AMPL_WIDTH),
		17896 => to_signed(32423, LUT_AMPL_WIDTH),
		17897 => to_signed(32423, LUT_AMPL_WIDTH),
		17898 => to_signed(32422, LUT_AMPL_WIDTH),
		17899 => to_signed(32422, LUT_AMPL_WIDTH),
		17900 => to_signed(32422, LUT_AMPL_WIDTH),
		17901 => to_signed(32421, LUT_AMPL_WIDTH),
		17902 => to_signed(32421, LUT_AMPL_WIDTH),
		17903 => to_signed(32420, LUT_AMPL_WIDTH),
		17904 => to_signed(32420, LUT_AMPL_WIDTH),
		17905 => to_signed(32419, LUT_AMPL_WIDTH),
		17906 => to_signed(32419, LUT_AMPL_WIDTH),
		17907 => to_signed(32418, LUT_AMPL_WIDTH),
		17908 => to_signed(32418, LUT_AMPL_WIDTH),
		17909 => to_signed(32417, LUT_AMPL_WIDTH),
		17910 => to_signed(32417, LUT_AMPL_WIDTH),
		17911 => to_signed(32416, LUT_AMPL_WIDTH),
		17912 => to_signed(32416, LUT_AMPL_WIDTH),
		17913 => to_signed(32416, LUT_AMPL_WIDTH),
		17914 => to_signed(32415, LUT_AMPL_WIDTH),
		17915 => to_signed(32415, LUT_AMPL_WIDTH),
		17916 => to_signed(32414, LUT_AMPL_WIDTH),
		17917 => to_signed(32414, LUT_AMPL_WIDTH),
		17918 => to_signed(32413, LUT_AMPL_WIDTH),
		17919 => to_signed(32413, LUT_AMPL_WIDTH),
		17920 => to_signed(32412, LUT_AMPL_WIDTH),
		17921 => to_signed(32412, LUT_AMPL_WIDTH),
		17922 => to_signed(32411, LUT_AMPL_WIDTH),
		17923 => to_signed(32411, LUT_AMPL_WIDTH),
		17924 => to_signed(32411, LUT_AMPL_WIDTH),
		17925 => to_signed(32410, LUT_AMPL_WIDTH),
		17926 => to_signed(32410, LUT_AMPL_WIDTH),
		17927 => to_signed(32409, LUT_AMPL_WIDTH),
		17928 => to_signed(32409, LUT_AMPL_WIDTH),
		17929 => to_signed(32408, LUT_AMPL_WIDTH),
		17930 => to_signed(32408, LUT_AMPL_WIDTH),
		17931 => to_signed(32407, LUT_AMPL_WIDTH),
		17932 => to_signed(32407, LUT_AMPL_WIDTH),
		17933 => to_signed(32406, LUT_AMPL_WIDTH),
		17934 => to_signed(32406, LUT_AMPL_WIDTH),
		17935 => to_signed(32405, LUT_AMPL_WIDTH),
		17936 => to_signed(32405, LUT_AMPL_WIDTH),
		17937 => to_signed(32404, LUT_AMPL_WIDTH),
		17938 => to_signed(32404, LUT_AMPL_WIDTH),
		17939 => to_signed(32404, LUT_AMPL_WIDTH),
		17940 => to_signed(32403, LUT_AMPL_WIDTH),
		17941 => to_signed(32403, LUT_AMPL_WIDTH),
		17942 => to_signed(32402, LUT_AMPL_WIDTH),
		17943 => to_signed(32402, LUT_AMPL_WIDTH),
		17944 => to_signed(32401, LUT_AMPL_WIDTH),
		17945 => to_signed(32401, LUT_AMPL_WIDTH),
		17946 => to_signed(32400, LUT_AMPL_WIDTH),
		17947 => to_signed(32400, LUT_AMPL_WIDTH),
		17948 => to_signed(32399, LUT_AMPL_WIDTH),
		17949 => to_signed(32399, LUT_AMPL_WIDTH),
		17950 => to_signed(32398, LUT_AMPL_WIDTH),
		17951 => to_signed(32398, LUT_AMPL_WIDTH),
		17952 => to_signed(32397, LUT_AMPL_WIDTH),
		17953 => to_signed(32397, LUT_AMPL_WIDTH),
		17954 => to_signed(32397, LUT_AMPL_WIDTH),
		17955 => to_signed(32396, LUT_AMPL_WIDTH),
		17956 => to_signed(32396, LUT_AMPL_WIDTH),
		17957 => to_signed(32395, LUT_AMPL_WIDTH),
		17958 => to_signed(32395, LUT_AMPL_WIDTH),
		17959 => to_signed(32394, LUT_AMPL_WIDTH),
		17960 => to_signed(32394, LUT_AMPL_WIDTH),
		17961 => to_signed(32393, LUT_AMPL_WIDTH),
		17962 => to_signed(32393, LUT_AMPL_WIDTH),
		17963 => to_signed(32392, LUT_AMPL_WIDTH),
		17964 => to_signed(32392, LUT_AMPL_WIDTH),
		17965 => to_signed(32391, LUT_AMPL_WIDTH),
		17966 => to_signed(32391, LUT_AMPL_WIDTH),
		17967 => to_signed(32390, LUT_AMPL_WIDTH),
		17968 => to_signed(32390, LUT_AMPL_WIDTH),
		17969 => to_signed(32389, LUT_AMPL_WIDTH),
		17970 => to_signed(32389, LUT_AMPL_WIDTH),
		17971 => to_signed(32388, LUT_AMPL_WIDTH),
		17972 => to_signed(32388, LUT_AMPL_WIDTH),
		17973 => to_signed(32387, LUT_AMPL_WIDTH),
		17974 => to_signed(32387, LUT_AMPL_WIDTH),
		17975 => to_signed(32387, LUT_AMPL_WIDTH),
		17976 => to_signed(32386, LUT_AMPL_WIDTH),
		17977 => to_signed(32386, LUT_AMPL_WIDTH),
		17978 => to_signed(32385, LUT_AMPL_WIDTH),
		17979 => to_signed(32385, LUT_AMPL_WIDTH),
		17980 => to_signed(32384, LUT_AMPL_WIDTH),
		17981 => to_signed(32384, LUT_AMPL_WIDTH),
		17982 => to_signed(32383, LUT_AMPL_WIDTH),
		17983 => to_signed(32383, LUT_AMPL_WIDTH),
		17984 => to_signed(32382, LUT_AMPL_WIDTH),
		17985 => to_signed(32382, LUT_AMPL_WIDTH),
		17986 => to_signed(32381, LUT_AMPL_WIDTH),
		17987 => to_signed(32381, LUT_AMPL_WIDTH),
		17988 => to_signed(32380, LUT_AMPL_WIDTH),
		17989 => to_signed(32380, LUT_AMPL_WIDTH),
		17990 => to_signed(32379, LUT_AMPL_WIDTH),
		17991 => to_signed(32379, LUT_AMPL_WIDTH),
		17992 => to_signed(32378, LUT_AMPL_WIDTH),
		17993 => to_signed(32378, LUT_AMPL_WIDTH),
		17994 => to_signed(32377, LUT_AMPL_WIDTH),
		17995 => to_signed(32377, LUT_AMPL_WIDTH),
		17996 => to_signed(32376, LUT_AMPL_WIDTH),
		17997 => to_signed(32376, LUT_AMPL_WIDTH),
		17998 => to_signed(32375, LUT_AMPL_WIDTH),
		17999 => to_signed(32375, LUT_AMPL_WIDTH),
		18000 => to_signed(32375, LUT_AMPL_WIDTH),
		18001 => to_signed(32374, LUT_AMPL_WIDTH),
		18002 => to_signed(32374, LUT_AMPL_WIDTH),
		18003 => to_signed(32373, LUT_AMPL_WIDTH),
		18004 => to_signed(32373, LUT_AMPL_WIDTH),
		18005 => to_signed(32372, LUT_AMPL_WIDTH),
		18006 => to_signed(32372, LUT_AMPL_WIDTH),
		18007 => to_signed(32371, LUT_AMPL_WIDTH),
		18008 => to_signed(32371, LUT_AMPL_WIDTH),
		18009 => to_signed(32370, LUT_AMPL_WIDTH),
		18010 => to_signed(32370, LUT_AMPL_WIDTH),
		18011 => to_signed(32369, LUT_AMPL_WIDTH),
		18012 => to_signed(32369, LUT_AMPL_WIDTH),
		18013 => to_signed(32368, LUT_AMPL_WIDTH),
		18014 => to_signed(32368, LUT_AMPL_WIDTH),
		18015 => to_signed(32367, LUT_AMPL_WIDTH),
		18016 => to_signed(32367, LUT_AMPL_WIDTH),
		18017 => to_signed(32366, LUT_AMPL_WIDTH),
		18018 => to_signed(32366, LUT_AMPL_WIDTH),
		18019 => to_signed(32365, LUT_AMPL_WIDTH),
		18020 => to_signed(32365, LUT_AMPL_WIDTH),
		18021 => to_signed(32364, LUT_AMPL_WIDTH),
		18022 => to_signed(32364, LUT_AMPL_WIDTH),
		18023 => to_signed(32363, LUT_AMPL_WIDTH),
		18024 => to_signed(32363, LUT_AMPL_WIDTH),
		18025 => to_signed(32362, LUT_AMPL_WIDTH),
		18026 => to_signed(32362, LUT_AMPL_WIDTH),
		18027 => to_signed(32361, LUT_AMPL_WIDTH),
		18028 => to_signed(32361, LUT_AMPL_WIDTH),
		18029 => to_signed(32360, LUT_AMPL_WIDTH),
		18030 => to_signed(32360, LUT_AMPL_WIDTH),
		18031 => to_signed(32359, LUT_AMPL_WIDTH),
		18032 => to_signed(32359, LUT_AMPL_WIDTH),
		18033 => to_signed(32358, LUT_AMPL_WIDTH),
		18034 => to_signed(32358, LUT_AMPL_WIDTH),
		18035 => to_signed(32357, LUT_AMPL_WIDTH),
		18036 => to_signed(32357, LUT_AMPL_WIDTH),
		18037 => to_signed(32356, LUT_AMPL_WIDTH),
		18038 => to_signed(32356, LUT_AMPL_WIDTH),
		18039 => to_signed(32355, LUT_AMPL_WIDTH),
		18040 => to_signed(32355, LUT_AMPL_WIDTH),
		18041 => to_signed(32354, LUT_AMPL_WIDTH),
		18042 => to_signed(32354, LUT_AMPL_WIDTH),
		18043 => to_signed(32353, LUT_AMPL_WIDTH),
		18044 => to_signed(32353, LUT_AMPL_WIDTH),
		18045 => to_signed(32352, LUT_AMPL_WIDTH),
		18046 => to_signed(32352, LUT_AMPL_WIDTH),
		18047 => to_signed(32351, LUT_AMPL_WIDTH),
		18048 => to_signed(32351, LUT_AMPL_WIDTH),
		18049 => to_signed(32350, LUT_AMPL_WIDTH),
		18050 => to_signed(32350, LUT_AMPL_WIDTH),
		18051 => to_signed(32349, LUT_AMPL_WIDTH),
		18052 => to_signed(32349, LUT_AMPL_WIDTH),
		18053 => to_signed(32348, LUT_AMPL_WIDTH),
		18054 => to_signed(32348, LUT_AMPL_WIDTH),
		18055 => to_signed(32347, LUT_AMPL_WIDTH),
		18056 => to_signed(32347, LUT_AMPL_WIDTH),
		18057 => to_signed(32346, LUT_AMPL_WIDTH),
		18058 => to_signed(32346, LUT_AMPL_WIDTH),
		18059 => to_signed(32345, LUT_AMPL_WIDTH),
		18060 => to_signed(32345, LUT_AMPL_WIDTH),
		18061 => to_signed(32344, LUT_AMPL_WIDTH),
		18062 => to_signed(32344, LUT_AMPL_WIDTH),
		18063 => to_signed(32343, LUT_AMPL_WIDTH),
		18064 => to_signed(32343, LUT_AMPL_WIDTH),
		18065 => to_signed(32342, LUT_AMPL_WIDTH),
		18066 => to_signed(32342, LUT_AMPL_WIDTH),
		18067 => to_signed(32341, LUT_AMPL_WIDTH),
		18068 => to_signed(32341, LUT_AMPL_WIDTH),
		18069 => to_signed(32340, LUT_AMPL_WIDTH),
		18070 => to_signed(32340, LUT_AMPL_WIDTH),
		18071 => to_signed(32339, LUT_AMPL_WIDTH),
		18072 => to_signed(32339, LUT_AMPL_WIDTH),
		18073 => to_signed(32338, LUT_AMPL_WIDTH),
		18074 => to_signed(32338, LUT_AMPL_WIDTH),
		18075 => to_signed(32337, LUT_AMPL_WIDTH),
		18076 => to_signed(32337, LUT_AMPL_WIDTH),
		18077 => to_signed(32336, LUT_AMPL_WIDTH),
		18078 => to_signed(32336, LUT_AMPL_WIDTH),
		18079 => to_signed(32335, LUT_AMPL_WIDTH),
		18080 => to_signed(32335, LUT_AMPL_WIDTH),
		18081 => to_signed(32334, LUT_AMPL_WIDTH),
		18082 => to_signed(32334, LUT_AMPL_WIDTH),
		18083 => to_signed(32333, LUT_AMPL_WIDTH),
		18084 => to_signed(32333, LUT_AMPL_WIDTH),
		18085 => to_signed(32332, LUT_AMPL_WIDTH),
		18086 => to_signed(32332, LUT_AMPL_WIDTH),
		18087 => to_signed(32331, LUT_AMPL_WIDTH),
		18088 => to_signed(32331, LUT_AMPL_WIDTH),
		18089 => to_signed(32330, LUT_AMPL_WIDTH),
		18090 => to_signed(32330, LUT_AMPL_WIDTH),
		18091 => to_signed(32329, LUT_AMPL_WIDTH),
		18092 => to_signed(32329, LUT_AMPL_WIDTH),
		18093 => to_signed(32328, LUT_AMPL_WIDTH),
		18094 => to_signed(32328, LUT_AMPL_WIDTH),
		18095 => to_signed(32327, LUT_AMPL_WIDTH),
		18096 => to_signed(32327, LUT_AMPL_WIDTH),
		18097 => to_signed(32326, LUT_AMPL_WIDTH),
		18098 => to_signed(32326, LUT_AMPL_WIDTH),
		18099 => to_signed(32325, LUT_AMPL_WIDTH),
		18100 => to_signed(32325, LUT_AMPL_WIDTH),
		18101 => to_signed(32324, LUT_AMPL_WIDTH),
		18102 => to_signed(32324, LUT_AMPL_WIDTH),
		18103 => to_signed(32323, LUT_AMPL_WIDTH),
		18104 => to_signed(32322, LUT_AMPL_WIDTH),
		18105 => to_signed(32322, LUT_AMPL_WIDTH),
		18106 => to_signed(32321, LUT_AMPL_WIDTH),
		18107 => to_signed(32321, LUT_AMPL_WIDTH),
		18108 => to_signed(32320, LUT_AMPL_WIDTH),
		18109 => to_signed(32320, LUT_AMPL_WIDTH),
		18110 => to_signed(32319, LUT_AMPL_WIDTH),
		18111 => to_signed(32319, LUT_AMPL_WIDTH),
		18112 => to_signed(32318, LUT_AMPL_WIDTH),
		18113 => to_signed(32318, LUT_AMPL_WIDTH),
		18114 => to_signed(32317, LUT_AMPL_WIDTH),
		18115 => to_signed(32317, LUT_AMPL_WIDTH),
		18116 => to_signed(32316, LUT_AMPL_WIDTH),
		18117 => to_signed(32316, LUT_AMPL_WIDTH),
		18118 => to_signed(32315, LUT_AMPL_WIDTH),
		18119 => to_signed(32315, LUT_AMPL_WIDTH),
		18120 => to_signed(32314, LUT_AMPL_WIDTH),
		18121 => to_signed(32314, LUT_AMPL_WIDTH),
		18122 => to_signed(32313, LUT_AMPL_WIDTH),
		18123 => to_signed(32313, LUT_AMPL_WIDTH),
		18124 => to_signed(32312, LUT_AMPL_WIDTH),
		18125 => to_signed(32312, LUT_AMPL_WIDTH),
		18126 => to_signed(32311, LUT_AMPL_WIDTH),
		18127 => to_signed(32311, LUT_AMPL_WIDTH),
		18128 => to_signed(32310, LUT_AMPL_WIDTH),
		18129 => to_signed(32310, LUT_AMPL_WIDTH),
		18130 => to_signed(32309, LUT_AMPL_WIDTH),
		18131 => to_signed(32308, LUT_AMPL_WIDTH),
		18132 => to_signed(32308, LUT_AMPL_WIDTH),
		18133 => to_signed(32307, LUT_AMPL_WIDTH),
		18134 => to_signed(32307, LUT_AMPL_WIDTH),
		18135 => to_signed(32306, LUT_AMPL_WIDTH),
		18136 => to_signed(32306, LUT_AMPL_WIDTH),
		18137 => to_signed(32305, LUT_AMPL_WIDTH),
		18138 => to_signed(32305, LUT_AMPL_WIDTH),
		18139 => to_signed(32304, LUT_AMPL_WIDTH),
		18140 => to_signed(32304, LUT_AMPL_WIDTH),
		18141 => to_signed(32303, LUT_AMPL_WIDTH),
		18142 => to_signed(32303, LUT_AMPL_WIDTH),
		18143 => to_signed(32302, LUT_AMPL_WIDTH),
		18144 => to_signed(32302, LUT_AMPL_WIDTH),
		18145 => to_signed(32301, LUT_AMPL_WIDTH),
		18146 => to_signed(32301, LUT_AMPL_WIDTH),
		18147 => to_signed(32300, LUT_AMPL_WIDTH),
		18148 => to_signed(32300, LUT_AMPL_WIDTH),
		18149 => to_signed(32299, LUT_AMPL_WIDTH),
		18150 => to_signed(32298, LUT_AMPL_WIDTH),
		18151 => to_signed(32298, LUT_AMPL_WIDTH),
		18152 => to_signed(32297, LUT_AMPL_WIDTH),
		18153 => to_signed(32297, LUT_AMPL_WIDTH),
		18154 => to_signed(32296, LUT_AMPL_WIDTH),
		18155 => to_signed(32296, LUT_AMPL_WIDTH),
		18156 => to_signed(32295, LUT_AMPL_WIDTH),
		18157 => to_signed(32295, LUT_AMPL_WIDTH),
		18158 => to_signed(32294, LUT_AMPL_WIDTH),
		18159 => to_signed(32294, LUT_AMPL_WIDTH),
		18160 => to_signed(32293, LUT_AMPL_WIDTH),
		18161 => to_signed(32293, LUT_AMPL_WIDTH),
		18162 => to_signed(32292, LUT_AMPL_WIDTH),
		18163 => to_signed(32292, LUT_AMPL_WIDTH),
		18164 => to_signed(32291, LUT_AMPL_WIDTH),
		18165 => to_signed(32290, LUT_AMPL_WIDTH),
		18166 => to_signed(32290, LUT_AMPL_WIDTH),
		18167 => to_signed(32289, LUT_AMPL_WIDTH),
		18168 => to_signed(32289, LUT_AMPL_WIDTH),
		18169 => to_signed(32288, LUT_AMPL_WIDTH),
		18170 => to_signed(32288, LUT_AMPL_WIDTH),
		18171 => to_signed(32287, LUT_AMPL_WIDTH),
		18172 => to_signed(32287, LUT_AMPL_WIDTH),
		18173 => to_signed(32286, LUT_AMPL_WIDTH),
		18174 => to_signed(32286, LUT_AMPL_WIDTH),
		18175 => to_signed(32285, LUT_AMPL_WIDTH),
		18176 => to_signed(32285, LUT_AMPL_WIDTH),
		18177 => to_signed(32284, LUT_AMPL_WIDTH),
		18178 => to_signed(32284, LUT_AMPL_WIDTH),
		18179 => to_signed(32283, LUT_AMPL_WIDTH),
		18180 => to_signed(32282, LUT_AMPL_WIDTH),
		18181 => to_signed(32282, LUT_AMPL_WIDTH),
		18182 => to_signed(32281, LUT_AMPL_WIDTH),
		18183 => to_signed(32281, LUT_AMPL_WIDTH),
		18184 => to_signed(32280, LUT_AMPL_WIDTH),
		18185 => to_signed(32280, LUT_AMPL_WIDTH),
		18186 => to_signed(32279, LUT_AMPL_WIDTH),
		18187 => to_signed(32279, LUT_AMPL_WIDTH),
		18188 => to_signed(32278, LUT_AMPL_WIDTH),
		18189 => to_signed(32278, LUT_AMPL_WIDTH),
		18190 => to_signed(32277, LUT_AMPL_WIDTH),
		18191 => to_signed(32277, LUT_AMPL_WIDTH),
		18192 => to_signed(32276, LUT_AMPL_WIDTH),
		18193 => to_signed(32275, LUT_AMPL_WIDTH),
		18194 => to_signed(32275, LUT_AMPL_WIDTH),
		18195 => to_signed(32274, LUT_AMPL_WIDTH),
		18196 => to_signed(32274, LUT_AMPL_WIDTH),
		18197 => to_signed(32273, LUT_AMPL_WIDTH),
		18198 => to_signed(32273, LUT_AMPL_WIDTH),
		18199 => to_signed(32272, LUT_AMPL_WIDTH),
		18200 => to_signed(32272, LUT_AMPL_WIDTH),
		18201 => to_signed(32271, LUT_AMPL_WIDTH),
		18202 => to_signed(32271, LUT_AMPL_WIDTH),
		18203 => to_signed(32270, LUT_AMPL_WIDTH),
		18204 => to_signed(32269, LUT_AMPL_WIDTH),
		18205 => to_signed(32269, LUT_AMPL_WIDTH),
		18206 => to_signed(32268, LUT_AMPL_WIDTH),
		18207 => to_signed(32268, LUT_AMPL_WIDTH),
		18208 => to_signed(32267, LUT_AMPL_WIDTH),
		18209 => to_signed(32267, LUT_AMPL_WIDTH),
		18210 => to_signed(32266, LUT_AMPL_WIDTH),
		18211 => to_signed(32266, LUT_AMPL_WIDTH),
		18212 => to_signed(32265, LUT_AMPL_WIDTH),
		18213 => to_signed(32265, LUT_AMPL_WIDTH),
		18214 => to_signed(32264, LUT_AMPL_WIDTH),
		18215 => to_signed(32263, LUT_AMPL_WIDTH),
		18216 => to_signed(32263, LUT_AMPL_WIDTH),
		18217 => to_signed(32262, LUT_AMPL_WIDTH),
		18218 => to_signed(32262, LUT_AMPL_WIDTH),
		18219 => to_signed(32261, LUT_AMPL_WIDTH),
		18220 => to_signed(32261, LUT_AMPL_WIDTH),
		18221 => to_signed(32260, LUT_AMPL_WIDTH),
		18222 => to_signed(32260, LUT_AMPL_WIDTH),
		18223 => to_signed(32259, LUT_AMPL_WIDTH),
		18224 => to_signed(32258, LUT_AMPL_WIDTH),
		18225 => to_signed(32258, LUT_AMPL_WIDTH),
		18226 => to_signed(32257, LUT_AMPL_WIDTH),
		18227 => to_signed(32257, LUT_AMPL_WIDTH),
		18228 => to_signed(32256, LUT_AMPL_WIDTH),
		18229 => to_signed(32256, LUT_AMPL_WIDTH),
		18230 => to_signed(32255, LUT_AMPL_WIDTH),
		18231 => to_signed(32255, LUT_AMPL_WIDTH),
		18232 => to_signed(32254, LUT_AMPL_WIDTH),
		18233 => to_signed(32253, LUT_AMPL_WIDTH),
		18234 => to_signed(32253, LUT_AMPL_WIDTH),
		18235 => to_signed(32252, LUT_AMPL_WIDTH),
		18236 => to_signed(32252, LUT_AMPL_WIDTH),
		18237 => to_signed(32251, LUT_AMPL_WIDTH),
		18238 => to_signed(32251, LUT_AMPL_WIDTH),
		18239 => to_signed(32250, LUT_AMPL_WIDTH),
		18240 => to_signed(32250, LUT_AMPL_WIDTH),
		18241 => to_signed(32249, LUT_AMPL_WIDTH),
		18242 => to_signed(32248, LUT_AMPL_WIDTH),
		18243 => to_signed(32248, LUT_AMPL_WIDTH),
		18244 => to_signed(32247, LUT_AMPL_WIDTH),
		18245 => to_signed(32247, LUT_AMPL_WIDTH),
		18246 => to_signed(32246, LUT_AMPL_WIDTH),
		18247 => to_signed(32246, LUT_AMPL_WIDTH),
		18248 => to_signed(32245, LUT_AMPL_WIDTH),
		18249 => to_signed(32245, LUT_AMPL_WIDTH),
		18250 => to_signed(32244, LUT_AMPL_WIDTH),
		18251 => to_signed(32243, LUT_AMPL_WIDTH),
		18252 => to_signed(32243, LUT_AMPL_WIDTH),
		18253 => to_signed(32242, LUT_AMPL_WIDTH),
		18254 => to_signed(32242, LUT_AMPL_WIDTH),
		18255 => to_signed(32241, LUT_AMPL_WIDTH),
		18256 => to_signed(32241, LUT_AMPL_WIDTH),
		18257 => to_signed(32240, LUT_AMPL_WIDTH),
		18258 => to_signed(32240, LUT_AMPL_WIDTH),
		18259 => to_signed(32239, LUT_AMPL_WIDTH),
		18260 => to_signed(32238, LUT_AMPL_WIDTH),
		18261 => to_signed(32238, LUT_AMPL_WIDTH),
		18262 => to_signed(32237, LUT_AMPL_WIDTH),
		18263 => to_signed(32237, LUT_AMPL_WIDTH),
		18264 => to_signed(32236, LUT_AMPL_WIDTH),
		18265 => to_signed(32236, LUT_AMPL_WIDTH),
		18266 => to_signed(32235, LUT_AMPL_WIDTH),
		18267 => to_signed(32234, LUT_AMPL_WIDTH),
		18268 => to_signed(32234, LUT_AMPL_WIDTH),
		18269 => to_signed(32233, LUT_AMPL_WIDTH),
		18270 => to_signed(32233, LUT_AMPL_WIDTH),
		18271 => to_signed(32232, LUT_AMPL_WIDTH),
		18272 => to_signed(32232, LUT_AMPL_WIDTH),
		18273 => to_signed(32231, LUT_AMPL_WIDTH),
		18274 => to_signed(32231, LUT_AMPL_WIDTH),
		18275 => to_signed(32230, LUT_AMPL_WIDTH),
		18276 => to_signed(32229, LUT_AMPL_WIDTH),
		18277 => to_signed(32229, LUT_AMPL_WIDTH),
		18278 => to_signed(32228, LUT_AMPL_WIDTH),
		18279 => to_signed(32228, LUT_AMPL_WIDTH),
		18280 => to_signed(32227, LUT_AMPL_WIDTH),
		18281 => to_signed(32227, LUT_AMPL_WIDTH),
		18282 => to_signed(32226, LUT_AMPL_WIDTH),
		18283 => to_signed(32225, LUT_AMPL_WIDTH),
		18284 => to_signed(32225, LUT_AMPL_WIDTH),
		18285 => to_signed(32224, LUT_AMPL_WIDTH),
		18286 => to_signed(32224, LUT_AMPL_WIDTH),
		18287 => to_signed(32223, LUT_AMPL_WIDTH),
		18288 => to_signed(32223, LUT_AMPL_WIDTH),
		18289 => to_signed(32222, LUT_AMPL_WIDTH),
		18290 => to_signed(32221, LUT_AMPL_WIDTH),
		18291 => to_signed(32221, LUT_AMPL_WIDTH),
		18292 => to_signed(32220, LUT_AMPL_WIDTH),
		18293 => to_signed(32220, LUT_AMPL_WIDTH),
		18294 => to_signed(32219, LUT_AMPL_WIDTH),
		18295 => to_signed(32219, LUT_AMPL_WIDTH),
		18296 => to_signed(32218, LUT_AMPL_WIDTH),
		18297 => to_signed(32217, LUT_AMPL_WIDTH),
		18298 => to_signed(32217, LUT_AMPL_WIDTH),
		18299 => to_signed(32216, LUT_AMPL_WIDTH),
		18300 => to_signed(32216, LUT_AMPL_WIDTH),
		18301 => to_signed(32215, LUT_AMPL_WIDTH),
		18302 => to_signed(32215, LUT_AMPL_WIDTH),
		18303 => to_signed(32214, LUT_AMPL_WIDTH),
		18304 => to_signed(32213, LUT_AMPL_WIDTH),
		18305 => to_signed(32213, LUT_AMPL_WIDTH),
		18306 => to_signed(32212, LUT_AMPL_WIDTH),
		18307 => to_signed(32212, LUT_AMPL_WIDTH),
		18308 => to_signed(32211, LUT_AMPL_WIDTH),
		18309 => to_signed(32211, LUT_AMPL_WIDTH),
		18310 => to_signed(32210, LUT_AMPL_WIDTH),
		18311 => to_signed(32209, LUT_AMPL_WIDTH),
		18312 => to_signed(32209, LUT_AMPL_WIDTH),
		18313 => to_signed(32208, LUT_AMPL_WIDTH),
		18314 => to_signed(32208, LUT_AMPL_WIDTH),
		18315 => to_signed(32207, LUT_AMPL_WIDTH),
		18316 => to_signed(32206, LUT_AMPL_WIDTH),
		18317 => to_signed(32206, LUT_AMPL_WIDTH),
		18318 => to_signed(32205, LUT_AMPL_WIDTH),
		18319 => to_signed(32205, LUT_AMPL_WIDTH),
		18320 => to_signed(32204, LUT_AMPL_WIDTH),
		18321 => to_signed(32204, LUT_AMPL_WIDTH),
		18322 => to_signed(32203, LUT_AMPL_WIDTH),
		18323 => to_signed(32202, LUT_AMPL_WIDTH),
		18324 => to_signed(32202, LUT_AMPL_WIDTH),
		18325 => to_signed(32201, LUT_AMPL_WIDTH),
		18326 => to_signed(32201, LUT_AMPL_WIDTH),
		18327 => to_signed(32200, LUT_AMPL_WIDTH),
		18328 => to_signed(32200, LUT_AMPL_WIDTH),
		18329 => to_signed(32199, LUT_AMPL_WIDTH),
		18330 => to_signed(32198, LUT_AMPL_WIDTH),
		18331 => to_signed(32198, LUT_AMPL_WIDTH),
		18332 => to_signed(32197, LUT_AMPL_WIDTH),
		18333 => to_signed(32197, LUT_AMPL_WIDTH),
		18334 => to_signed(32196, LUT_AMPL_WIDTH),
		18335 => to_signed(32195, LUT_AMPL_WIDTH),
		18336 => to_signed(32195, LUT_AMPL_WIDTH),
		18337 => to_signed(32194, LUT_AMPL_WIDTH),
		18338 => to_signed(32194, LUT_AMPL_WIDTH),
		18339 => to_signed(32193, LUT_AMPL_WIDTH),
		18340 => to_signed(32193, LUT_AMPL_WIDTH),
		18341 => to_signed(32192, LUT_AMPL_WIDTH),
		18342 => to_signed(32191, LUT_AMPL_WIDTH),
		18343 => to_signed(32191, LUT_AMPL_WIDTH),
		18344 => to_signed(32190, LUT_AMPL_WIDTH),
		18345 => to_signed(32190, LUT_AMPL_WIDTH),
		18346 => to_signed(32189, LUT_AMPL_WIDTH),
		18347 => to_signed(32188, LUT_AMPL_WIDTH),
		18348 => to_signed(32188, LUT_AMPL_WIDTH),
		18349 => to_signed(32187, LUT_AMPL_WIDTH),
		18350 => to_signed(32187, LUT_AMPL_WIDTH),
		18351 => to_signed(32186, LUT_AMPL_WIDTH),
		18352 => to_signed(32185, LUT_AMPL_WIDTH),
		18353 => to_signed(32185, LUT_AMPL_WIDTH),
		18354 => to_signed(32184, LUT_AMPL_WIDTH),
		18355 => to_signed(32184, LUT_AMPL_WIDTH),
		18356 => to_signed(32183, LUT_AMPL_WIDTH),
		18357 => to_signed(32183, LUT_AMPL_WIDTH),
		18358 => to_signed(32182, LUT_AMPL_WIDTH),
		18359 => to_signed(32181, LUT_AMPL_WIDTH),
		18360 => to_signed(32181, LUT_AMPL_WIDTH),
		18361 => to_signed(32180, LUT_AMPL_WIDTH),
		18362 => to_signed(32180, LUT_AMPL_WIDTH),
		18363 => to_signed(32179, LUT_AMPL_WIDTH),
		18364 => to_signed(32178, LUT_AMPL_WIDTH),
		18365 => to_signed(32178, LUT_AMPL_WIDTH),
		18366 => to_signed(32177, LUT_AMPL_WIDTH),
		18367 => to_signed(32177, LUT_AMPL_WIDTH),
		18368 => to_signed(32176, LUT_AMPL_WIDTH),
		18369 => to_signed(32175, LUT_AMPL_WIDTH),
		18370 => to_signed(32175, LUT_AMPL_WIDTH),
		18371 => to_signed(32174, LUT_AMPL_WIDTH),
		18372 => to_signed(32174, LUT_AMPL_WIDTH),
		18373 => to_signed(32173, LUT_AMPL_WIDTH),
		18374 => to_signed(32172, LUT_AMPL_WIDTH),
		18375 => to_signed(32172, LUT_AMPL_WIDTH),
		18376 => to_signed(32171, LUT_AMPL_WIDTH),
		18377 => to_signed(32171, LUT_AMPL_WIDTH),
		18378 => to_signed(32170, LUT_AMPL_WIDTH),
		18379 => to_signed(32169, LUT_AMPL_WIDTH),
		18380 => to_signed(32169, LUT_AMPL_WIDTH),
		18381 => to_signed(32168, LUT_AMPL_WIDTH),
		18382 => to_signed(32168, LUT_AMPL_WIDTH),
		18383 => to_signed(32167, LUT_AMPL_WIDTH),
		18384 => to_signed(32166, LUT_AMPL_WIDTH),
		18385 => to_signed(32166, LUT_AMPL_WIDTH),
		18386 => to_signed(32165, LUT_AMPL_WIDTH),
		18387 => to_signed(32165, LUT_AMPL_WIDTH),
		18388 => to_signed(32164, LUT_AMPL_WIDTH),
		18389 => to_signed(32163, LUT_AMPL_WIDTH),
		18390 => to_signed(32163, LUT_AMPL_WIDTH),
		18391 => to_signed(32162, LUT_AMPL_WIDTH),
		18392 => to_signed(32162, LUT_AMPL_WIDTH),
		18393 => to_signed(32161, LUT_AMPL_WIDTH),
		18394 => to_signed(32160, LUT_AMPL_WIDTH),
		18395 => to_signed(32160, LUT_AMPL_WIDTH),
		18396 => to_signed(32159, LUT_AMPL_WIDTH),
		18397 => to_signed(32159, LUT_AMPL_WIDTH),
		18398 => to_signed(32158, LUT_AMPL_WIDTH),
		18399 => to_signed(32157, LUT_AMPL_WIDTH),
		18400 => to_signed(32157, LUT_AMPL_WIDTH),
		18401 => to_signed(32156, LUT_AMPL_WIDTH),
		18402 => to_signed(32156, LUT_AMPL_WIDTH),
		18403 => to_signed(32155, LUT_AMPL_WIDTH),
		18404 => to_signed(32154, LUT_AMPL_WIDTH),
		18405 => to_signed(32154, LUT_AMPL_WIDTH),
		18406 => to_signed(32153, LUT_AMPL_WIDTH),
		18407 => to_signed(32153, LUT_AMPL_WIDTH),
		18408 => to_signed(32152, LUT_AMPL_WIDTH),
		18409 => to_signed(32151, LUT_AMPL_WIDTH),
		18410 => to_signed(32151, LUT_AMPL_WIDTH),
		18411 => to_signed(32150, LUT_AMPL_WIDTH),
		18412 => to_signed(32150, LUT_AMPL_WIDTH),
		18413 => to_signed(32149, LUT_AMPL_WIDTH),
		18414 => to_signed(32148, LUT_AMPL_WIDTH),
		18415 => to_signed(32148, LUT_AMPL_WIDTH),
		18416 => to_signed(32147, LUT_AMPL_WIDTH),
		18417 => to_signed(32147, LUT_AMPL_WIDTH),
		18418 => to_signed(32146, LUT_AMPL_WIDTH),
		18419 => to_signed(32145, LUT_AMPL_WIDTH),
		18420 => to_signed(32145, LUT_AMPL_WIDTH),
		18421 => to_signed(32144, LUT_AMPL_WIDTH),
		18422 => to_signed(32144, LUT_AMPL_WIDTH),
		18423 => to_signed(32143, LUT_AMPL_WIDTH),
		18424 => to_signed(32142, LUT_AMPL_WIDTH),
		18425 => to_signed(32142, LUT_AMPL_WIDTH),
		18426 => to_signed(32141, LUT_AMPL_WIDTH),
		18427 => to_signed(32140, LUT_AMPL_WIDTH),
		18428 => to_signed(32140, LUT_AMPL_WIDTH),
		18429 => to_signed(32139, LUT_AMPL_WIDTH),
		18430 => to_signed(32139, LUT_AMPL_WIDTH),
		18431 => to_signed(32138, LUT_AMPL_WIDTH),
		18432 => to_signed(32137, LUT_AMPL_WIDTH),
		18433 => to_signed(32137, LUT_AMPL_WIDTH),
		18434 => to_signed(32136, LUT_AMPL_WIDTH),
		18435 => to_signed(32136, LUT_AMPL_WIDTH),
		18436 => to_signed(32135, LUT_AMPL_WIDTH),
		18437 => to_signed(32134, LUT_AMPL_WIDTH),
		18438 => to_signed(32134, LUT_AMPL_WIDTH),
		18439 => to_signed(32133, LUT_AMPL_WIDTH),
		18440 => to_signed(32132, LUT_AMPL_WIDTH),
		18441 => to_signed(32132, LUT_AMPL_WIDTH),
		18442 => to_signed(32131, LUT_AMPL_WIDTH),
		18443 => to_signed(32131, LUT_AMPL_WIDTH),
		18444 => to_signed(32130, LUT_AMPL_WIDTH),
		18445 => to_signed(32129, LUT_AMPL_WIDTH),
		18446 => to_signed(32129, LUT_AMPL_WIDTH),
		18447 => to_signed(32128, LUT_AMPL_WIDTH),
		18448 => to_signed(32128, LUT_AMPL_WIDTH),
		18449 => to_signed(32127, LUT_AMPL_WIDTH),
		18450 => to_signed(32126, LUT_AMPL_WIDTH),
		18451 => to_signed(32126, LUT_AMPL_WIDTH),
		18452 => to_signed(32125, LUT_AMPL_WIDTH),
		18453 => to_signed(32124, LUT_AMPL_WIDTH),
		18454 => to_signed(32124, LUT_AMPL_WIDTH),
		18455 => to_signed(32123, LUT_AMPL_WIDTH),
		18456 => to_signed(32123, LUT_AMPL_WIDTH),
		18457 => to_signed(32122, LUT_AMPL_WIDTH),
		18458 => to_signed(32121, LUT_AMPL_WIDTH),
		18459 => to_signed(32121, LUT_AMPL_WIDTH),
		18460 => to_signed(32120, LUT_AMPL_WIDTH),
		18461 => to_signed(32119, LUT_AMPL_WIDTH),
		18462 => to_signed(32119, LUT_AMPL_WIDTH),
		18463 => to_signed(32118, LUT_AMPL_WIDTH),
		18464 => to_signed(32118, LUT_AMPL_WIDTH),
		18465 => to_signed(32117, LUT_AMPL_WIDTH),
		18466 => to_signed(32116, LUT_AMPL_WIDTH),
		18467 => to_signed(32116, LUT_AMPL_WIDTH),
		18468 => to_signed(32115, LUT_AMPL_WIDTH),
		18469 => to_signed(32115, LUT_AMPL_WIDTH),
		18470 => to_signed(32114, LUT_AMPL_WIDTH),
		18471 => to_signed(32113, LUT_AMPL_WIDTH),
		18472 => to_signed(32113, LUT_AMPL_WIDTH),
		18473 => to_signed(32112, LUT_AMPL_WIDTH),
		18474 => to_signed(32111, LUT_AMPL_WIDTH),
		18475 => to_signed(32111, LUT_AMPL_WIDTH),
		18476 => to_signed(32110, LUT_AMPL_WIDTH),
		18477 => to_signed(32110, LUT_AMPL_WIDTH),
		18478 => to_signed(32109, LUT_AMPL_WIDTH),
		18479 => to_signed(32108, LUT_AMPL_WIDTH),
		18480 => to_signed(32108, LUT_AMPL_WIDTH),
		18481 => to_signed(32107, LUT_AMPL_WIDTH),
		18482 => to_signed(32106, LUT_AMPL_WIDTH),
		18483 => to_signed(32106, LUT_AMPL_WIDTH),
		18484 => to_signed(32105, LUT_AMPL_WIDTH),
		18485 => to_signed(32104, LUT_AMPL_WIDTH),
		18486 => to_signed(32104, LUT_AMPL_WIDTH),
		18487 => to_signed(32103, LUT_AMPL_WIDTH),
		18488 => to_signed(32103, LUT_AMPL_WIDTH),
		18489 => to_signed(32102, LUT_AMPL_WIDTH),
		18490 => to_signed(32101, LUT_AMPL_WIDTH),
		18491 => to_signed(32101, LUT_AMPL_WIDTH),
		18492 => to_signed(32100, LUT_AMPL_WIDTH),
		18493 => to_signed(32099, LUT_AMPL_WIDTH),
		18494 => to_signed(32099, LUT_AMPL_WIDTH),
		18495 => to_signed(32098, LUT_AMPL_WIDTH),
		18496 => to_signed(32098, LUT_AMPL_WIDTH),
		18497 => to_signed(32097, LUT_AMPL_WIDTH),
		18498 => to_signed(32096, LUT_AMPL_WIDTH),
		18499 => to_signed(32096, LUT_AMPL_WIDTH),
		18500 => to_signed(32095, LUT_AMPL_WIDTH),
		18501 => to_signed(32094, LUT_AMPL_WIDTH),
		18502 => to_signed(32094, LUT_AMPL_WIDTH),
		18503 => to_signed(32093, LUT_AMPL_WIDTH),
		18504 => to_signed(32092, LUT_AMPL_WIDTH),
		18505 => to_signed(32092, LUT_AMPL_WIDTH),
		18506 => to_signed(32091, LUT_AMPL_WIDTH),
		18507 => to_signed(32091, LUT_AMPL_WIDTH),
		18508 => to_signed(32090, LUT_AMPL_WIDTH),
		18509 => to_signed(32089, LUT_AMPL_WIDTH),
		18510 => to_signed(32089, LUT_AMPL_WIDTH),
		18511 => to_signed(32088, LUT_AMPL_WIDTH),
		18512 => to_signed(32087, LUT_AMPL_WIDTH),
		18513 => to_signed(32087, LUT_AMPL_WIDTH),
		18514 => to_signed(32086, LUT_AMPL_WIDTH),
		18515 => to_signed(32086, LUT_AMPL_WIDTH),
		18516 => to_signed(32085, LUT_AMPL_WIDTH),
		18517 => to_signed(32084, LUT_AMPL_WIDTH),
		18518 => to_signed(32084, LUT_AMPL_WIDTH),
		18519 => to_signed(32083, LUT_AMPL_WIDTH),
		18520 => to_signed(32082, LUT_AMPL_WIDTH),
		18521 => to_signed(32082, LUT_AMPL_WIDTH),
		18522 => to_signed(32081, LUT_AMPL_WIDTH),
		18523 => to_signed(32080, LUT_AMPL_WIDTH),
		18524 => to_signed(32080, LUT_AMPL_WIDTH),
		18525 => to_signed(32079, LUT_AMPL_WIDTH),
		18526 => to_signed(32078, LUT_AMPL_WIDTH),
		18527 => to_signed(32078, LUT_AMPL_WIDTH),
		18528 => to_signed(32077, LUT_AMPL_WIDTH),
		18529 => to_signed(32077, LUT_AMPL_WIDTH),
		18530 => to_signed(32076, LUT_AMPL_WIDTH),
		18531 => to_signed(32075, LUT_AMPL_WIDTH),
		18532 => to_signed(32075, LUT_AMPL_WIDTH),
		18533 => to_signed(32074, LUT_AMPL_WIDTH),
		18534 => to_signed(32073, LUT_AMPL_WIDTH),
		18535 => to_signed(32073, LUT_AMPL_WIDTH),
		18536 => to_signed(32072, LUT_AMPL_WIDTH),
		18537 => to_signed(32071, LUT_AMPL_WIDTH),
		18538 => to_signed(32071, LUT_AMPL_WIDTH),
		18539 => to_signed(32070, LUT_AMPL_WIDTH),
		18540 => to_signed(32069, LUT_AMPL_WIDTH),
		18541 => to_signed(32069, LUT_AMPL_WIDTH),
		18542 => to_signed(32068, LUT_AMPL_WIDTH),
		18543 => to_signed(32068, LUT_AMPL_WIDTH),
		18544 => to_signed(32067, LUT_AMPL_WIDTH),
		18545 => to_signed(32066, LUT_AMPL_WIDTH),
		18546 => to_signed(32066, LUT_AMPL_WIDTH),
		18547 => to_signed(32065, LUT_AMPL_WIDTH),
		18548 => to_signed(32064, LUT_AMPL_WIDTH),
		18549 => to_signed(32064, LUT_AMPL_WIDTH),
		18550 => to_signed(32063, LUT_AMPL_WIDTH),
		18551 => to_signed(32062, LUT_AMPL_WIDTH),
		18552 => to_signed(32062, LUT_AMPL_WIDTH),
		18553 => to_signed(32061, LUT_AMPL_WIDTH),
		18554 => to_signed(32060, LUT_AMPL_WIDTH),
		18555 => to_signed(32060, LUT_AMPL_WIDTH),
		18556 => to_signed(32059, LUT_AMPL_WIDTH),
		18557 => to_signed(32058, LUT_AMPL_WIDTH),
		18558 => to_signed(32058, LUT_AMPL_WIDTH),
		18559 => to_signed(32057, LUT_AMPL_WIDTH),
		18560 => to_signed(32057, LUT_AMPL_WIDTH),
		18561 => to_signed(32056, LUT_AMPL_WIDTH),
		18562 => to_signed(32055, LUT_AMPL_WIDTH),
		18563 => to_signed(32055, LUT_AMPL_WIDTH),
		18564 => to_signed(32054, LUT_AMPL_WIDTH),
		18565 => to_signed(32053, LUT_AMPL_WIDTH),
		18566 => to_signed(32053, LUT_AMPL_WIDTH),
		18567 => to_signed(32052, LUT_AMPL_WIDTH),
		18568 => to_signed(32051, LUT_AMPL_WIDTH),
		18569 => to_signed(32051, LUT_AMPL_WIDTH),
		18570 => to_signed(32050, LUT_AMPL_WIDTH),
		18571 => to_signed(32049, LUT_AMPL_WIDTH),
		18572 => to_signed(32049, LUT_AMPL_WIDTH),
		18573 => to_signed(32048, LUT_AMPL_WIDTH),
		18574 => to_signed(32047, LUT_AMPL_WIDTH),
		18575 => to_signed(32047, LUT_AMPL_WIDTH),
		18576 => to_signed(32046, LUT_AMPL_WIDTH),
		18577 => to_signed(32045, LUT_AMPL_WIDTH),
		18578 => to_signed(32045, LUT_AMPL_WIDTH),
		18579 => to_signed(32044, LUT_AMPL_WIDTH),
		18580 => to_signed(32043, LUT_AMPL_WIDTH),
		18581 => to_signed(32043, LUT_AMPL_WIDTH),
		18582 => to_signed(32042, LUT_AMPL_WIDTH),
		18583 => to_signed(32041, LUT_AMPL_WIDTH),
		18584 => to_signed(32041, LUT_AMPL_WIDTH),
		18585 => to_signed(32040, LUT_AMPL_WIDTH),
		18586 => to_signed(32040, LUT_AMPL_WIDTH),
		18587 => to_signed(32039, LUT_AMPL_WIDTH),
		18588 => to_signed(32038, LUT_AMPL_WIDTH),
		18589 => to_signed(32038, LUT_AMPL_WIDTH),
		18590 => to_signed(32037, LUT_AMPL_WIDTH),
		18591 => to_signed(32036, LUT_AMPL_WIDTH),
		18592 => to_signed(32036, LUT_AMPL_WIDTH),
		18593 => to_signed(32035, LUT_AMPL_WIDTH),
		18594 => to_signed(32034, LUT_AMPL_WIDTH),
		18595 => to_signed(32034, LUT_AMPL_WIDTH),
		18596 => to_signed(32033, LUT_AMPL_WIDTH),
		18597 => to_signed(32032, LUT_AMPL_WIDTH),
		18598 => to_signed(32032, LUT_AMPL_WIDTH),
		18599 => to_signed(32031, LUT_AMPL_WIDTH),
		18600 => to_signed(32030, LUT_AMPL_WIDTH),
		18601 => to_signed(32030, LUT_AMPL_WIDTH),
		18602 => to_signed(32029, LUT_AMPL_WIDTH),
		18603 => to_signed(32028, LUT_AMPL_WIDTH),
		18604 => to_signed(32028, LUT_AMPL_WIDTH),
		18605 => to_signed(32027, LUT_AMPL_WIDTH),
		18606 => to_signed(32026, LUT_AMPL_WIDTH),
		18607 => to_signed(32026, LUT_AMPL_WIDTH),
		18608 => to_signed(32025, LUT_AMPL_WIDTH),
		18609 => to_signed(32024, LUT_AMPL_WIDTH),
		18610 => to_signed(32024, LUT_AMPL_WIDTH),
		18611 => to_signed(32023, LUT_AMPL_WIDTH),
		18612 => to_signed(32022, LUT_AMPL_WIDTH),
		18613 => to_signed(32022, LUT_AMPL_WIDTH),
		18614 => to_signed(32021, LUT_AMPL_WIDTH),
		18615 => to_signed(32020, LUT_AMPL_WIDTH),
		18616 => to_signed(32020, LUT_AMPL_WIDTH),
		18617 => to_signed(32019, LUT_AMPL_WIDTH),
		18618 => to_signed(32018, LUT_AMPL_WIDTH),
		18619 => to_signed(32018, LUT_AMPL_WIDTH),
		18620 => to_signed(32017, LUT_AMPL_WIDTH),
		18621 => to_signed(32016, LUT_AMPL_WIDTH),
		18622 => to_signed(32016, LUT_AMPL_WIDTH),
		18623 => to_signed(32015, LUT_AMPL_WIDTH),
		18624 => to_signed(32014, LUT_AMPL_WIDTH),
		18625 => to_signed(32014, LUT_AMPL_WIDTH),
		18626 => to_signed(32013, LUT_AMPL_WIDTH),
		18627 => to_signed(32012, LUT_AMPL_WIDTH),
		18628 => to_signed(32012, LUT_AMPL_WIDTH),
		18629 => to_signed(32011, LUT_AMPL_WIDTH),
		18630 => to_signed(32010, LUT_AMPL_WIDTH),
		18631 => to_signed(32010, LUT_AMPL_WIDTH),
		18632 => to_signed(32009, LUT_AMPL_WIDTH),
		18633 => to_signed(32008, LUT_AMPL_WIDTH),
		18634 => to_signed(32008, LUT_AMPL_WIDTH),
		18635 => to_signed(32007, LUT_AMPL_WIDTH),
		18636 => to_signed(32006, LUT_AMPL_WIDTH),
		18637 => to_signed(32006, LUT_AMPL_WIDTH),
		18638 => to_signed(32005, LUT_AMPL_WIDTH),
		18639 => to_signed(32004, LUT_AMPL_WIDTH),
		18640 => to_signed(32004, LUT_AMPL_WIDTH),
		18641 => to_signed(32003, LUT_AMPL_WIDTH),
		18642 => to_signed(32002, LUT_AMPL_WIDTH),
		18643 => to_signed(32002, LUT_AMPL_WIDTH),
		18644 => to_signed(32001, LUT_AMPL_WIDTH),
		18645 => to_signed(32000, LUT_AMPL_WIDTH),
		18646 => to_signed(31999, LUT_AMPL_WIDTH),
		18647 => to_signed(31999, LUT_AMPL_WIDTH),
		18648 => to_signed(31998, LUT_AMPL_WIDTH),
		18649 => to_signed(31997, LUT_AMPL_WIDTH),
		18650 => to_signed(31997, LUT_AMPL_WIDTH),
		18651 => to_signed(31996, LUT_AMPL_WIDTH),
		18652 => to_signed(31995, LUT_AMPL_WIDTH),
		18653 => to_signed(31995, LUT_AMPL_WIDTH),
		18654 => to_signed(31994, LUT_AMPL_WIDTH),
		18655 => to_signed(31993, LUT_AMPL_WIDTH),
		18656 => to_signed(31993, LUT_AMPL_WIDTH),
		18657 => to_signed(31992, LUT_AMPL_WIDTH),
		18658 => to_signed(31991, LUT_AMPL_WIDTH),
		18659 => to_signed(31991, LUT_AMPL_WIDTH),
		18660 => to_signed(31990, LUT_AMPL_WIDTH),
		18661 => to_signed(31989, LUT_AMPL_WIDTH),
		18662 => to_signed(31989, LUT_AMPL_WIDTH),
		18663 => to_signed(31988, LUT_AMPL_WIDTH),
		18664 => to_signed(31987, LUT_AMPL_WIDTH),
		18665 => to_signed(31987, LUT_AMPL_WIDTH),
		18666 => to_signed(31986, LUT_AMPL_WIDTH),
		18667 => to_signed(31985, LUT_AMPL_WIDTH),
		18668 => to_signed(31985, LUT_AMPL_WIDTH),
		18669 => to_signed(31984, LUT_AMPL_WIDTH),
		18670 => to_signed(31983, LUT_AMPL_WIDTH),
		18671 => to_signed(31982, LUT_AMPL_WIDTH),
		18672 => to_signed(31982, LUT_AMPL_WIDTH),
		18673 => to_signed(31981, LUT_AMPL_WIDTH),
		18674 => to_signed(31980, LUT_AMPL_WIDTH),
		18675 => to_signed(31980, LUT_AMPL_WIDTH),
		18676 => to_signed(31979, LUT_AMPL_WIDTH),
		18677 => to_signed(31978, LUT_AMPL_WIDTH),
		18678 => to_signed(31978, LUT_AMPL_WIDTH),
		18679 => to_signed(31977, LUT_AMPL_WIDTH),
		18680 => to_signed(31976, LUT_AMPL_WIDTH),
		18681 => to_signed(31976, LUT_AMPL_WIDTH),
		18682 => to_signed(31975, LUT_AMPL_WIDTH),
		18683 => to_signed(31974, LUT_AMPL_WIDTH),
		18684 => to_signed(31974, LUT_AMPL_WIDTH),
		18685 => to_signed(31973, LUT_AMPL_WIDTH),
		18686 => to_signed(31972, LUT_AMPL_WIDTH),
		18687 => to_signed(31972, LUT_AMPL_WIDTH),
		18688 => to_signed(31971, LUT_AMPL_WIDTH),
		18689 => to_signed(31970, LUT_AMPL_WIDTH),
		18690 => to_signed(31969, LUT_AMPL_WIDTH),
		18691 => to_signed(31969, LUT_AMPL_WIDTH),
		18692 => to_signed(31968, LUT_AMPL_WIDTH),
		18693 => to_signed(31967, LUT_AMPL_WIDTH),
		18694 => to_signed(31967, LUT_AMPL_WIDTH),
		18695 => to_signed(31966, LUT_AMPL_WIDTH),
		18696 => to_signed(31965, LUT_AMPL_WIDTH),
		18697 => to_signed(31965, LUT_AMPL_WIDTH),
		18698 => to_signed(31964, LUT_AMPL_WIDTH),
		18699 => to_signed(31963, LUT_AMPL_WIDTH),
		18700 => to_signed(31963, LUT_AMPL_WIDTH),
		18701 => to_signed(31962, LUT_AMPL_WIDTH),
		18702 => to_signed(31961, LUT_AMPL_WIDTH),
		18703 => to_signed(31960, LUT_AMPL_WIDTH),
		18704 => to_signed(31960, LUT_AMPL_WIDTH),
		18705 => to_signed(31959, LUT_AMPL_WIDTH),
		18706 => to_signed(31958, LUT_AMPL_WIDTH),
		18707 => to_signed(31958, LUT_AMPL_WIDTH),
		18708 => to_signed(31957, LUT_AMPL_WIDTH),
		18709 => to_signed(31956, LUT_AMPL_WIDTH),
		18710 => to_signed(31956, LUT_AMPL_WIDTH),
		18711 => to_signed(31955, LUT_AMPL_WIDTH),
		18712 => to_signed(31954, LUT_AMPL_WIDTH),
		18713 => to_signed(31954, LUT_AMPL_WIDTH),
		18714 => to_signed(31953, LUT_AMPL_WIDTH),
		18715 => to_signed(31952, LUT_AMPL_WIDTH),
		18716 => to_signed(31951, LUT_AMPL_WIDTH),
		18717 => to_signed(31951, LUT_AMPL_WIDTH),
		18718 => to_signed(31950, LUT_AMPL_WIDTH),
		18719 => to_signed(31949, LUT_AMPL_WIDTH),
		18720 => to_signed(31949, LUT_AMPL_WIDTH),
		18721 => to_signed(31948, LUT_AMPL_WIDTH),
		18722 => to_signed(31947, LUT_AMPL_WIDTH),
		18723 => to_signed(31947, LUT_AMPL_WIDTH),
		18724 => to_signed(31946, LUT_AMPL_WIDTH),
		18725 => to_signed(31945, LUT_AMPL_WIDTH),
		18726 => to_signed(31944, LUT_AMPL_WIDTH),
		18727 => to_signed(31944, LUT_AMPL_WIDTH),
		18728 => to_signed(31943, LUT_AMPL_WIDTH),
		18729 => to_signed(31942, LUT_AMPL_WIDTH),
		18730 => to_signed(31942, LUT_AMPL_WIDTH),
		18731 => to_signed(31941, LUT_AMPL_WIDTH),
		18732 => to_signed(31940, LUT_AMPL_WIDTH),
		18733 => to_signed(31940, LUT_AMPL_WIDTH),
		18734 => to_signed(31939, LUT_AMPL_WIDTH),
		18735 => to_signed(31938, LUT_AMPL_WIDTH),
		18736 => to_signed(31937, LUT_AMPL_WIDTH),
		18737 => to_signed(31937, LUT_AMPL_WIDTH),
		18738 => to_signed(31936, LUT_AMPL_WIDTH),
		18739 => to_signed(31935, LUT_AMPL_WIDTH),
		18740 => to_signed(31935, LUT_AMPL_WIDTH),
		18741 => to_signed(31934, LUT_AMPL_WIDTH),
		18742 => to_signed(31933, LUT_AMPL_WIDTH),
		18743 => to_signed(31933, LUT_AMPL_WIDTH),
		18744 => to_signed(31932, LUT_AMPL_WIDTH),
		18745 => to_signed(31931, LUT_AMPL_WIDTH),
		18746 => to_signed(31930, LUT_AMPL_WIDTH),
		18747 => to_signed(31930, LUT_AMPL_WIDTH),
		18748 => to_signed(31929, LUT_AMPL_WIDTH),
		18749 => to_signed(31928, LUT_AMPL_WIDTH),
		18750 => to_signed(31928, LUT_AMPL_WIDTH),
		18751 => to_signed(31927, LUT_AMPL_WIDTH),
		18752 => to_signed(31926, LUT_AMPL_WIDTH),
		18753 => to_signed(31925, LUT_AMPL_WIDTH),
		18754 => to_signed(31925, LUT_AMPL_WIDTH),
		18755 => to_signed(31924, LUT_AMPL_WIDTH),
		18756 => to_signed(31923, LUT_AMPL_WIDTH),
		18757 => to_signed(31923, LUT_AMPL_WIDTH),
		18758 => to_signed(31922, LUT_AMPL_WIDTH),
		18759 => to_signed(31921, LUT_AMPL_WIDTH),
		18760 => to_signed(31921, LUT_AMPL_WIDTH),
		18761 => to_signed(31920, LUT_AMPL_WIDTH),
		18762 => to_signed(31919, LUT_AMPL_WIDTH),
		18763 => to_signed(31918, LUT_AMPL_WIDTH),
		18764 => to_signed(31918, LUT_AMPL_WIDTH),
		18765 => to_signed(31917, LUT_AMPL_WIDTH),
		18766 => to_signed(31916, LUT_AMPL_WIDTH),
		18767 => to_signed(31916, LUT_AMPL_WIDTH),
		18768 => to_signed(31915, LUT_AMPL_WIDTH),
		18769 => to_signed(31914, LUT_AMPL_WIDTH),
		18770 => to_signed(31913, LUT_AMPL_WIDTH),
		18771 => to_signed(31913, LUT_AMPL_WIDTH),
		18772 => to_signed(31912, LUT_AMPL_WIDTH),
		18773 => to_signed(31911, LUT_AMPL_WIDTH),
		18774 => to_signed(31911, LUT_AMPL_WIDTH),
		18775 => to_signed(31910, LUT_AMPL_WIDTH),
		18776 => to_signed(31909, LUT_AMPL_WIDTH),
		18777 => to_signed(31908, LUT_AMPL_WIDTH),
		18778 => to_signed(31908, LUT_AMPL_WIDTH),
		18779 => to_signed(31907, LUT_AMPL_WIDTH),
		18780 => to_signed(31906, LUT_AMPL_WIDTH),
		18781 => to_signed(31906, LUT_AMPL_WIDTH),
		18782 => to_signed(31905, LUT_AMPL_WIDTH),
		18783 => to_signed(31904, LUT_AMPL_WIDTH),
		18784 => to_signed(31903, LUT_AMPL_WIDTH),
		18785 => to_signed(31903, LUT_AMPL_WIDTH),
		18786 => to_signed(31902, LUT_AMPL_WIDTH),
		18787 => to_signed(31901, LUT_AMPL_WIDTH),
		18788 => to_signed(31901, LUT_AMPL_WIDTH),
		18789 => to_signed(31900, LUT_AMPL_WIDTH),
		18790 => to_signed(31899, LUT_AMPL_WIDTH),
		18791 => to_signed(31898, LUT_AMPL_WIDTH),
		18792 => to_signed(31898, LUT_AMPL_WIDTH),
		18793 => to_signed(31897, LUT_AMPL_WIDTH),
		18794 => to_signed(31896, LUT_AMPL_WIDTH),
		18795 => to_signed(31896, LUT_AMPL_WIDTH),
		18796 => to_signed(31895, LUT_AMPL_WIDTH),
		18797 => to_signed(31894, LUT_AMPL_WIDTH),
		18798 => to_signed(31893, LUT_AMPL_WIDTH),
		18799 => to_signed(31893, LUT_AMPL_WIDTH),
		18800 => to_signed(31892, LUT_AMPL_WIDTH),
		18801 => to_signed(31891, LUT_AMPL_WIDTH),
		18802 => to_signed(31890, LUT_AMPL_WIDTH),
		18803 => to_signed(31890, LUT_AMPL_WIDTH),
		18804 => to_signed(31889, LUT_AMPL_WIDTH),
		18805 => to_signed(31888, LUT_AMPL_WIDTH),
		18806 => to_signed(31888, LUT_AMPL_WIDTH),
		18807 => to_signed(31887, LUT_AMPL_WIDTH),
		18808 => to_signed(31886, LUT_AMPL_WIDTH),
		18809 => to_signed(31885, LUT_AMPL_WIDTH),
		18810 => to_signed(31885, LUT_AMPL_WIDTH),
		18811 => to_signed(31884, LUT_AMPL_WIDTH),
		18812 => to_signed(31883, LUT_AMPL_WIDTH),
		18813 => to_signed(31882, LUT_AMPL_WIDTH),
		18814 => to_signed(31882, LUT_AMPL_WIDTH),
		18815 => to_signed(31881, LUT_AMPL_WIDTH),
		18816 => to_signed(31880, LUT_AMPL_WIDTH),
		18817 => to_signed(31880, LUT_AMPL_WIDTH),
		18818 => to_signed(31879, LUT_AMPL_WIDTH),
		18819 => to_signed(31878, LUT_AMPL_WIDTH),
		18820 => to_signed(31877, LUT_AMPL_WIDTH),
		18821 => to_signed(31877, LUT_AMPL_WIDTH),
		18822 => to_signed(31876, LUT_AMPL_WIDTH),
		18823 => to_signed(31875, LUT_AMPL_WIDTH),
		18824 => to_signed(31875, LUT_AMPL_WIDTH),
		18825 => to_signed(31874, LUT_AMPL_WIDTH),
		18826 => to_signed(31873, LUT_AMPL_WIDTH),
		18827 => to_signed(31872, LUT_AMPL_WIDTH),
		18828 => to_signed(31872, LUT_AMPL_WIDTH),
		18829 => to_signed(31871, LUT_AMPL_WIDTH),
		18830 => to_signed(31870, LUT_AMPL_WIDTH),
		18831 => to_signed(31869, LUT_AMPL_WIDTH),
		18832 => to_signed(31869, LUT_AMPL_WIDTH),
		18833 => to_signed(31868, LUT_AMPL_WIDTH),
		18834 => to_signed(31867, LUT_AMPL_WIDTH),
		18835 => to_signed(31866, LUT_AMPL_WIDTH),
		18836 => to_signed(31866, LUT_AMPL_WIDTH),
		18837 => to_signed(31865, LUT_AMPL_WIDTH),
		18838 => to_signed(31864, LUT_AMPL_WIDTH),
		18839 => to_signed(31864, LUT_AMPL_WIDTH),
		18840 => to_signed(31863, LUT_AMPL_WIDTH),
		18841 => to_signed(31862, LUT_AMPL_WIDTH),
		18842 => to_signed(31861, LUT_AMPL_WIDTH),
		18843 => to_signed(31861, LUT_AMPL_WIDTH),
		18844 => to_signed(31860, LUT_AMPL_WIDTH),
		18845 => to_signed(31859, LUT_AMPL_WIDTH),
		18846 => to_signed(31858, LUT_AMPL_WIDTH),
		18847 => to_signed(31858, LUT_AMPL_WIDTH),
		18848 => to_signed(31857, LUT_AMPL_WIDTH),
		18849 => to_signed(31856, LUT_AMPL_WIDTH),
		18850 => to_signed(31855, LUT_AMPL_WIDTH),
		18851 => to_signed(31855, LUT_AMPL_WIDTH),
		18852 => to_signed(31854, LUT_AMPL_WIDTH),
		18853 => to_signed(31853, LUT_AMPL_WIDTH),
		18854 => to_signed(31853, LUT_AMPL_WIDTH),
		18855 => to_signed(31852, LUT_AMPL_WIDTH),
		18856 => to_signed(31851, LUT_AMPL_WIDTH),
		18857 => to_signed(31850, LUT_AMPL_WIDTH),
		18858 => to_signed(31850, LUT_AMPL_WIDTH),
		18859 => to_signed(31849, LUT_AMPL_WIDTH),
		18860 => to_signed(31848, LUT_AMPL_WIDTH),
		18861 => to_signed(31847, LUT_AMPL_WIDTH),
		18862 => to_signed(31847, LUT_AMPL_WIDTH),
		18863 => to_signed(31846, LUT_AMPL_WIDTH),
		18864 => to_signed(31845, LUT_AMPL_WIDTH),
		18865 => to_signed(31844, LUT_AMPL_WIDTH),
		18866 => to_signed(31844, LUT_AMPL_WIDTH),
		18867 => to_signed(31843, LUT_AMPL_WIDTH),
		18868 => to_signed(31842, LUT_AMPL_WIDTH),
		18869 => to_signed(31841, LUT_AMPL_WIDTH),
		18870 => to_signed(31841, LUT_AMPL_WIDTH),
		18871 => to_signed(31840, LUT_AMPL_WIDTH),
		18872 => to_signed(31839, LUT_AMPL_WIDTH),
		18873 => to_signed(31838, LUT_AMPL_WIDTH),
		18874 => to_signed(31838, LUT_AMPL_WIDTH),
		18875 => to_signed(31837, LUT_AMPL_WIDTH),
		18876 => to_signed(31836, LUT_AMPL_WIDTH),
		18877 => to_signed(31836, LUT_AMPL_WIDTH),
		18878 => to_signed(31835, LUT_AMPL_WIDTH),
		18879 => to_signed(31834, LUT_AMPL_WIDTH),
		18880 => to_signed(31833, LUT_AMPL_WIDTH),
		18881 => to_signed(31833, LUT_AMPL_WIDTH),
		18882 => to_signed(31832, LUT_AMPL_WIDTH),
		18883 => to_signed(31831, LUT_AMPL_WIDTH),
		18884 => to_signed(31830, LUT_AMPL_WIDTH),
		18885 => to_signed(31830, LUT_AMPL_WIDTH),
		18886 => to_signed(31829, LUT_AMPL_WIDTH),
		18887 => to_signed(31828, LUT_AMPL_WIDTH),
		18888 => to_signed(31827, LUT_AMPL_WIDTH),
		18889 => to_signed(31827, LUT_AMPL_WIDTH),
		18890 => to_signed(31826, LUT_AMPL_WIDTH),
		18891 => to_signed(31825, LUT_AMPL_WIDTH),
		18892 => to_signed(31824, LUT_AMPL_WIDTH),
		18893 => to_signed(31824, LUT_AMPL_WIDTH),
		18894 => to_signed(31823, LUT_AMPL_WIDTH),
		18895 => to_signed(31822, LUT_AMPL_WIDTH),
		18896 => to_signed(31821, LUT_AMPL_WIDTH),
		18897 => to_signed(31821, LUT_AMPL_WIDTH),
		18898 => to_signed(31820, LUT_AMPL_WIDTH),
		18899 => to_signed(31819, LUT_AMPL_WIDTH),
		18900 => to_signed(31818, LUT_AMPL_WIDTH),
		18901 => to_signed(31818, LUT_AMPL_WIDTH),
		18902 => to_signed(31817, LUT_AMPL_WIDTH),
		18903 => to_signed(31816, LUT_AMPL_WIDTH),
		18904 => to_signed(31815, LUT_AMPL_WIDTH),
		18905 => to_signed(31815, LUT_AMPL_WIDTH),
		18906 => to_signed(31814, LUT_AMPL_WIDTH),
		18907 => to_signed(31813, LUT_AMPL_WIDTH),
		18908 => to_signed(31812, LUT_AMPL_WIDTH),
		18909 => to_signed(31812, LUT_AMPL_WIDTH),
		18910 => to_signed(31811, LUT_AMPL_WIDTH),
		18911 => to_signed(31810, LUT_AMPL_WIDTH),
		18912 => to_signed(31809, LUT_AMPL_WIDTH),
		18913 => to_signed(31809, LUT_AMPL_WIDTH),
		18914 => to_signed(31808, LUT_AMPL_WIDTH),
		18915 => to_signed(31807, LUT_AMPL_WIDTH),
		18916 => to_signed(31806, LUT_AMPL_WIDTH),
		18917 => to_signed(31806, LUT_AMPL_WIDTH),
		18918 => to_signed(31805, LUT_AMPL_WIDTH),
		18919 => to_signed(31804, LUT_AMPL_WIDTH),
		18920 => to_signed(31803, LUT_AMPL_WIDTH),
		18921 => to_signed(31802, LUT_AMPL_WIDTH),
		18922 => to_signed(31802, LUT_AMPL_WIDTH),
		18923 => to_signed(31801, LUT_AMPL_WIDTH),
		18924 => to_signed(31800, LUT_AMPL_WIDTH),
		18925 => to_signed(31799, LUT_AMPL_WIDTH),
		18926 => to_signed(31799, LUT_AMPL_WIDTH),
		18927 => to_signed(31798, LUT_AMPL_WIDTH),
		18928 => to_signed(31797, LUT_AMPL_WIDTH),
		18929 => to_signed(31796, LUT_AMPL_WIDTH),
		18930 => to_signed(31796, LUT_AMPL_WIDTH),
		18931 => to_signed(31795, LUT_AMPL_WIDTH),
		18932 => to_signed(31794, LUT_AMPL_WIDTH),
		18933 => to_signed(31793, LUT_AMPL_WIDTH),
		18934 => to_signed(31793, LUT_AMPL_WIDTH),
		18935 => to_signed(31792, LUT_AMPL_WIDTH),
		18936 => to_signed(31791, LUT_AMPL_WIDTH),
		18937 => to_signed(31790, LUT_AMPL_WIDTH),
		18938 => to_signed(31790, LUT_AMPL_WIDTH),
		18939 => to_signed(31789, LUT_AMPL_WIDTH),
		18940 => to_signed(31788, LUT_AMPL_WIDTH),
		18941 => to_signed(31787, LUT_AMPL_WIDTH),
		18942 => to_signed(31787, LUT_AMPL_WIDTH),
		18943 => to_signed(31786, LUT_AMPL_WIDTH),
		18944 => to_signed(31785, LUT_AMPL_WIDTH),
		18945 => to_signed(31784, LUT_AMPL_WIDTH),
		18946 => to_signed(31783, LUT_AMPL_WIDTH),
		18947 => to_signed(31783, LUT_AMPL_WIDTH),
		18948 => to_signed(31782, LUT_AMPL_WIDTH),
		18949 => to_signed(31781, LUT_AMPL_WIDTH),
		18950 => to_signed(31780, LUT_AMPL_WIDTH),
		18951 => to_signed(31780, LUT_AMPL_WIDTH),
		18952 => to_signed(31779, LUT_AMPL_WIDTH),
		18953 => to_signed(31778, LUT_AMPL_WIDTH),
		18954 => to_signed(31777, LUT_AMPL_WIDTH),
		18955 => to_signed(31777, LUT_AMPL_WIDTH),
		18956 => to_signed(31776, LUT_AMPL_WIDTH),
		18957 => to_signed(31775, LUT_AMPL_WIDTH),
		18958 => to_signed(31774, LUT_AMPL_WIDTH),
		18959 => to_signed(31774, LUT_AMPL_WIDTH),
		18960 => to_signed(31773, LUT_AMPL_WIDTH),
		18961 => to_signed(31772, LUT_AMPL_WIDTH),
		18962 => to_signed(31771, LUT_AMPL_WIDTH),
		18963 => to_signed(31770, LUT_AMPL_WIDTH),
		18964 => to_signed(31770, LUT_AMPL_WIDTH),
		18965 => to_signed(31769, LUT_AMPL_WIDTH),
		18966 => to_signed(31768, LUT_AMPL_WIDTH),
		18967 => to_signed(31767, LUT_AMPL_WIDTH),
		18968 => to_signed(31767, LUT_AMPL_WIDTH),
		18969 => to_signed(31766, LUT_AMPL_WIDTH),
		18970 => to_signed(31765, LUT_AMPL_WIDTH),
		18971 => to_signed(31764, LUT_AMPL_WIDTH),
		18972 => to_signed(31764, LUT_AMPL_WIDTH),
		18973 => to_signed(31763, LUT_AMPL_WIDTH),
		18974 => to_signed(31762, LUT_AMPL_WIDTH),
		18975 => to_signed(31761, LUT_AMPL_WIDTH),
		18976 => to_signed(31760, LUT_AMPL_WIDTH),
		18977 => to_signed(31760, LUT_AMPL_WIDTH),
		18978 => to_signed(31759, LUT_AMPL_WIDTH),
		18979 => to_signed(31758, LUT_AMPL_WIDTH),
		18980 => to_signed(31757, LUT_AMPL_WIDTH),
		18981 => to_signed(31757, LUT_AMPL_WIDTH),
		18982 => to_signed(31756, LUT_AMPL_WIDTH),
		18983 => to_signed(31755, LUT_AMPL_WIDTH),
		18984 => to_signed(31754, LUT_AMPL_WIDTH),
		18985 => to_signed(31753, LUT_AMPL_WIDTH),
		18986 => to_signed(31753, LUT_AMPL_WIDTH),
		18987 => to_signed(31752, LUT_AMPL_WIDTH),
		18988 => to_signed(31751, LUT_AMPL_WIDTH),
		18989 => to_signed(31750, LUT_AMPL_WIDTH),
		18990 => to_signed(31750, LUT_AMPL_WIDTH),
		18991 => to_signed(31749, LUT_AMPL_WIDTH),
		18992 => to_signed(31748, LUT_AMPL_WIDTH),
		18993 => to_signed(31747, LUT_AMPL_WIDTH),
		18994 => to_signed(31746, LUT_AMPL_WIDTH),
		18995 => to_signed(31746, LUT_AMPL_WIDTH),
		18996 => to_signed(31745, LUT_AMPL_WIDTH),
		18997 => to_signed(31744, LUT_AMPL_WIDTH),
		18998 => to_signed(31743, LUT_AMPL_WIDTH),
		18999 => to_signed(31743, LUT_AMPL_WIDTH),
		19000 => to_signed(31742, LUT_AMPL_WIDTH),
		19001 => to_signed(31741, LUT_AMPL_WIDTH),
		19002 => to_signed(31740, LUT_AMPL_WIDTH),
		19003 => to_signed(31739, LUT_AMPL_WIDTH),
		19004 => to_signed(31739, LUT_AMPL_WIDTH),
		19005 => to_signed(31738, LUT_AMPL_WIDTH),
		19006 => to_signed(31737, LUT_AMPL_WIDTH),
		19007 => to_signed(31736, LUT_AMPL_WIDTH),
		19008 => to_signed(31736, LUT_AMPL_WIDTH),
		19009 => to_signed(31735, LUT_AMPL_WIDTH),
		19010 => to_signed(31734, LUT_AMPL_WIDTH),
		19011 => to_signed(31733, LUT_AMPL_WIDTH),
		19012 => to_signed(31732, LUT_AMPL_WIDTH),
		19013 => to_signed(31732, LUT_AMPL_WIDTH),
		19014 => to_signed(31731, LUT_AMPL_WIDTH),
		19015 => to_signed(31730, LUT_AMPL_WIDTH),
		19016 => to_signed(31729, LUT_AMPL_WIDTH),
		19017 => to_signed(31729, LUT_AMPL_WIDTH),
		19018 => to_signed(31728, LUT_AMPL_WIDTH),
		19019 => to_signed(31727, LUT_AMPL_WIDTH),
		19020 => to_signed(31726, LUT_AMPL_WIDTH),
		19021 => to_signed(31725, LUT_AMPL_WIDTH),
		19022 => to_signed(31725, LUT_AMPL_WIDTH),
		19023 => to_signed(31724, LUT_AMPL_WIDTH),
		19024 => to_signed(31723, LUT_AMPL_WIDTH),
		19025 => to_signed(31722, LUT_AMPL_WIDTH),
		19026 => to_signed(31721, LUT_AMPL_WIDTH),
		19027 => to_signed(31721, LUT_AMPL_WIDTH),
		19028 => to_signed(31720, LUT_AMPL_WIDTH),
		19029 => to_signed(31719, LUT_AMPL_WIDTH),
		19030 => to_signed(31718, LUT_AMPL_WIDTH),
		19031 => to_signed(31718, LUT_AMPL_WIDTH),
		19032 => to_signed(31717, LUT_AMPL_WIDTH),
		19033 => to_signed(31716, LUT_AMPL_WIDTH),
		19034 => to_signed(31715, LUT_AMPL_WIDTH),
		19035 => to_signed(31714, LUT_AMPL_WIDTH),
		19036 => to_signed(31714, LUT_AMPL_WIDTH),
		19037 => to_signed(31713, LUT_AMPL_WIDTH),
		19038 => to_signed(31712, LUT_AMPL_WIDTH),
		19039 => to_signed(31711, LUT_AMPL_WIDTH),
		19040 => to_signed(31710, LUT_AMPL_WIDTH),
		19041 => to_signed(31710, LUT_AMPL_WIDTH),
		19042 => to_signed(31709, LUT_AMPL_WIDTH),
		19043 => to_signed(31708, LUT_AMPL_WIDTH),
		19044 => to_signed(31707, LUT_AMPL_WIDTH),
		19045 => to_signed(31706, LUT_AMPL_WIDTH),
		19046 => to_signed(31706, LUT_AMPL_WIDTH),
		19047 => to_signed(31705, LUT_AMPL_WIDTH),
		19048 => to_signed(31704, LUT_AMPL_WIDTH),
		19049 => to_signed(31703, LUT_AMPL_WIDTH),
		19050 => to_signed(31702, LUT_AMPL_WIDTH),
		19051 => to_signed(31702, LUT_AMPL_WIDTH),
		19052 => to_signed(31701, LUT_AMPL_WIDTH),
		19053 => to_signed(31700, LUT_AMPL_WIDTH),
		19054 => to_signed(31699, LUT_AMPL_WIDTH),
		19055 => to_signed(31698, LUT_AMPL_WIDTH),
		19056 => to_signed(31698, LUT_AMPL_WIDTH),
		19057 => to_signed(31697, LUT_AMPL_WIDTH),
		19058 => to_signed(31696, LUT_AMPL_WIDTH),
		19059 => to_signed(31695, LUT_AMPL_WIDTH),
		19060 => to_signed(31695, LUT_AMPL_WIDTH),
		19061 => to_signed(31694, LUT_AMPL_WIDTH),
		19062 => to_signed(31693, LUT_AMPL_WIDTH),
		19063 => to_signed(31692, LUT_AMPL_WIDTH),
		19064 => to_signed(31691, LUT_AMPL_WIDTH),
		19065 => to_signed(31691, LUT_AMPL_WIDTH),
		19066 => to_signed(31690, LUT_AMPL_WIDTH),
		19067 => to_signed(31689, LUT_AMPL_WIDTH),
		19068 => to_signed(31688, LUT_AMPL_WIDTH),
		19069 => to_signed(31687, LUT_AMPL_WIDTH),
		19070 => to_signed(31687, LUT_AMPL_WIDTH),
		19071 => to_signed(31686, LUT_AMPL_WIDTH),
		19072 => to_signed(31685, LUT_AMPL_WIDTH),
		19073 => to_signed(31684, LUT_AMPL_WIDTH),
		19074 => to_signed(31683, LUT_AMPL_WIDTH),
		19075 => to_signed(31683, LUT_AMPL_WIDTH),
		19076 => to_signed(31682, LUT_AMPL_WIDTH),
		19077 => to_signed(31681, LUT_AMPL_WIDTH),
		19078 => to_signed(31680, LUT_AMPL_WIDTH),
		19079 => to_signed(31679, LUT_AMPL_WIDTH),
		19080 => to_signed(31679, LUT_AMPL_WIDTH),
		19081 => to_signed(31678, LUT_AMPL_WIDTH),
		19082 => to_signed(31677, LUT_AMPL_WIDTH),
		19083 => to_signed(31676, LUT_AMPL_WIDTH),
		19084 => to_signed(31675, LUT_AMPL_WIDTH),
		19085 => to_signed(31674, LUT_AMPL_WIDTH),
		19086 => to_signed(31674, LUT_AMPL_WIDTH),
		19087 => to_signed(31673, LUT_AMPL_WIDTH),
		19088 => to_signed(31672, LUT_AMPL_WIDTH),
		19089 => to_signed(31671, LUT_AMPL_WIDTH),
		19090 => to_signed(31670, LUT_AMPL_WIDTH),
		19091 => to_signed(31670, LUT_AMPL_WIDTH),
		19092 => to_signed(31669, LUT_AMPL_WIDTH),
		19093 => to_signed(31668, LUT_AMPL_WIDTH),
		19094 => to_signed(31667, LUT_AMPL_WIDTH),
		19095 => to_signed(31666, LUT_AMPL_WIDTH),
		19096 => to_signed(31666, LUT_AMPL_WIDTH),
		19097 => to_signed(31665, LUT_AMPL_WIDTH),
		19098 => to_signed(31664, LUT_AMPL_WIDTH),
		19099 => to_signed(31663, LUT_AMPL_WIDTH),
		19100 => to_signed(31662, LUT_AMPL_WIDTH),
		19101 => to_signed(31662, LUT_AMPL_WIDTH),
		19102 => to_signed(31661, LUT_AMPL_WIDTH),
		19103 => to_signed(31660, LUT_AMPL_WIDTH),
		19104 => to_signed(31659, LUT_AMPL_WIDTH),
		19105 => to_signed(31658, LUT_AMPL_WIDTH),
		19106 => to_signed(31658, LUT_AMPL_WIDTH),
		19107 => to_signed(31657, LUT_AMPL_WIDTH),
		19108 => to_signed(31656, LUT_AMPL_WIDTH),
		19109 => to_signed(31655, LUT_AMPL_WIDTH),
		19110 => to_signed(31654, LUT_AMPL_WIDTH),
		19111 => to_signed(31653, LUT_AMPL_WIDTH),
		19112 => to_signed(31653, LUT_AMPL_WIDTH),
		19113 => to_signed(31652, LUT_AMPL_WIDTH),
		19114 => to_signed(31651, LUT_AMPL_WIDTH),
		19115 => to_signed(31650, LUT_AMPL_WIDTH),
		19116 => to_signed(31649, LUT_AMPL_WIDTH),
		19117 => to_signed(31649, LUT_AMPL_WIDTH),
		19118 => to_signed(31648, LUT_AMPL_WIDTH),
		19119 => to_signed(31647, LUT_AMPL_WIDTH),
		19120 => to_signed(31646, LUT_AMPL_WIDTH),
		19121 => to_signed(31645, LUT_AMPL_WIDTH),
		19122 => to_signed(31645, LUT_AMPL_WIDTH),
		19123 => to_signed(31644, LUT_AMPL_WIDTH),
		19124 => to_signed(31643, LUT_AMPL_WIDTH),
		19125 => to_signed(31642, LUT_AMPL_WIDTH),
		19126 => to_signed(31641, LUT_AMPL_WIDTH),
		19127 => to_signed(31640, LUT_AMPL_WIDTH),
		19128 => to_signed(31640, LUT_AMPL_WIDTH),
		19129 => to_signed(31639, LUT_AMPL_WIDTH),
		19130 => to_signed(31638, LUT_AMPL_WIDTH),
		19131 => to_signed(31637, LUT_AMPL_WIDTH),
		19132 => to_signed(31636, LUT_AMPL_WIDTH),
		19133 => to_signed(31636, LUT_AMPL_WIDTH),
		19134 => to_signed(31635, LUT_AMPL_WIDTH),
		19135 => to_signed(31634, LUT_AMPL_WIDTH),
		19136 => to_signed(31633, LUT_AMPL_WIDTH),
		19137 => to_signed(31632, LUT_AMPL_WIDTH),
		19138 => to_signed(31631, LUT_AMPL_WIDTH),
		19139 => to_signed(31631, LUT_AMPL_WIDTH),
		19140 => to_signed(31630, LUT_AMPL_WIDTH),
		19141 => to_signed(31629, LUT_AMPL_WIDTH),
		19142 => to_signed(31628, LUT_AMPL_WIDTH),
		19143 => to_signed(31627, LUT_AMPL_WIDTH),
		19144 => to_signed(31627, LUT_AMPL_WIDTH),
		19145 => to_signed(31626, LUT_AMPL_WIDTH),
		19146 => to_signed(31625, LUT_AMPL_WIDTH),
		19147 => to_signed(31624, LUT_AMPL_WIDTH),
		19148 => to_signed(31623, LUT_AMPL_WIDTH),
		19149 => to_signed(31622, LUT_AMPL_WIDTH),
		19150 => to_signed(31622, LUT_AMPL_WIDTH),
		19151 => to_signed(31621, LUT_AMPL_WIDTH),
		19152 => to_signed(31620, LUT_AMPL_WIDTH),
		19153 => to_signed(31619, LUT_AMPL_WIDTH),
		19154 => to_signed(31618, LUT_AMPL_WIDTH),
		19155 => to_signed(31617, LUT_AMPL_WIDTH),
		19156 => to_signed(31617, LUT_AMPL_WIDTH),
		19157 => to_signed(31616, LUT_AMPL_WIDTH),
		19158 => to_signed(31615, LUT_AMPL_WIDTH),
		19159 => to_signed(31614, LUT_AMPL_WIDTH),
		19160 => to_signed(31613, LUT_AMPL_WIDTH),
		19161 => to_signed(31613, LUT_AMPL_WIDTH),
		19162 => to_signed(31612, LUT_AMPL_WIDTH),
		19163 => to_signed(31611, LUT_AMPL_WIDTH),
		19164 => to_signed(31610, LUT_AMPL_WIDTH),
		19165 => to_signed(31609, LUT_AMPL_WIDTH),
		19166 => to_signed(31608, LUT_AMPL_WIDTH),
		19167 => to_signed(31608, LUT_AMPL_WIDTH),
		19168 => to_signed(31607, LUT_AMPL_WIDTH),
		19169 => to_signed(31606, LUT_AMPL_WIDTH),
		19170 => to_signed(31605, LUT_AMPL_WIDTH),
		19171 => to_signed(31604, LUT_AMPL_WIDTH),
		19172 => to_signed(31603, LUT_AMPL_WIDTH),
		19173 => to_signed(31603, LUT_AMPL_WIDTH),
		19174 => to_signed(31602, LUT_AMPL_WIDTH),
		19175 => to_signed(31601, LUT_AMPL_WIDTH),
		19176 => to_signed(31600, LUT_AMPL_WIDTH),
		19177 => to_signed(31599, LUT_AMPL_WIDTH),
		19178 => to_signed(31598, LUT_AMPL_WIDTH),
		19179 => to_signed(31598, LUT_AMPL_WIDTH),
		19180 => to_signed(31597, LUT_AMPL_WIDTH),
		19181 => to_signed(31596, LUT_AMPL_WIDTH),
		19182 => to_signed(31595, LUT_AMPL_WIDTH),
		19183 => to_signed(31594, LUT_AMPL_WIDTH),
		19184 => to_signed(31593, LUT_AMPL_WIDTH),
		19185 => to_signed(31593, LUT_AMPL_WIDTH),
		19186 => to_signed(31592, LUT_AMPL_WIDTH),
		19187 => to_signed(31591, LUT_AMPL_WIDTH),
		19188 => to_signed(31590, LUT_AMPL_WIDTH),
		19189 => to_signed(31589, LUT_AMPL_WIDTH),
		19190 => to_signed(31588, LUT_AMPL_WIDTH),
		19191 => to_signed(31588, LUT_AMPL_WIDTH),
		19192 => to_signed(31587, LUT_AMPL_WIDTH),
		19193 => to_signed(31586, LUT_AMPL_WIDTH),
		19194 => to_signed(31585, LUT_AMPL_WIDTH),
		19195 => to_signed(31584, LUT_AMPL_WIDTH),
		19196 => to_signed(31583, LUT_AMPL_WIDTH),
		19197 => to_signed(31583, LUT_AMPL_WIDTH),
		19198 => to_signed(31582, LUT_AMPL_WIDTH),
		19199 => to_signed(31581, LUT_AMPL_WIDTH),
		19200 => to_signed(31580, LUT_AMPL_WIDTH),
		19201 => to_signed(31579, LUT_AMPL_WIDTH),
		19202 => to_signed(31578, LUT_AMPL_WIDTH),
		19203 => to_signed(31578, LUT_AMPL_WIDTH),
		19204 => to_signed(31577, LUT_AMPL_WIDTH),
		19205 => to_signed(31576, LUT_AMPL_WIDTH),
		19206 => to_signed(31575, LUT_AMPL_WIDTH),
		19207 => to_signed(31574, LUT_AMPL_WIDTH),
		19208 => to_signed(31573, LUT_AMPL_WIDTH),
		19209 => to_signed(31572, LUT_AMPL_WIDTH),
		19210 => to_signed(31572, LUT_AMPL_WIDTH),
		19211 => to_signed(31571, LUT_AMPL_WIDTH),
		19212 => to_signed(31570, LUT_AMPL_WIDTH),
		19213 => to_signed(31569, LUT_AMPL_WIDTH),
		19214 => to_signed(31568, LUT_AMPL_WIDTH),
		19215 => to_signed(31567, LUT_AMPL_WIDTH),
		19216 => to_signed(31567, LUT_AMPL_WIDTH),
		19217 => to_signed(31566, LUT_AMPL_WIDTH),
		19218 => to_signed(31565, LUT_AMPL_WIDTH),
		19219 => to_signed(31564, LUT_AMPL_WIDTH),
		19220 => to_signed(31563, LUT_AMPL_WIDTH),
		19221 => to_signed(31562, LUT_AMPL_WIDTH),
		19222 => to_signed(31562, LUT_AMPL_WIDTH),
		19223 => to_signed(31561, LUT_AMPL_WIDTH),
		19224 => to_signed(31560, LUT_AMPL_WIDTH),
		19225 => to_signed(31559, LUT_AMPL_WIDTH),
		19226 => to_signed(31558, LUT_AMPL_WIDTH),
		19227 => to_signed(31557, LUT_AMPL_WIDTH),
		19228 => to_signed(31556, LUT_AMPL_WIDTH),
		19229 => to_signed(31556, LUT_AMPL_WIDTH),
		19230 => to_signed(31555, LUT_AMPL_WIDTH),
		19231 => to_signed(31554, LUT_AMPL_WIDTH),
		19232 => to_signed(31553, LUT_AMPL_WIDTH),
		19233 => to_signed(31552, LUT_AMPL_WIDTH),
		19234 => to_signed(31551, LUT_AMPL_WIDTH),
		19235 => to_signed(31551, LUT_AMPL_WIDTH),
		19236 => to_signed(31550, LUT_AMPL_WIDTH),
		19237 => to_signed(31549, LUT_AMPL_WIDTH),
		19238 => to_signed(31548, LUT_AMPL_WIDTH),
		19239 => to_signed(31547, LUT_AMPL_WIDTH),
		19240 => to_signed(31546, LUT_AMPL_WIDTH),
		19241 => to_signed(31545, LUT_AMPL_WIDTH),
		19242 => to_signed(31545, LUT_AMPL_WIDTH),
		19243 => to_signed(31544, LUT_AMPL_WIDTH),
		19244 => to_signed(31543, LUT_AMPL_WIDTH),
		19245 => to_signed(31542, LUT_AMPL_WIDTH),
		19246 => to_signed(31541, LUT_AMPL_WIDTH),
		19247 => to_signed(31540, LUT_AMPL_WIDTH),
		19248 => to_signed(31539, LUT_AMPL_WIDTH),
		19249 => to_signed(31539, LUT_AMPL_WIDTH),
		19250 => to_signed(31538, LUT_AMPL_WIDTH),
		19251 => to_signed(31537, LUT_AMPL_WIDTH),
		19252 => to_signed(31536, LUT_AMPL_WIDTH),
		19253 => to_signed(31535, LUT_AMPL_WIDTH),
		19254 => to_signed(31534, LUT_AMPL_WIDTH),
		19255 => to_signed(31534, LUT_AMPL_WIDTH),
		19256 => to_signed(31533, LUT_AMPL_WIDTH),
		19257 => to_signed(31532, LUT_AMPL_WIDTH),
		19258 => to_signed(31531, LUT_AMPL_WIDTH),
		19259 => to_signed(31530, LUT_AMPL_WIDTH),
		19260 => to_signed(31529, LUT_AMPL_WIDTH),
		19261 => to_signed(31528, LUT_AMPL_WIDTH),
		19262 => to_signed(31528, LUT_AMPL_WIDTH),
		19263 => to_signed(31527, LUT_AMPL_WIDTH),
		19264 => to_signed(31526, LUT_AMPL_WIDTH),
		19265 => to_signed(31525, LUT_AMPL_WIDTH),
		19266 => to_signed(31524, LUT_AMPL_WIDTH),
		19267 => to_signed(31523, LUT_AMPL_WIDTH),
		19268 => to_signed(31522, LUT_AMPL_WIDTH),
		19269 => to_signed(31522, LUT_AMPL_WIDTH),
		19270 => to_signed(31521, LUT_AMPL_WIDTH),
		19271 => to_signed(31520, LUT_AMPL_WIDTH),
		19272 => to_signed(31519, LUT_AMPL_WIDTH),
		19273 => to_signed(31518, LUT_AMPL_WIDTH),
		19274 => to_signed(31517, LUT_AMPL_WIDTH),
		19275 => to_signed(31516, LUT_AMPL_WIDTH),
		19276 => to_signed(31516, LUT_AMPL_WIDTH),
		19277 => to_signed(31515, LUT_AMPL_WIDTH),
		19278 => to_signed(31514, LUT_AMPL_WIDTH),
		19279 => to_signed(31513, LUT_AMPL_WIDTH),
		19280 => to_signed(31512, LUT_AMPL_WIDTH),
		19281 => to_signed(31511, LUT_AMPL_WIDTH),
		19282 => to_signed(31510, LUT_AMPL_WIDTH),
		19283 => to_signed(31510, LUT_AMPL_WIDTH),
		19284 => to_signed(31509, LUT_AMPL_WIDTH),
		19285 => to_signed(31508, LUT_AMPL_WIDTH),
		19286 => to_signed(31507, LUT_AMPL_WIDTH),
		19287 => to_signed(31506, LUT_AMPL_WIDTH),
		19288 => to_signed(31505, LUT_AMPL_WIDTH),
		19289 => to_signed(31504, LUT_AMPL_WIDTH),
		19290 => to_signed(31503, LUT_AMPL_WIDTH),
		19291 => to_signed(31503, LUT_AMPL_WIDTH),
		19292 => to_signed(31502, LUT_AMPL_WIDTH),
		19293 => to_signed(31501, LUT_AMPL_WIDTH),
		19294 => to_signed(31500, LUT_AMPL_WIDTH),
		19295 => to_signed(31499, LUT_AMPL_WIDTH),
		19296 => to_signed(31498, LUT_AMPL_WIDTH),
		19297 => to_signed(31497, LUT_AMPL_WIDTH),
		19298 => to_signed(31497, LUT_AMPL_WIDTH),
		19299 => to_signed(31496, LUT_AMPL_WIDTH),
		19300 => to_signed(31495, LUT_AMPL_WIDTH),
		19301 => to_signed(31494, LUT_AMPL_WIDTH),
		19302 => to_signed(31493, LUT_AMPL_WIDTH),
		19303 => to_signed(31492, LUT_AMPL_WIDTH),
		19304 => to_signed(31491, LUT_AMPL_WIDTH),
		19305 => to_signed(31490, LUT_AMPL_WIDTH),
		19306 => to_signed(31490, LUT_AMPL_WIDTH),
		19307 => to_signed(31489, LUT_AMPL_WIDTH),
		19308 => to_signed(31488, LUT_AMPL_WIDTH),
		19309 => to_signed(31487, LUT_AMPL_WIDTH),
		19310 => to_signed(31486, LUT_AMPL_WIDTH),
		19311 => to_signed(31485, LUT_AMPL_WIDTH),
		19312 => to_signed(31484, LUT_AMPL_WIDTH),
		19313 => to_signed(31484, LUT_AMPL_WIDTH),
		19314 => to_signed(31483, LUT_AMPL_WIDTH),
		19315 => to_signed(31482, LUT_AMPL_WIDTH),
		19316 => to_signed(31481, LUT_AMPL_WIDTH),
		19317 => to_signed(31480, LUT_AMPL_WIDTH),
		19318 => to_signed(31479, LUT_AMPL_WIDTH),
		19319 => to_signed(31478, LUT_AMPL_WIDTH),
		19320 => to_signed(31477, LUT_AMPL_WIDTH),
		19321 => to_signed(31477, LUT_AMPL_WIDTH),
		19322 => to_signed(31476, LUT_AMPL_WIDTH),
		19323 => to_signed(31475, LUT_AMPL_WIDTH),
		19324 => to_signed(31474, LUT_AMPL_WIDTH),
		19325 => to_signed(31473, LUT_AMPL_WIDTH),
		19326 => to_signed(31472, LUT_AMPL_WIDTH),
		19327 => to_signed(31471, LUT_AMPL_WIDTH),
		19328 => to_signed(31470, LUT_AMPL_WIDTH),
		19329 => to_signed(31470, LUT_AMPL_WIDTH),
		19330 => to_signed(31469, LUT_AMPL_WIDTH),
		19331 => to_signed(31468, LUT_AMPL_WIDTH),
		19332 => to_signed(31467, LUT_AMPL_WIDTH),
		19333 => to_signed(31466, LUT_AMPL_WIDTH),
		19334 => to_signed(31465, LUT_AMPL_WIDTH),
		19335 => to_signed(31464, LUT_AMPL_WIDTH),
		19336 => to_signed(31463, LUT_AMPL_WIDTH),
		19337 => to_signed(31463, LUT_AMPL_WIDTH),
		19338 => to_signed(31462, LUT_AMPL_WIDTH),
		19339 => to_signed(31461, LUT_AMPL_WIDTH),
		19340 => to_signed(31460, LUT_AMPL_WIDTH),
		19341 => to_signed(31459, LUT_AMPL_WIDTH),
		19342 => to_signed(31458, LUT_AMPL_WIDTH),
		19343 => to_signed(31457, LUT_AMPL_WIDTH),
		19344 => to_signed(31456, LUT_AMPL_WIDTH),
		19345 => to_signed(31456, LUT_AMPL_WIDTH),
		19346 => to_signed(31455, LUT_AMPL_WIDTH),
		19347 => to_signed(31454, LUT_AMPL_WIDTH),
		19348 => to_signed(31453, LUT_AMPL_WIDTH),
		19349 => to_signed(31452, LUT_AMPL_WIDTH),
		19350 => to_signed(31451, LUT_AMPL_WIDTH),
		19351 => to_signed(31450, LUT_AMPL_WIDTH),
		19352 => to_signed(31449, LUT_AMPL_WIDTH),
		19353 => to_signed(31448, LUT_AMPL_WIDTH),
		19354 => to_signed(31448, LUT_AMPL_WIDTH),
		19355 => to_signed(31447, LUT_AMPL_WIDTH),
		19356 => to_signed(31446, LUT_AMPL_WIDTH),
		19357 => to_signed(31445, LUT_AMPL_WIDTH),
		19358 => to_signed(31444, LUT_AMPL_WIDTH),
		19359 => to_signed(31443, LUT_AMPL_WIDTH),
		19360 => to_signed(31442, LUT_AMPL_WIDTH),
		19361 => to_signed(31441, LUT_AMPL_WIDTH),
		19362 => to_signed(31441, LUT_AMPL_WIDTH),
		19363 => to_signed(31440, LUT_AMPL_WIDTH),
		19364 => to_signed(31439, LUT_AMPL_WIDTH),
		19365 => to_signed(31438, LUT_AMPL_WIDTH),
		19366 => to_signed(31437, LUT_AMPL_WIDTH),
		19367 => to_signed(31436, LUT_AMPL_WIDTH),
		19368 => to_signed(31435, LUT_AMPL_WIDTH),
		19369 => to_signed(31434, LUT_AMPL_WIDTH),
		19370 => to_signed(31433, LUT_AMPL_WIDTH),
		19371 => to_signed(31433, LUT_AMPL_WIDTH),
		19372 => to_signed(31432, LUT_AMPL_WIDTH),
		19373 => to_signed(31431, LUT_AMPL_WIDTH),
		19374 => to_signed(31430, LUT_AMPL_WIDTH),
		19375 => to_signed(31429, LUT_AMPL_WIDTH),
		19376 => to_signed(31428, LUT_AMPL_WIDTH),
		19377 => to_signed(31427, LUT_AMPL_WIDTH),
		19378 => to_signed(31426, LUT_AMPL_WIDTH),
		19379 => to_signed(31425, LUT_AMPL_WIDTH),
		19380 => to_signed(31425, LUT_AMPL_WIDTH),
		19381 => to_signed(31424, LUT_AMPL_WIDTH),
		19382 => to_signed(31423, LUT_AMPL_WIDTH),
		19383 => to_signed(31422, LUT_AMPL_WIDTH),
		19384 => to_signed(31421, LUT_AMPL_WIDTH),
		19385 => to_signed(31420, LUT_AMPL_WIDTH),
		19386 => to_signed(31419, LUT_AMPL_WIDTH),
		19387 => to_signed(31418, LUT_AMPL_WIDTH),
		19388 => to_signed(31417, LUT_AMPL_WIDTH),
		19389 => to_signed(31417, LUT_AMPL_WIDTH),
		19390 => to_signed(31416, LUT_AMPL_WIDTH),
		19391 => to_signed(31415, LUT_AMPL_WIDTH),
		19392 => to_signed(31414, LUT_AMPL_WIDTH),
		19393 => to_signed(31413, LUT_AMPL_WIDTH),
		19394 => to_signed(31412, LUT_AMPL_WIDTH),
		19395 => to_signed(31411, LUT_AMPL_WIDTH),
		19396 => to_signed(31410, LUT_AMPL_WIDTH),
		19397 => to_signed(31409, LUT_AMPL_WIDTH),
		19398 => to_signed(31408, LUT_AMPL_WIDTH),
		19399 => to_signed(31408, LUT_AMPL_WIDTH),
		19400 => to_signed(31407, LUT_AMPL_WIDTH),
		19401 => to_signed(31406, LUT_AMPL_WIDTH),
		19402 => to_signed(31405, LUT_AMPL_WIDTH),
		19403 => to_signed(31404, LUT_AMPL_WIDTH),
		19404 => to_signed(31403, LUT_AMPL_WIDTH),
		19405 => to_signed(31402, LUT_AMPL_WIDTH),
		19406 => to_signed(31401, LUT_AMPL_WIDTH),
		19407 => to_signed(31400, LUT_AMPL_WIDTH),
		19408 => to_signed(31400, LUT_AMPL_WIDTH),
		19409 => to_signed(31399, LUT_AMPL_WIDTH),
		19410 => to_signed(31398, LUT_AMPL_WIDTH),
		19411 => to_signed(31397, LUT_AMPL_WIDTH),
		19412 => to_signed(31396, LUT_AMPL_WIDTH),
		19413 => to_signed(31395, LUT_AMPL_WIDTH),
		19414 => to_signed(31394, LUT_AMPL_WIDTH),
		19415 => to_signed(31393, LUT_AMPL_WIDTH),
		19416 => to_signed(31392, LUT_AMPL_WIDTH),
		19417 => to_signed(31391, LUT_AMPL_WIDTH),
		19418 => to_signed(31391, LUT_AMPL_WIDTH),
		19419 => to_signed(31390, LUT_AMPL_WIDTH),
		19420 => to_signed(31389, LUT_AMPL_WIDTH),
		19421 => to_signed(31388, LUT_AMPL_WIDTH),
		19422 => to_signed(31387, LUT_AMPL_WIDTH),
		19423 => to_signed(31386, LUT_AMPL_WIDTH),
		19424 => to_signed(31385, LUT_AMPL_WIDTH),
		19425 => to_signed(31384, LUT_AMPL_WIDTH),
		19426 => to_signed(31383, LUT_AMPL_WIDTH),
		19427 => to_signed(31382, LUT_AMPL_WIDTH),
		19428 => to_signed(31381, LUT_AMPL_WIDTH),
		19429 => to_signed(31381, LUT_AMPL_WIDTH),
		19430 => to_signed(31380, LUT_AMPL_WIDTH),
		19431 => to_signed(31379, LUT_AMPL_WIDTH),
		19432 => to_signed(31378, LUT_AMPL_WIDTH),
		19433 => to_signed(31377, LUT_AMPL_WIDTH),
		19434 => to_signed(31376, LUT_AMPL_WIDTH),
		19435 => to_signed(31375, LUT_AMPL_WIDTH),
		19436 => to_signed(31374, LUT_AMPL_WIDTH),
		19437 => to_signed(31373, LUT_AMPL_WIDTH),
		19438 => to_signed(31372, LUT_AMPL_WIDTH),
		19439 => to_signed(31372, LUT_AMPL_WIDTH),
		19440 => to_signed(31371, LUT_AMPL_WIDTH),
		19441 => to_signed(31370, LUT_AMPL_WIDTH),
		19442 => to_signed(31369, LUT_AMPL_WIDTH),
		19443 => to_signed(31368, LUT_AMPL_WIDTH),
		19444 => to_signed(31367, LUT_AMPL_WIDTH),
		19445 => to_signed(31366, LUT_AMPL_WIDTH),
		19446 => to_signed(31365, LUT_AMPL_WIDTH),
		19447 => to_signed(31364, LUT_AMPL_WIDTH),
		19448 => to_signed(31363, LUT_AMPL_WIDTH),
		19449 => to_signed(31362, LUT_AMPL_WIDTH),
		19450 => to_signed(31362, LUT_AMPL_WIDTH),
		19451 => to_signed(31361, LUT_AMPL_WIDTH),
		19452 => to_signed(31360, LUT_AMPL_WIDTH),
		19453 => to_signed(31359, LUT_AMPL_WIDTH),
		19454 => to_signed(31358, LUT_AMPL_WIDTH),
		19455 => to_signed(31357, LUT_AMPL_WIDTH),
		19456 => to_signed(31356, LUT_AMPL_WIDTH),
		19457 => to_signed(31355, LUT_AMPL_WIDTH),
		19458 => to_signed(31354, LUT_AMPL_WIDTH),
		19459 => to_signed(31353, LUT_AMPL_WIDTH),
		19460 => to_signed(31352, LUT_AMPL_WIDTH),
		19461 => to_signed(31352, LUT_AMPL_WIDTH),
		19462 => to_signed(31351, LUT_AMPL_WIDTH),
		19463 => to_signed(31350, LUT_AMPL_WIDTH),
		19464 => to_signed(31349, LUT_AMPL_WIDTH),
		19465 => to_signed(31348, LUT_AMPL_WIDTH),
		19466 => to_signed(31347, LUT_AMPL_WIDTH),
		19467 => to_signed(31346, LUT_AMPL_WIDTH),
		19468 => to_signed(31345, LUT_AMPL_WIDTH),
		19469 => to_signed(31344, LUT_AMPL_WIDTH),
		19470 => to_signed(31343, LUT_AMPL_WIDTH),
		19471 => to_signed(31342, LUT_AMPL_WIDTH),
		19472 => to_signed(31341, LUT_AMPL_WIDTH),
		19473 => to_signed(31341, LUT_AMPL_WIDTH),
		19474 => to_signed(31340, LUT_AMPL_WIDTH),
		19475 => to_signed(31339, LUT_AMPL_WIDTH),
		19476 => to_signed(31338, LUT_AMPL_WIDTH),
		19477 => to_signed(31337, LUT_AMPL_WIDTH),
		19478 => to_signed(31336, LUT_AMPL_WIDTH),
		19479 => to_signed(31335, LUT_AMPL_WIDTH),
		19480 => to_signed(31334, LUT_AMPL_WIDTH),
		19481 => to_signed(31333, LUT_AMPL_WIDTH),
		19482 => to_signed(31332, LUT_AMPL_WIDTH),
		19483 => to_signed(31331, LUT_AMPL_WIDTH),
		19484 => to_signed(31330, LUT_AMPL_WIDTH),
		19485 => to_signed(31329, LUT_AMPL_WIDTH),
		19486 => to_signed(31329, LUT_AMPL_WIDTH),
		19487 => to_signed(31328, LUT_AMPL_WIDTH),
		19488 => to_signed(31327, LUT_AMPL_WIDTH),
		19489 => to_signed(31326, LUT_AMPL_WIDTH),
		19490 => to_signed(31325, LUT_AMPL_WIDTH),
		19491 => to_signed(31324, LUT_AMPL_WIDTH),
		19492 => to_signed(31323, LUT_AMPL_WIDTH),
		19493 => to_signed(31322, LUT_AMPL_WIDTH),
		19494 => to_signed(31321, LUT_AMPL_WIDTH),
		19495 => to_signed(31320, LUT_AMPL_WIDTH),
		19496 => to_signed(31319, LUT_AMPL_WIDTH),
		19497 => to_signed(31318, LUT_AMPL_WIDTH),
		19498 => to_signed(31318, LUT_AMPL_WIDTH),
		19499 => to_signed(31317, LUT_AMPL_WIDTH),
		19500 => to_signed(31316, LUT_AMPL_WIDTH),
		19501 => to_signed(31315, LUT_AMPL_WIDTH),
		19502 => to_signed(31314, LUT_AMPL_WIDTH),
		19503 => to_signed(31313, LUT_AMPL_WIDTH),
		19504 => to_signed(31312, LUT_AMPL_WIDTH),
		19505 => to_signed(31311, LUT_AMPL_WIDTH),
		19506 => to_signed(31310, LUT_AMPL_WIDTH),
		19507 => to_signed(31309, LUT_AMPL_WIDTH),
		19508 => to_signed(31308, LUT_AMPL_WIDTH),
		19509 => to_signed(31307, LUT_AMPL_WIDTH),
		19510 => to_signed(31306, LUT_AMPL_WIDTH),
		19511 => to_signed(31305, LUT_AMPL_WIDTH),
		19512 => to_signed(31305, LUT_AMPL_WIDTH),
		19513 => to_signed(31304, LUT_AMPL_WIDTH),
		19514 => to_signed(31303, LUT_AMPL_WIDTH),
		19515 => to_signed(31302, LUT_AMPL_WIDTH),
		19516 => to_signed(31301, LUT_AMPL_WIDTH),
		19517 => to_signed(31300, LUT_AMPL_WIDTH),
		19518 => to_signed(31299, LUT_AMPL_WIDTH),
		19519 => to_signed(31298, LUT_AMPL_WIDTH),
		19520 => to_signed(31297, LUT_AMPL_WIDTH),
		19521 => to_signed(31296, LUT_AMPL_WIDTH),
		19522 => to_signed(31295, LUT_AMPL_WIDTH),
		19523 => to_signed(31294, LUT_AMPL_WIDTH),
		19524 => to_signed(31293, LUT_AMPL_WIDTH),
		19525 => to_signed(31292, LUT_AMPL_WIDTH),
		19526 => to_signed(31292, LUT_AMPL_WIDTH),
		19527 => to_signed(31291, LUT_AMPL_WIDTH),
		19528 => to_signed(31290, LUT_AMPL_WIDTH),
		19529 => to_signed(31289, LUT_AMPL_WIDTH),
		19530 => to_signed(31288, LUT_AMPL_WIDTH),
		19531 => to_signed(31287, LUT_AMPL_WIDTH),
		19532 => to_signed(31286, LUT_AMPL_WIDTH),
		19533 => to_signed(31285, LUT_AMPL_WIDTH),
		19534 => to_signed(31284, LUT_AMPL_WIDTH),
		19535 => to_signed(31283, LUT_AMPL_WIDTH),
		19536 => to_signed(31282, LUT_AMPL_WIDTH),
		19537 => to_signed(31281, LUT_AMPL_WIDTH),
		19538 => to_signed(31280, LUT_AMPL_WIDTH),
		19539 => to_signed(31279, LUT_AMPL_WIDTH),
		19540 => to_signed(31278, LUT_AMPL_WIDTH),
		19541 => to_signed(31278, LUT_AMPL_WIDTH),
		19542 => to_signed(31277, LUT_AMPL_WIDTH),
		19543 => to_signed(31276, LUT_AMPL_WIDTH),
		19544 => to_signed(31275, LUT_AMPL_WIDTH),
		19545 => to_signed(31274, LUT_AMPL_WIDTH),
		19546 => to_signed(31273, LUT_AMPL_WIDTH),
		19547 => to_signed(31272, LUT_AMPL_WIDTH),
		19548 => to_signed(31271, LUT_AMPL_WIDTH),
		19549 => to_signed(31270, LUT_AMPL_WIDTH),
		19550 => to_signed(31269, LUT_AMPL_WIDTH),
		19551 => to_signed(31268, LUT_AMPL_WIDTH),
		19552 => to_signed(31267, LUT_AMPL_WIDTH),
		19553 => to_signed(31266, LUT_AMPL_WIDTH),
		19554 => to_signed(31265, LUT_AMPL_WIDTH),
		19555 => to_signed(31264, LUT_AMPL_WIDTH),
		19556 => to_signed(31263, LUT_AMPL_WIDTH),
		19557 => to_signed(31262, LUT_AMPL_WIDTH),
		19558 => to_signed(31262, LUT_AMPL_WIDTH),
		19559 => to_signed(31261, LUT_AMPL_WIDTH),
		19560 => to_signed(31260, LUT_AMPL_WIDTH),
		19561 => to_signed(31259, LUT_AMPL_WIDTH),
		19562 => to_signed(31258, LUT_AMPL_WIDTH),
		19563 => to_signed(31257, LUT_AMPL_WIDTH),
		19564 => to_signed(31256, LUT_AMPL_WIDTH),
		19565 => to_signed(31255, LUT_AMPL_WIDTH),
		19566 => to_signed(31254, LUT_AMPL_WIDTH),
		19567 => to_signed(31253, LUT_AMPL_WIDTH),
		19568 => to_signed(31252, LUT_AMPL_WIDTH),
		19569 => to_signed(31251, LUT_AMPL_WIDTH),
		19570 => to_signed(31250, LUT_AMPL_WIDTH),
		19571 => to_signed(31249, LUT_AMPL_WIDTH),
		19572 => to_signed(31248, LUT_AMPL_WIDTH),
		19573 => to_signed(31247, LUT_AMPL_WIDTH),
		19574 => to_signed(31246, LUT_AMPL_WIDTH),
		19575 => to_signed(31246, LUT_AMPL_WIDTH),
		19576 => to_signed(31245, LUT_AMPL_WIDTH),
		19577 => to_signed(31244, LUT_AMPL_WIDTH),
		19578 => to_signed(31243, LUT_AMPL_WIDTH),
		19579 => to_signed(31242, LUT_AMPL_WIDTH),
		19580 => to_signed(31241, LUT_AMPL_WIDTH),
		19581 => to_signed(31240, LUT_AMPL_WIDTH),
		19582 => to_signed(31239, LUT_AMPL_WIDTH),
		19583 => to_signed(31238, LUT_AMPL_WIDTH),
		19584 => to_signed(31237, LUT_AMPL_WIDTH),
		19585 => to_signed(31236, LUT_AMPL_WIDTH),
		19586 => to_signed(31235, LUT_AMPL_WIDTH),
		19587 => to_signed(31234, LUT_AMPL_WIDTH),
		19588 => to_signed(31233, LUT_AMPL_WIDTH),
		19589 => to_signed(31232, LUT_AMPL_WIDTH),
		19590 => to_signed(31231, LUT_AMPL_WIDTH),
		19591 => to_signed(31230, LUT_AMPL_WIDTH),
		19592 => to_signed(31229, LUT_AMPL_WIDTH),
		19593 => to_signed(31228, LUT_AMPL_WIDTH),
		19594 => to_signed(31227, LUT_AMPL_WIDTH),
		19595 => to_signed(31227, LUT_AMPL_WIDTH),
		19596 => to_signed(31226, LUT_AMPL_WIDTH),
		19597 => to_signed(31225, LUT_AMPL_WIDTH),
		19598 => to_signed(31224, LUT_AMPL_WIDTH),
		19599 => to_signed(31223, LUT_AMPL_WIDTH),
		19600 => to_signed(31222, LUT_AMPL_WIDTH),
		19601 => to_signed(31221, LUT_AMPL_WIDTH),
		19602 => to_signed(31220, LUT_AMPL_WIDTH),
		19603 => to_signed(31219, LUT_AMPL_WIDTH),
		19604 => to_signed(31218, LUT_AMPL_WIDTH),
		19605 => to_signed(31217, LUT_AMPL_WIDTH),
		19606 => to_signed(31216, LUT_AMPL_WIDTH),
		19607 => to_signed(31215, LUT_AMPL_WIDTH),
		19608 => to_signed(31214, LUT_AMPL_WIDTH),
		19609 => to_signed(31213, LUT_AMPL_WIDTH),
		19610 => to_signed(31212, LUT_AMPL_WIDTH),
		19611 => to_signed(31211, LUT_AMPL_WIDTH),
		19612 => to_signed(31210, LUT_AMPL_WIDTH),
		19613 => to_signed(31209, LUT_AMPL_WIDTH),
		19614 => to_signed(31208, LUT_AMPL_WIDTH),
		19615 => to_signed(31207, LUT_AMPL_WIDTH),
		19616 => to_signed(31206, LUT_AMPL_WIDTH),
		19617 => to_signed(31206, LUT_AMPL_WIDTH),
		19618 => to_signed(31205, LUT_AMPL_WIDTH),
		19619 => to_signed(31204, LUT_AMPL_WIDTH),
		19620 => to_signed(31203, LUT_AMPL_WIDTH),
		19621 => to_signed(31202, LUT_AMPL_WIDTH),
		19622 => to_signed(31201, LUT_AMPL_WIDTH),
		19623 => to_signed(31200, LUT_AMPL_WIDTH),
		19624 => to_signed(31199, LUT_AMPL_WIDTH),
		19625 => to_signed(31198, LUT_AMPL_WIDTH),
		19626 => to_signed(31197, LUT_AMPL_WIDTH),
		19627 => to_signed(31196, LUT_AMPL_WIDTH),
		19628 => to_signed(31195, LUT_AMPL_WIDTH),
		19629 => to_signed(31194, LUT_AMPL_WIDTH),
		19630 => to_signed(31193, LUT_AMPL_WIDTH),
		19631 => to_signed(31192, LUT_AMPL_WIDTH),
		19632 => to_signed(31191, LUT_AMPL_WIDTH),
		19633 => to_signed(31190, LUT_AMPL_WIDTH),
		19634 => to_signed(31189, LUT_AMPL_WIDTH),
		19635 => to_signed(31188, LUT_AMPL_WIDTH),
		19636 => to_signed(31187, LUT_AMPL_WIDTH),
		19637 => to_signed(31186, LUT_AMPL_WIDTH),
		19638 => to_signed(31185, LUT_AMPL_WIDTH),
		19639 => to_signed(31184, LUT_AMPL_WIDTH),
		19640 => to_signed(31183, LUT_AMPL_WIDTH),
		19641 => to_signed(31182, LUT_AMPL_WIDTH),
		19642 => to_signed(31181, LUT_AMPL_WIDTH),
		19643 => to_signed(31181, LUT_AMPL_WIDTH),
		19644 => to_signed(31180, LUT_AMPL_WIDTH),
		19645 => to_signed(31179, LUT_AMPL_WIDTH),
		19646 => to_signed(31178, LUT_AMPL_WIDTH),
		19647 => to_signed(31177, LUT_AMPL_WIDTH),
		19648 => to_signed(31176, LUT_AMPL_WIDTH),
		19649 => to_signed(31175, LUT_AMPL_WIDTH),
		19650 => to_signed(31174, LUT_AMPL_WIDTH),
		19651 => to_signed(31173, LUT_AMPL_WIDTH),
		19652 => to_signed(31172, LUT_AMPL_WIDTH),
		19653 => to_signed(31171, LUT_AMPL_WIDTH),
		19654 => to_signed(31170, LUT_AMPL_WIDTH),
		19655 => to_signed(31169, LUT_AMPL_WIDTH),
		19656 => to_signed(31168, LUT_AMPL_WIDTH),
		19657 => to_signed(31167, LUT_AMPL_WIDTH),
		19658 => to_signed(31166, LUT_AMPL_WIDTH),
		19659 => to_signed(31165, LUT_AMPL_WIDTH),
		19660 => to_signed(31164, LUT_AMPL_WIDTH),
		19661 => to_signed(31163, LUT_AMPL_WIDTH),
		19662 => to_signed(31162, LUT_AMPL_WIDTH),
		19663 => to_signed(31161, LUT_AMPL_WIDTH),
		19664 => to_signed(31160, LUT_AMPL_WIDTH),
		19665 => to_signed(31159, LUT_AMPL_WIDTH),
		19666 => to_signed(31158, LUT_AMPL_WIDTH),
		19667 => to_signed(31157, LUT_AMPL_WIDTH),
		19668 => to_signed(31156, LUT_AMPL_WIDTH),
		19669 => to_signed(31155, LUT_AMPL_WIDTH),
		19670 => to_signed(31154, LUT_AMPL_WIDTH),
		19671 => to_signed(31153, LUT_AMPL_WIDTH),
		19672 => to_signed(31152, LUT_AMPL_WIDTH),
		19673 => to_signed(31151, LUT_AMPL_WIDTH),
		19674 => to_signed(31150, LUT_AMPL_WIDTH),
		19675 => to_signed(31149, LUT_AMPL_WIDTH),
		19676 => to_signed(31148, LUT_AMPL_WIDTH),
		19677 => to_signed(31148, LUT_AMPL_WIDTH),
		19678 => to_signed(31147, LUT_AMPL_WIDTH),
		19679 => to_signed(31146, LUT_AMPL_WIDTH),
		19680 => to_signed(31145, LUT_AMPL_WIDTH),
		19681 => to_signed(31144, LUT_AMPL_WIDTH),
		19682 => to_signed(31143, LUT_AMPL_WIDTH),
		19683 => to_signed(31142, LUT_AMPL_WIDTH),
		19684 => to_signed(31141, LUT_AMPL_WIDTH),
		19685 => to_signed(31140, LUT_AMPL_WIDTH),
		19686 => to_signed(31139, LUT_AMPL_WIDTH),
		19687 => to_signed(31138, LUT_AMPL_WIDTH),
		19688 => to_signed(31137, LUT_AMPL_WIDTH),
		19689 => to_signed(31136, LUT_AMPL_WIDTH),
		19690 => to_signed(31135, LUT_AMPL_WIDTH),
		19691 => to_signed(31134, LUT_AMPL_WIDTH),
		19692 => to_signed(31133, LUT_AMPL_WIDTH),
		19693 => to_signed(31132, LUT_AMPL_WIDTH),
		19694 => to_signed(31131, LUT_AMPL_WIDTH),
		19695 => to_signed(31130, LUT_AMPL_WIDTH),
		19696 => to_signed(31129, LUT_AMPL_WIDTH),
		19697 => to_signed(31128, LUT_AMPL_WIDTH),
		19698 => to_signed(31127, LUT_AMPL_WIDTH),
		19699 => to_signed(31126, LUT_AMPL_WIDTH),
		19700 => to_signed(31125, LUT_AMPL_WIDTH),
		19701 => to_signed(31124, LUT_AMPL_WIDTH),
		19702 => to_signed(31123, LUT_AMPL_WIDTH),
		19703 => to_signed(31122, LUT_AMPL_WIDTH),
		19704 => to_signed(31121, LUT_AMPL_WIDTH),
		19705 => to_signed(31120, LUT_AMPL_WIDTH),
		19706 => to_signed(31119, LUT_AMPL_WIDTH),
		19707 => to_signed(31118, LUT_AMPL_WIDTH),
		19708 => to_signed(31117, LUT_AMPL_WIDTH),
		19709 => to_signed(31116, LUT_AMPL_WIDTH),
		19710 => to_signed(31115, LUT_AMPL_WIDTH),
		19711 => to_signed(31114, LUT_AMPL_WIDTH),
		19712 => to_signed(31113, LUT_AMPL_WIDTH),
		19713 => to_signed(31112, LUT_AMPL_WIDTH),
		19714 => to_signed(31111, LUT_AMPL_WIDTH),
		19715 => to_signed(31110, LUT_AMPL_WIDTH),
		19716 => to_signed(31109, LUT_AMPL_WIDTH),
		19717 => to_signed(31108, LUT_AMPL_WIDTH),
		19718 => to_signed(31107, LUT_AMPL_WIDTH),
		19719 => to_signed(31106, LUT_AMPL_WIDTH),
		19720 => to_signed(31105, LUT_AMPL_WIDTH),
		19721 => to_signed(31104, LUT_AMPL_WIDTH),
		19722 => to_signed(31103, LUT_AMPL_WIDTH),
		19723 => to_signed(31102, LUT_AMPL_WIDTH),
		19724 => to_signed(31101, LUT_AMPL_WIDTH),
		19725 => to_signed(31100, LUT_AMPL_WIDTH),
		19726 => to_signed(31099, LUT_AMPL_WIDTH),
		19727 => to_signed(31098, LUT_AMPL_WIDTH),
		19728 => to_signed(31097, LUT_AMPL_WIDTH),
		19729 => to_signed(31096, LUT_AMPL_WIDTH),
		19730 => to_signed(31095, LUT_AMPL_WIDTH),
		19731 => to_signed(31094, LUT_AMPL_WIDTH),
		19732 => to_signed(31093, LUT_AMPL_WIDTH),
		19733 => to_signed(31092, LUT_AMPL_WIDTH),
		19734 => to_signed(31091, LUT_AMPL_WIDTH),
		19735 => to_signed(31090, LUT_AMPL_WIDTH),
		19736 => to_signed(31089, LUT_AMPL_WIDTH),
		19737 => to_signed(31088, LUT_AMPL_WIDTH),
		19738 => to_signed(31087, LUT_AMPL_WIDTH),
		19739 => to_signed(31086, LUT_AMPL_WIDTH),
		19740 => to_signed(31085, LUT_AMPL_WIDTH),
		19741 => to_signed(31084, LUT_AMPL_WIDTH),
		19742 => to_signed(31083, LUT_AMPL_WIDTH),
		19743 => to_signed(31083, LUT_AMPL_WIDTH),
		19744 => to_signed(31082, LUT_AMPL_WIDTH),
		19745 => to_signed(31081, LUT_AMPL_WIDTH),
		19746 => to_signed(31080, LUT_AMPL_WIDTH),
		19747 => to_signed(31079, LUT_AMPL_WIDTH),
		19748 => to_signed(31078, LUT_AMPL_WIDTH),
		19749 => to_signed(31077, LUT_AMPL_WIDTH),
		19750 => to_signed(31076, LUT_AMPL_WIDTH),
		19751 => to_signed(31075, LUT_AMPL_WIDTH),
		19752 => to_signed(31074, LUT_AMPL_WIDTH),
		19753 => to_signed(31073, LUT_AMPL_WIDTH),
		19754 => to_signed(31072, LUT_AMPL_WIDTH),
		19755 => to_signed(31071, LUT_AMPL_WIDTH),
		19756 => to_signed(31070, LUT_AMPL_WIDTH),
		19757 => to_signed(31069, LUT_AMPL_WIDTH),
		19758 => to_signed(31068, LUT_AMPL_WIDTH),
		19759 => to_signed(31067, LUT_AMPL_WIDTH),
		19760 => to_signed(31066, LUT_AMPL_WIDTH),
		19761 => to_signed(31065, LUT_AMPL_WIDTH),
		19762 => to_signed(31064, LUT_AMPL_WIDTH),
		19763 => to_signed(31063, LUT_AMPL_WIDTH),
		19764 => to_signed(31062, LUT_AMPL_WIDTH),
		19765 => to_signed(31061, LUT_AMPL_WIDTH),
		19766 => to_signed(31060, LUT_AMPL_WIDTH),
		19767 => to_signed(31059, LUT_AMPL_WIDTH),
		19768 => to_signed(31058, LUT_AMPL_WIDTH),
		19769 => to_signed(31057, LUT_AMPL_WIDTH),
		19770 => to_signed(31056, LUT_AMPL_WIDTH),
		19771 => to_signed(31055, LUT_AMPL_WIDTH),
		19772 => to_signed(31054, LUT_AMPL_WIDTH),
		19773 => to_signed(31053, LUT_AMPL_WIDTH),
		19774 => to_signed(31052, LUT_AMPL_WIDTH),
		19775 => to_signed(31051, LUT_AMPL_WIDTH),
		19776 => to_signed(31050, LUT_AMPL_WIDTH),
		19777 => to_signed(31049, LUT_AMPL_WIDTH),
		19778 => to_signed(31048, LUT_AMPL_WIDTH),
		19779 => to_signed(31047, LUT_AMPL_WIDTH),
		19780 => to_signed(31046, LUT_AMPL_WIDTH),
		19781 => to_signed(31045, LUT_AMPL_WIDTH),
		19782 => to_signed(31044, LUT_AMPL_WIDTH),
		19783 => to_signed(31043, LUT_AMPL_WIDTH),
		19784 => to_signed(31041, LUT_AMPL_WIDTH),
		19785 => to_signed(31040, LUT_AMPL_WIDTH),
		19786 => to_signed(31039, LUT_AMPL_WIDTH),
		19787 => to_signed(31038, LUT_AMPL_WIDTH),
		19788 => to_signed(31037, LUT_AMPL_WIDTH),
		19789 => to_signed(31036, LUT_AMPL_WIDTH),
		19790 => to_signed(31035, LUT_AMPL_WIDTH),
		19791 => to_signed(31034, LUT_AMPL_WIDTH),
		19792 => to_signed(31033, LUT_AMPL_WIDTH),
		19793 => to_signed(31032, LUT_AMPL_WIDTH),
		19794 => to_signed(31031, LUT_AMPL_WIDTH),
		19795 => to_signed(31030, LUT_AMPL_WIDTH),
		19796 => to_signed(31029, LUT_AMPL_WIDTH),
		19797 => to_signed(31028, LUT_AMPL_WIDTH),
		19798 => to_signed(31027, LUT_AMPL_WIDTH),
		19799 => to_signed(31026, LUT_AMPL_WIDTH),
		19800 => to_signed(31025, LUT_AMPL_WIDTH),
		19801 => to_signed(31024, LUT_AMPL_WIDTH),
		19802 => to_signed(31023, LUT_AMPL_WIDTH),
		19803 => to_signed(31022, LUT_AMPL_WIDTH),
		19804 => to_signed(31021, LUT_AMPL_WIDTH),
		19805 => to_signed(31020, LUT_AMPL_WIDTH),
		19806 => to_signed(31019, LUT_AMPL_WIDTH),
		19807 => to_signed(31018, LUT_AMPL_WIDTH),
		19808 => to_signed(31017, LUT_AMPL_WIDTH),
		19809 => to_signed(31016, LUT_AMPL_WIDTH),
		19810 => to_signed(31015, LUT_AMPL_WIDTH),
		19811 => to_signed(31014, LUT_AMPL_WIDTH),
		19812 => to_signed(31013, LUT_AMPL_WIDTH),
		19813 => to_signed(31012, LUT_AMPL_WIDTH),
		19814 => to_signed(31011, LUT_AMPL_WIDTH),
		19815 => to_signed(31010, LUT_AMPL_WIDTH),
		19816 => to_signed(31009, LUT_AMPL_WIDTH),
		19817 => to_signed(31008, LUT_AMPL_WIDTH),
		19818 => to_signed(31007, LUT_AMPL_WIDTH),
		19819 => to_signed(31006, LUT_AMPL_WIDTH),
		19820 => to_signed(31005, LUT_AMPL_WIDTH),
		19821 => to_signed(31004, LUT_AMPL_WIDTH),
		19822 => to_signed(31003, LUT_AMPL_WIDTH),
		19823 => to_signed(31002, LUT_AMPL_WIDTH),
		19824 => to_signed(31001, LUT_AMPL_WIDTH),
		19825 => to_signed(31000, LUT_AMPL_WIDTH),
		19826 => to_signed(30999, LUT_AMPL_WIDTH),
		19827 => to_signed(30998, LUT_AMPL_WIDTH),
		19828 => to_signed(30997, LUT_AMPL_WIDTH),
		19829 => to_signed(30996, LUT_AMPL_WIDTH),
		19830 => to_signed(30995, LUT_AMPL_WIDTH),
		19831 => to_signed(30994, LUT_AMPL_WIDTH),
		19832 => to_signed(30993, LUT_AMPL_WIDTH),
		19833 => to_signed(30992, LUT_AMPL_WIDTH),
		19834 => to_signed(30991, LUT_AMPL_WIDTH),
		19835 => to_signed(30990, LUT_AMPL_WIDTH),
		19836 => to_signed(30989, LUT_AMPL_WIDTH),
		19837 => to_signed(30988, LUT_AMPL_WIDTH),
		19838 => to_signed(30987, LUT_AMPL_WIDTH),
		19839 => to_signed(30986, LUT_AMPL_WIDTH),
		19840 => to_signed(30985, LUT_AMPL_WIDTH),
		19841 => to_signed(30984, LUT_AMPL_WIDTH),
		19842 => to_signed(30983, LUT_AMPL_WIDTH),
		19843 => to_signed(30982, LUT_AMPL_WIDTH),
		19844 => to_signed(30981, LUT_AMPL_WIDTH),
		19845 => to_signed(30980, LUT_AMPL_WIDTH),
		19846 => to_signed(30979, LUT_AMPL_WIDTH),
		19847 => to_signed(30978, LUT_AMPL_WIDTH),
		19848 => to_signed(30977, LUT_AMPL_WIDTH),
		19849 => to_signed(30976, LUT_AMPL_WIDTH),
		19850 => to_signed(30974, LUT_AMPL_WIDTH),
		19851 => to_signed(30973, LUT_AMPL_WIDTH),
		19852 => to_signed(30972, LUT_AMPL_WIDTH),
		19853 => to_signed(30971, LUT_AMPL_WIDTH),
		19854 => to_signed(30970, LUT_AMPL_WIDTH),
		19855 => to_signed(30969, LUT_AMPL_WIDTH),
		19856 => to_signed(30968, LUT_AMPL_WIDTH),
		19857 => to_signed(30967, LUT_AMPL_WIDTH),
		19858 => to_signed(30966, LUT_AMPL_WIDTH),
		19859 => to_signed(30965, LUT_AMPL_WIDTH),
		19860 => to_signed(30964, LUT_AMPL_WIDTH),
		19861 => to_signed(30963, LUT_AMPL_WIDTH),
		19862 => to_signed(30962, LUT_AMPL_WIDTH),
		19863 => to_signed(30961, LUT_AMPL_WIDTH),
		19864 => to_signed(30960, LUT_AMPL_WIDTH),
		19865 => to_signed(30959, LUT_AMPL_WIDTH),
		19866 => to_signed(30958, LUT_AMPL_WIDTH),
		19867 => to_signed(30957, LUT_AMPL_WIDTH),
		19868 => to_signed(30956, LUT_AMPL_WIDTH),
		19869 => to_signed(30955, LUT_AMPL_WIDTH),
		19870 => to_signed(30954, LUT_AMPL_WIDTH),
		19871 => to_signed(30953, LUT_AMPL_WIDTH),
		19872 => to_signed(30952, LUT_AMPL_WIDTH),
		19873 => to_signed(30951, LUT_AMPL_WIDTH),
		19874 => to_signed(30950, LUT_AMPL_WIDTH),
		19875 => to_signed(30949, LUT_AMPL_WIDTH),
		19876 => to_signed(30948, LUT_AMPL_WIDTH),
		19877 => to_signed(30947, LUT_AMPL_WIDTH),
		19878 => to_signed(30946, LUT_AMPL_WIDTH),
		19879 => to_signed(30945, LUT_AMPL_WIDTH),
		19880 => to_signed(30944, LUT_AMPL_WIDTH),
		19881 => to_signed(30943, LUT_AMPL_WIDTH),
		19882 => to_signed(30942, LUT_AMPL_WIDTH),
		19883 => to_signed(30941, LUT_AMPL_WIDTH),
		19884 => to_signed(30939, LUT_AMPL_WIDTH),
		19885 => to_signed(30938, LUT_AMPL_WIDTH),
		19886 => to_signed(30937, LUT_AMPL_WIDTH),
		19887 => to_signed(30936, LUT_AMPL_WIDTH),
		19888 => to_signed(30935, LUT_AMPL_WIDTH),
		19889 => to_signed(30934, LUT_AMPL_WIDTH),
		19890 => to_signed(30933, LUT_AMPL_WIDTH),
		19891 => to_signed(30932, LUT_AMPL_WIDTH),
		19892 => to_signed(30931, LUT_AMPL_WIDTH),
		19893 => to_signed(30930, LUT_AMPL_WIDTH),
		19894 => to_signed(30929, LUT_AMPL_WIDTH),
		19895 => to_signed(30928, LUT_AMPL_WIDTH),
		19896 => to_signed(30927, LUT_AMPL_WIDTH),
		19897 => to_signed(30926, LUT_AMPL_WIDTH),
		19898 => to_signed(30925, LUT_AMPL_WIDTH),
		19899 => to_signed(30924, LUT_AMPL_WIDTH),
		19900 => to_signed(30923, LUT_AMPL_WIDTH),
		19901 => to_signed(30922, LUT_AMPL_WIDTH),
		19902 => to_signed(30921, LUT_AMPL_WIDTH),
		19903 => to_signed(30920, LUT_AMPL_WIDTH),
		19904 => to_signed(30919, LUT_AMPL_WIDTH),
		19905 => to_signed(30918, LUT_AMPL_WIDTH),
		19906 => to_signed(30917, LUT_AMPL_WIDTH),
		19907 => to_signed(30916, LUT_AMPL_WIDTH),
		19908 => to_signed(30915, LUT_AMPL_WIDTH),
		19909 => to_signed(30914, LUT_AMPL_WIDTH),
		19910 => to_signed(30912, LUT_AMPL_WIDTH),
		19911 => to_signed(30911, LUT_AMPL_WIDTH),
		19912 => to_signed(30910, LUT_AMPL_WIDTH),
		19913 => to_signed(30909, LUT_AMPL_WIDTH),
		19914 => to_signed(30908, LUT_AMPL_WIDTH),
		19915 => to_signed(30907, LUT_AMPL_WIDTH),
		19916 => to_signed(30906, LUT_AMPL_WIDTH),
		19917 => to_signed(30905, LUT_AMPL_WIDTH),
		19918 => to_signed(30904, LUT_AMPL_WIDTH),
		19919 => to_signed(30903, LUT_AMPL_WIDTH),
		19920 => to_signed(30902, LUT_AMPL_WIDTH),
		19921 => to_signed(30901, LUT_AMPL_WIDTH),
		19922 => to_signed(30900, LUT_AMPL_WIDTH),
		19923 => to_signed(30899, LUT_AMPL_WIDTH),
		19924 => to_signed(30898, LUT_AMPL_WIDTH),
		19925 => to_signed(30897, LUT_AMPL_WIDTH),
		19926 => to_signed(30896, LUT_AMPL_WIDTH),
		19927 => to_signed(30895, LUT_AMPL_WIDTH),
		19928 => to_signed(30894, LUT_AMPL_WIDTH),
		19929 => to_signed(30893, LUT_AMPL_WIDTH),
		19930 => to_signed(30892, LUT_AMPL_WIDTH),
		19931 => to_signed(30891, LUT_AMPL_WIDTH),
		19932 => to_signed(30889, LUT_AMPL_WIDTH),
		19933 => to_signed(30888, LUT_AMPL_WIDTH),
		19934 => to_signed(30887, LUT_AMPL_WIDTH),
		19935 => to_signed(30886, LUT_AMPL_WIDTH),
		19936 => to_signed(30885, LUT_AMPL_WIDTH),
		19937 => to_signed(30884, LUT_AMPL_WIDTH),
		19938 => to_signed(30883, LUT_AMPL_WIDTH),
		19939 => to_signed(30882, LUT_AMPL_WIDTH),
		19940 => to_signed(30881, LUT_AMPL_WIDTH),
		19941 => to_signed(30880, LUT_AMPL_WIDTH),
		19942 => to_signed(30879, LUT_AMPL_WIDTH),
		19943 => to_signed(30878, LUT_AMPL_WIDTH),
		19944 => to_signed(30877, LUT_AMPL_WIDTH),
		19945 => to_signed(30876, LUT_AMPL_WIDTH),
		19946 => to_signed(30875, LUT_AMPL_WIDTH),
		19947 => to_signed(30874, LUT_AMPL_WIDTH),
		19948 => to_signed(30873, LUT_AMPL_WIDTH),
		19949 => to_signed(30872, LUT_AMPL_WIDTH),
		19950 => to_signed(30871, LUT_AMPL_WIDTH),
		19951 => to_signed(30870, LUT_AMPL_WIDTH),
		19952 => to_signed(30868, LUT_AMPL_WIDTH),
		19953 => to_signed(30867, LUT_AMPL_WIDTH),
		19954 => to_signed(30866, LUT_AMPL_WIDTH),
		19955 => to_signed(30865, LUT_AMPL_WIDTH),
		19956 => to_signed(30864, LUT_AMPL_WIDTH),
		19957 => to_signed(30863, LUT_AMPL_WIDTH),
		19958 => to_signed(30862, LUT_AMPL_WIDTH),
		19959 => to_signed(30861, LUT_AMPL_WIDTH),
		19960 => to_signed(30860, LUT_AMPL_WIDTH),
		19961 => to_signed(30859, LUT_AMPL_WIDTH),
		19962 => to_signed(30858, LUT_AMPL_WIDTH),
		19963 => to_signed(30857, LUT_AMPL_WIDTH),
		19964 => to_signed(30856, LUT_AMPL_WIDTH),
		19965 => to_signed(30855, LUT_AMPL_WIDTH),
		19966 => to_signed(30854, LUT_AMPL_WIDTH),
		19967 => to_signed(30853, LUT_AMPL_WIDTH),
		19968 => to_signed(30852, LUT_AMPL_WIDTH),
		19969 => to_signed(30851, LUT_AMPL_WIDTH),
		19970 => to_signed(30849, LUT_AMPL_WIDTH),
		19971 => to_signed(30848, LUT_AMPL_WIDTH),
		19972 => to_signed(30847, LUT_AMPL_WIDTH),
		19973 => to_signed(30846, LUT_AMPL_WIDTH),
		19974 => to_signed(30845, LUT_AMPL_WIDTH),
		19975 => to_signed(30844, LUT_AMPL_WIDTH),
		19976 => to_signed(30843, LUT_AMPL_WIDTH),
		19977 => to_signed(30842, LUT_AMPL_WIDTH),
		19978 => to_signed(30841, LUT_AMPL_WIDTH),
		19979 => to_signed(30840, LUT_AMPL_WIDTH),
		19980 => to_signed(30839, LUT_AMPL_WIDTH),
		19981 => to_signed(30838, LUT_AMPL_WIDTH),
		19982 => to_signed(30837, LUT_AMPL_WIDTH),
		19983 => to_signed(30836, LUT_AMPL_WIDTH),
		19984 => to_signed(30835, LUT_AMPL_WIDTH),
		19985 => to_signed(30834, LUT_AMPL_WIDTH),
		19986 => to_signed(30832, LUT_AMPL_WIDTH),
		19987 => to_signed(30831, LUT_AMPL_WIDTH),
		19988 => to_signed(30830, LUT_AMPL_WIDTH),
		19989 => to_signed(30829, LUT_AMPL_WIDTH),
		19990 => to_signed(30828, LUT_AMPL_WIDTH),
		19991 => to_signed(30827, LUT_AMPL_WIDTH),
		19992 => to_signed(30826, LUT_AMPL_WIDTH),
		19993 => to_signed(30825, LUT_AMPL_WIDTH),
		19994 => to_signed(30824, LUT_AMPL_WIDTH),
		19995 => to_signed(30823, LUT_AMPL_WIDTH),
		19996 => to_signed(30822, LUT_AMPL_WIDTH),
		19997 => to_signed(30821, LUT_AMPL_WIDTH),
		19998 => to_signed(30820, LUT_AMPL_WIDTH),
		19999 => to_signed(30819, LUT_AMPL_WIDTH),
		20000 => to_signed(30818, LUT_AMPL_WIDTH),
		20001 => to_signed(30816, LUT_AMPL_WIDTH),
		20002 => to_signed(30815, LUT_AMPL_WIDTH),
		20003 => to_signed(30814, LUT_AMPL_WIDTH),
		20004 => to_signed(30813, LUT_AMPL_WIDTH),
		20005 => to_signed(30812, LUT_AMPL_WIDTH),
		20006 => to_signed(30811, LUT_AMPL_WIDTH),
		20007 => to_signed(30810, LUT_AMPL_WIDTH),
		20008 => to_signed(30809, LUT_AMPL_WIDTH),
		20009 => to_signed(30808, LUT_AMPL_WIDTH),
		20010 => to_signed(30807, LUT_AMPL_WIDTH),
		20011 => to_signed(30806, LUT_AMPL_WIDTH),
		20012 => to_signed(30805, LUT_AMPL_WIDTH),
		20013 => to_signed(30804, LUT_AMPL_WIDTH),
		20014 => to_signed(30803, LUT_AMPL_WIDTH),
		20015 => to_signed(30802, LUT_AMPL_WIDTH),
		20016 => to_signed(30800, LUT_AMPL_WIDTH),
		20017 => to_signed(30799, LUT_AMPL_WIDTH),
		20018 => to_signed(30798, LUT_AMPL_WIDTH),
		20019 => to_signed(30797, LUT_AMPL_WIDTH),
		20020 => to_signed(30796, LUT_AMPL_WIDTH),
		20021 => to_signed(30795, LUT_AMPL_WIDTH),
		20022 => to_signed(30794, LUT_AMPL_WIDTH),
		20023 => to_signed(30793, LUT_AMPL_WIDTH),
		20024 => to_signed(30792, LUT_AMPL_WIDTH),
		20025 => to_signed(30791, LUT_AMPL_WIDTH),
		20026 => to_signed(30790, LUT_AMPL_WIDTH),
		20027 => to_signed(30789, LUT_AMPL_WIDTH),
		20028 => to_signed(30788, LUT_AMPL_WIDTH),
		20029 => to_signed(30786, LUT_AMPL_WIDTH),
		20030 => to_signed(30785, LUT_AMPL_WIDTH),
		20031 => to_signed(30784, LUT_AMPL_WIDTH),
		20032 => to_signed(30783, LUT_AMPL_WIDTH),
		20033 => to_signed(30782, LUT_AMPL_WIDTH),
		20034 => to_signed(30781, LUT_AMPL_WIDTH),
		20035 => to_signed(30780, LUT_AMPL_WIDTH),
		20036 => to_signed(30779, LUT_AMPL_WIDTH),
		20037 => to_signed(30778, LUT_AMPL_WIDTH),
		20038 => to_signed(30777, LUT_AMPL_WIDTH),
		20039 => to_signed(30776, LUT_AMPL_WIDTH),
		20040 => to_signed(30775, LUT_AMPL_WIDTH),
		20041 => to_signed(30774, LUT_AMPL_WIDTH),
		20042 => to_signed(30772, LUT_AMPL_WIDTH),
		20043 => to_signed(30771, LUT_AMPL_WIDTH),
		20044 => to_signed(30770, LUT_AMPL_WIDTH),
		20045 => to_signed(30769, LUT_AMPL_WIDTH),
		20046 => to_signed(30768, LUT_AMPL_WIDTH),
		20047 => to_signed(30767, LUT_AMPL_WIDTH),
		20048 => to_signed(30766, LUT_AMPL_WIDTH),
		20049 => to_signed(30765, LUT_AMPL_WIDTH),
		20050 => to_signed(30764, LUT_AMPL_WIDTH),
		20051 => to_signed(30763, LUT_AMPL_WIDTH),
		20052 => to_signed(30762, LUT_AMPL_WIDTH),
		20053 => to_signed(30761, LUT_AMPL_WIDTH),
		20054 => to_signed(30760, LUT_AMPL_WIDTH),
		20055 => to_signed(30758, LUT_AMPL_WIDTH),
		20056 => to_signed(30757, LUT_AMPL_WIDTH),
		20057 => to_signed(30756, LUT_AMPL_WIDTH),
		20058 => to_signed(30755, LUT_AMPL_WIDTH),
		20059 => to_signed(30754, LUT_AMPL_WIDTH),
		20060 => to_signed(30753, LUT_AMPL_WIDTH),
		20061 => to_signed(30752, LUT_AMPL_WIDTH),
		20062 => to_signed(30751, LUT_AMPL_WIDTH),
		20063 => to_signed(30750, LUT_AMPL_WIDTH),
		20064 => to_signed(30749, LUT_AMPL_WIDTH),
		20065 => to_signed(30748, LUT_AMPL_WIDTH),
		20066 => to_signed(30746, LUT_AMPL_WIDTH),
		20067 => to_signed(30745, LUT_AMPL_WIDTH),
		20068 => to_signed(30744, LUT_AMPL_WIDTH),
		20069 => to_signed(30743, LUT_AMPL_WIDTH),
		20070 => to_signed(30742, LUT_AMPL_WIDTH),
		20071 => to_signed(30741, LUT_AMPL_WIDTH),
		20072 => to_signed(30740, LUT_AMPL_WIDTH),
		20073 => to_signed(30739, LUT_AMPL_WIDTH),
		20074 => to_signed(30738, LUT_AMPL_WIDTH),
		20075 => to_signed(30737, LUT_AMPL_WIDTH),
		20076 => to_signed(30736, LUT_AMPL_WIDTH),
		20077 => to_signed(30735, LUT_AMPL_WIDTH),
		20078 => to_signed(30733, LUT_AMPL_WIDTH),
		20079 => to_signed(30732, LUT_AMPL_WIDTH),
		20080 => to_signed(30731, LUT_AMPL_WIDTH),
		20081 => to_signed(30730, LUT_AMPL_WIDTH),
		20082 => to_signed(30729, LUT_AMPL_WIDTH),
		20083 => to_signed(30728, LUT_AMPL_WIDTH),
		20084 => to_signed(30727, LUT_AMPL_WIDTH),
		20085 => to_signed(30726, LUT_AMPL_WIDTH),
		20086 => to_signed(30725, LUT_AMPL_WIDTH),
		20087 => to_signed(30724, LUT_AMPL_WIDTH),
		20088 => to_signed(30723, LUT_AMPL_WIDTH),
		20089 => to_signed(30721, LUT_AMPL_WIDTH),
		20090 => to_signed(30720, LUT_AMPL_WIDTH),
		20091 => to_signed(30719, LUT_AMPL_WIDTH),
		20092 => to_signed(30718, LUT_AMPL_WIDTH),
		20093 => to_signed(30717, LUT_AMPL_WIDTH),
		20094 => to_signed(30716, LUT_AMPL_WIDTH),
		20095 => to_signed(30715, LUT_AMPL_WIDTH),
		20096 => to_signed(30714, LUT_AMPL_WIDTH),
		20097 => to_signed(30713, LUT_AMPL_WIDTH),
		20098 => to_signed(30712, LUT_AMPL_WIDTH),
		20099 => to_signed(30711, LUT_AMPL_WIDTH),
		20100 => to_signed(30709, LUT_AMPL_WIDTH),
		20101 => to_signed(30708, LUT_AMPL_WIDTH),
		20102 => to_signed(30707, LUT_AMPL_WIDTH),
		20103 => to_signed(30706, LUT_AMPL_WIDTH),
		20104 => to_signed(30705, LUT_AMPL_WIDTH),
		20105 => to_signed(30704, LUT_AMPL_WIDTH),
		20106 => to_signed(30703, LUT_AMPL_WIDTH),
		20107 => to_signed(30702, LUT_AMPL_WIDTH),
		20108 => to_signed(30701, LUT_AMPL_WIDTH),
		20109 => to_signed(30700, LUT_AMPL_WIDTH),
		20110 => to_signed(30698, LUT_AMPL_WIDTH),
		20111 => to_signed(30697, LUT_AMPL_WIDTH),
		20112 => to_signed(30696, LUT_AMPL_WIDTH),
		20113 => to_signed(30695, LUT_AMPL_WIDTH),
		20114 => to_signed(30694, LUT_AMPL_WIDTH),
		20115 => to_signed(30693, LUT_AMPL_WIDTH),
		20116 => to_signed(30692, LUT_AMPL_WIDTH),
		20117 => to_signed(30691, LUT_AMPL_WIDTH),
		20118 => to_signed(30690, LUT_AMPL_WIDTH),
		20119 => to_signed(30689, LUT_AMPL_WIDTH),
		20120 => to_signed(30687, LUT_AMPL_WIDTH),
		20121 => to_signed(30686, LUT_AMPL_WIDTH),
		20122 => to_signed(30685, LUT_AMPL_WIDTH),
		20123 => to_signed(30684, LUT_AMPL_WIDTH),
		20124 => to_signed(30683, LUT_AMPL_WIDTH),
		20125 => to_signed(30682, LUT_AMPL_WIDTH),
		20126 => to_signed(30681, LUT_AMPL_WIDTH),
		20127 => to_signed(30680, LUT_AMPL_WIDTH),
		20128 => to_signed(30679, LUT_AMPL_WIDTH),
		20129 => to_signed(30678, LUT_AMPL_WIDTH),
		20130 => to_signed(30676, LUT_AMPL_WIDTH),
		20131 => to_signed(30675, LUT_AMPL_WIDTH),
		20132 => to_signed(30674, LUT_AMPL_WIDTH),
		20133 => to_signed(30673, LUT_AMPL_WIDTH),
		20134 => to_signed(30672, LUT_AMPL_WIDTH),
		20135 => to_signed(30671, LUT_AMPL_WIDTH),
		20136 => to_signed(30670, LUT_AMPL_WIDTH),
		20137 => to_signed(30669, LUT_AMPL_WIDTH),
		20138 => to_signed(30668, LUT_AMPL_WIDTH),
		20139 => to_signed(30666, LUT_AMPL_WIDTH),
		20140 => to_signed(30665, LUT_AMPL_WIDTH),
		20141 => to_signed(30664, LUT_AMPL_WIDTH),
		20142 => to_signed(30663, LUT_AMPL_WIDTH),
		20143 => to_signed(30662, LUT_AMPL_WIDTH),
		20144 => to_signed(30661, LUT_AMPL_WIDTH),
		20145 => to_signed(30660, LUT_AMPL_WIDTH),
		20146 => to_signed(30659, LUT_AMPL_WIDTH),
		20147 => to_signed(30658, LUT_AMPL_WIDTH),
		20148 => to_signed(30656, LUT_AMPL_WIDTH),
		20149 => to_signed(30655, LUT_AMPL_WIDTH),
		20150 => to_signed(30654, LUT_AMPL_WIDTH),
		20151 => to_signed(30653, LUT_AMPL_WIDTH),
		20152 => to_signed(30652, LUT_AMPL_WIDTH),
		20153 => to_signed(30651, LUT_AMPL_WIDTH),
		20154 => to_signed(30650, LUT_AMPL_WIDTH),
		20155 => to_signed(30649, LUT_AMPL_WIDTH),
		20156 => to_signed(30648, LUT_AMPL_WIDTH),
		20157 => to_signed(30646, LUT_AMPL_WIDTH),
		20158 => to_signed(30645, LUT_AMPL_WIDTH),
		20159 => to_signed(30644, LUT_AMPL_WIDTH),
		20160 => to_signed(30643, LUT_AMPL_WIDTH),
		20161 => to_signed(30642, LUT_AMPL_WIDTH),
		20162 => to_signed(30641, LUT_AMPL_WIDTH),
		20163 => to_signed(30640, LUT_AMPL_WIDTH),
		20164 => to_signed(30639, LUT_AMPL_WIDTH),
		20165 => to_signed(30638, LUT_AMPL_WIDTH),
		20166 => to_signed(30636, LUT_AMPL_WIDTH),
		20167 => to_signed(30635, LUT_AMPL_WIDTH),
		20168 => to_signed(30634, LUT_AMPL_WIDTH),
		20169 => to_signed(30633, LUT_AMPL_WIDTH),
		20170 => to_signed(30632, LUT_AMPL_WIDTH),
		20171 => to_signed(30631, LUT_AMPL_WIDTH),
		20172 => to_signed(30630, LUT_AMPL_WIDTH),
		20173 => to_signed(30629, LUT_AMPL_WIDTH),
		20174 => to_signed(30628, LUT_AMPL_WIDTH),
		20175 => to_signed(30626, LUT_AMPL_WIDTH),
		20176 => to_signed(30625, LUT_AMPL_WIDTH),
		20177 => to_signed(30624, LUT_AMPL_WIDTH),
		20178 => to_signed(30623, LUT_AMPL_WIDTH),
		20179 => to_signed(30622, LUT_AMPL_WIDTH),
		20180 => to_signed(30621, LUT_AMPL_WIDTH),
		20181 => to_signed(30620, LUT_AMPL_WIDTH),
		20182 => to_signed(30619, LUT_AMPL_WIDTH),
		20183 => to_signed(30617, LUT_AMPL_WIDTH),
		20184 => to_signed(30616, LUT_AMPL_WIDTH),
		20185 => to_signed(30615, LUT_AMPL_WIDTH),
		20186 => to_signed(30614, LUT_AMPL_WIDTH),
		20187 => to_signed(30613, LUT_AMPL_WIDTH),
		20188 => to_signed(30612, LUT_AMPL_WIDTH),
		20189 => to_signed(30611, LUT_AMPL_WIDTH),
		20190 => to_signed(30610, LUT_AMPL_WIDTH),
		20191 => to_signed(30609, LUT_AMPL_WIDTH),
		20192 => to_signed(30607, LUT_AMPL_WIDTH),
		20193 => to_signed(30606, LUT_AMPL_WIDTH),
		20194 => to_signed(30605, LUT_AMPL_WIDTH),
		20195 => to_signed(30604, LUT_AMPL_WIDTH),
		20196 => to_signed(30603, LUT_AMPL_WIDTH),
		20197 => to_signed(30602, LUT_AMPL_WIDTH),
		20198 => to_signed(30601, LUT_AMPL_WIDTH),
		20199 => to_signed(30600, LUT_AMPL_WIDTH),
		20200 => to_signed(30598, LUT_AMPL_WIDTH),
		20201 => to_signed(30597, LUT_AMPL_WIDTH),
		20202 => to_signed(30596, LUT_AMPL_WIDTH),
		20203 => to_signed(30595, LUT_AMPL_WIDTH),
		20204 => to_signed(30594, LUT_AMPL_WIDTH),
		20205 => to_signed(30593, LUT_AMPL_WIDTH),
		20206 => to_signed(30592, LUT_AMPL_WIDTH),
		20207 => to_signed(30591, LUT_AMPL_WIDTH),
		20208 => to_signed(30589, LUT_AMPL_WIDTH),
		20209 => to_signed(30588, LUT_AMPL_WIDTH),
		20210 => to_signed(30587, LUT_AMPL_WIDTH),
		20211 => to_signed(30586, LUT_AMPL_WIDTH),
		20212 => to_signed(30585, LUT_AMPL_WIDTH),
		20213 => to_signed(30584, LUT_AMPL_WIDTH),
		20214 => to_signed(30583, LUT_AMPL_WIDTH),
		20215 => to_signed(30582, LUT_AMPL_WIDTH),
		20216 => to_signed(30580, LUT_AMPL_WIDTH),
		20217 => to_signed(30579, LUT_AMPL_WIDTH),
		20218 => to_signed(30578, LUT_AMPL_WIDTH),
		20219 => to_signed(30577, LUT_AMPL_WIDTH),
		20220 => to_signed(30576, LUT_AMPL_WIDTH),
		20221 => to_signed(30575, LUT_AMPL_WIDTH),
		20222 => to_signed(30574, LUT_AMPL_WIDTH),
		20223 => to_signed(30573, LUT_AMPL_WIDTH),
		20224 => to_signed(30571, LUT_AMPL_WIDTH),
		20225 => to_signed(30570, LUT_AMPL_WIDTH),
		20226 => to_signed(30569, LUT_AMPL_WIDTH),
		20227 => to_signed(30568, LUT_AMPL_WIDTH),
		20228 => to_signed(30567, LUT_AMPL_WIDTH),
		20229 => to_signed(30566, LUT_AMPL_WIDTH),
		20230 => to_signed(30565, LUT_AMPL_WIDTH),
		20231 => to_signed(30563, LUT_AMPL_WIDTH),
		20232 => to_signed(30562, LUT_AMPL_WIDTH),
		20233 => to_signed(30561, LUT_AMPL_WIDTH),
		20234 => to_signed(30560, LUT_AMPL_WIDTH),
		20235 => to_signed(30559, LUT_AMPL_WIDTH),
		20236 => to_signed(30558, LUT_AMPL_WIDTH),
		20237 => to_signed(30557, LUT_AMPL_WIDTH),
		20238 => to_signed(30556, LUT_AMPL_WIDTH),
		20239 => to_signed(30554, LUT_AMPL_WIDTH),
		20240 => to_signed(30553, LUT_AMPL_WIDTH),
		20241 => to_signed(30552, LUT_AMPL_WIDTH),
		20242 => to_signed(30551, LUT_AMPL_WIDTH),
		20243 => to_signed(30550, LUT_AMPL_WIDTH),
		20244 => to_signed(30549, LUT_AMPL_WIDTH),
		20245 => to_signed(30548, LUT_AMPL_WIDTH),
		20246 => to_signed(30546, LUT_AMPL_WIDTH),
		20247 => to_signed(30545, LUT_AMPL_WIDTH),
		20248 => to_signed(30544, LUT_AMPL_WIDTH),
		20249 => to_signed(30543, LUT_AMPL_WIDTH),
		20250 => to_signed(30542, LUT_AMPL_WIDTH),
		20251 => to_signed(30541, LUT_AMPL_WIDTH),
		20252 => to_signed(30540, LUT_AMPL_WIDTH),
		20253 => to_signed(30538, LUT_AMPL_WIDTH),
		20254 => to_signed(30537, LUT_AMPL_WIDTH),
		20255 => to_signed(30536, LUT_AMPL_WIDTH),
		20256 => to_signed(30535, LUT_AMPL_WIDTH),
		20257 => to_signed(30534, LUT_AMPL_WIDTH),
		20258 => to_signed(30533, LUT_AMPL_WIDTH),
		20259 => to_signed(30532, LUT_AMPL_WIDTH),
		20260 => to_signed(30530, LUT_AMPL_WIDTH),
		20261 => to_signed(30529, LUT_AMPL_WIDTH),
		20262 => to_signed(30528, LUT_AMPL_WIDTH),
		20263 => to_signed(30527, LUT_AMPL_WIDTH),
		20264 => to_signed(30526, LUT_AMPL_WIDTH),
		20265 => to_signed(30525, LUT_AMPL_WIDTH),
		20266 => to_signed(30524, LUT_AMPL_WIDTH),
		20267 => to_signed(30522, LUT_AMPL_WIDTH),
		20268 => to_signed(30521, LUT_AMPL_WIDTH),
		20269 => to_signed(30520, LUT_AMPL_WIDTH),
		20270 => to_signed(30519, LUT_AMPL_WIDTH),
		20271 => to_signed(30518, LUT_AMPL_WIDTH),
		20272 => to_signed(30517, LUT_AMPL_WIDTH),
		20273 => to_signed(30516, LUT_AMPL_WIDTH),
		20274 => to_signed(30514, LUT_AMPL_WIDTH),
		20275 => to_signed(30513, LUT_AMPL_WIDTH),
		20276 => to_signed(30512, LUT_AMPL_WIDTH),
		20277 => to_signed(30511, LUT_AMPL_WIDTH),
		20278 => to_signed(30510, LUT_AMPL_WIDTH),
		20279 => to_signed(30509, LUT_AMPL_WIDTH),
		20280 => to_signed(30508, LUT_AMPL_WIDTH),
		20281 => to_signed(30506, LUT_AMPL_WIDTH),
		20282 => to_signed(30505, LUT_AMPL_WIDTH),
		20283 => to_signed(30504, LUT_AMPL_WIDTH),
		20284 => to_signed(30503, LUT_AMPL_WIDTH),
		20285 => to_signed(30502, LUT_AMPL_WIDTH),
		20286 => to_signed(30501, LUT_AMPL_WIDTH),
		20287 => to_signed(30500, LUT_AMPL_WIDTH),
		20288 => to_signed(30498, LUT_AMPL_WIDTH),
		20289 => to_signed(30497, LUT_AMPL_WIDTH),
		20290 => to_signed(30496, LUT_AMPL_WIDTH),
		20291 => to_signed(30495, LUT_AMPL_WIDTH),
		20292 => to_signed(30494, LUT_AMPL_WIDTH),
		20293 => to_signed(30493, LUT_AMPL_WIDTH),
		20294 => to_signed(30492, LUT_AMPL_WIDTH),
		20295 => to_signed(30490, LUT_AMPL_WIDTH),
		20296 => to_signed(30489, LUT_AMPL_WIDTH),
		20297 => to_signed(30488, LUT_AMPL_WIDTH),
		20298 => to_signed(30487, LUT_AMPL_WIDTH),
		20299 => to_signed(30486, LUT_AMPL_WIDTH),
		20300 => to_signed(30485, LUT_AMPL_WIDTH),
		20301 => to_signed(30483, LUT_AMPL_WIDTH),
		20302 => to_signed(30482, LUT_AMPL_WIDTH),
		20303 => to_signed(30481, LUT_AMPL_WIDTH),
		20304 => to_signed(30480, LUT_AMPL_WIDTH),
		20305 => to_signed(30479, LUT_AMPL_WIDTH),
		20306 => to_signed(30478, LUT_AMPL_WIDTH),
		20307 => to_signed(30477, LUT_AMPL_WIDTH),
		20308 => to_signed(30475, LUT_AMPL_WIDTH),
		20309 => to_signed(30474, LUT_AMPL_WIDTH),
		20310 => to_signed(30473, LUT_AMPL_WIDTH),
		20311 => to_signed(30472, LUT_AMPL_WIDTH),
		20312 => to_signed(30471, LUT_AMPL_WIDTH),
		20313 => to_signed(30470, LUT_AMPL_WIDTH),
		20314 => to_signed(30468, LUT_AMPL_WIDTH),
		20315 => to_signed(30467, LUT_AMPL_WIDTH),
		20316 => to_signed(30466, LUT_AMPL_WIDTH),
		20317 => to_signed(30465, LUT_AMPL_WIDTH),
		20318 => to_signed(30464, LUT_AMPL_WIDTH),
		20319 => to_signed(30463, LUT_AMPL_WIDTH),
		20320 => to_signed(30462, LUT_AMPL_WIDTH),
		20321 => to_signed(30460, LUT_AMPL_WIDTH),
		20322 => to_signed(30459, LUT_AMPL_WIDTH),
		20323 => to_signed(30458, LUT_AMPL_WIDTH),
		20324 => to_signed(30457, LUT_AMPL_WIDTH),
		20325 => to_signed(30456, LUT_AMPL_WIDTH),
		20326 => to_signed(30455, LUT_AMPL_WIDTH),
		20327 => to_signed(30453, LUT_AMPL_WIDTH),
		20328 => to_signed(30452, LUT_AMPL_WIDTH),
		20329 => to_signed(30451, LUT_AMPL_WIDTH),
		20330 => to_signed(30450, LUT_AMPL_WIDTH),
		20331 => to_signed(30449, LUT_AMPL_WIDTH),
		20332 => to_signed(30448, LUT_AMPL_WIDTH),
		20333 => to_signed(30446, LUT_AMPL_WIDTH),
		20334 => to_signed(30445, LUT_AMPL_WIDTH),
		20335 => to_signed(30444, LUT_AMPL_WIDTH),
		20336 => to_signed(30443, LUT_AMPL_WIDTH),
		20337 => to_signed(30442, LUT_AMPL_WIDTH),
		20338 => to_signed(30441, LUT_AMPL_WIDTH),
		20339 => to_signed(30439, LUT_AMPL_WIDTH),
		20340 => to_signed(30438, LUT_AMPL_WIDTH),
		20341 => to_signed(30437, LUT_AMPL_WIDTH),
		20342 => to_signed(30436, LUT_AMPL_WIDTH),
		20343 => to_signed(30435, LUT_AMPL_WIDTH),
		20344 => to_signed(30434, LUT_AMPL_WIDTH),
		20345 => to_signed(30433, LUT_AMPL_WIDTH),
		20346 => to_signed(30431, LUT_AMPL_WIDTH),
		20347 => to_signed(30430, LUT_AMPL_WIDTH),
		20348 => to_signed(30429, LUT_AMPL_WIDTH),
		20349 => to_signed(30428, LUT_AMPL_WIDTH),
		20350 => to_signed(30427, LUT_AMPL_WIDTH),
		20351 => to_signed(30426, LUT_AMPL_WIDTH),
		20352 => to_signed(30424, LUT_AMPL_WIDTH),
		20353 => to_signed(30423, LUT_AMPL_WIDTH),
		20354 => to_signed(30422, LUT_AMPL_WIDTH),
		20355 => to_signed(30421, LUT_AMPL_WIDTH),
		20356 => to_signed(30420, LUT_AMPL_WIDTH),
		20357 => to_signed(30419, LUT_AMPL_WIDTH),
		20358 => to_signed(30417, LUT_AMPL_WIDTH),
		20359 => to_signed(30416, LUT_AMPL_WIDTH),
		20360 => to_signed(30415, LUT_AMPL_WIDTH),
		20361 => to_signed(30414, LUT_AMPL_WIDTH),
		20362 => to_signed(30413, LUT_AMPL_WIDTH),
		20363 => to_signed(30412, LUT_AMPL_WIDTH),
		20364 => to_signed(30410, LUT_AMPL_WIDTH),
		20365 => to_signed(30409, LUT_AMPL_WIDTH),
		20366 => to_signed(30408, LUT_AMPL_WIDTH),
		20367 => to_signed(30407, LUT_AMPL_WIDTH),
		20368 => to_signed(30406, LUT_AMPL_WIDTH),
		20369 => to_signed(30404, LUT_AMPL_WIDTH),
		20370 => to_signed(30403, LUT_AMPL_WIDTH),
		20371 => to_signed(30402, LUT_AMPL_WIDTH),
		20372 => to_signed(30401, LUT_AMPL_WIDTH),
		20373 => to_signed(30400, LUT_AMPL_WIDTH),
		20374 => to_signed(30399, LUT_AMPL_WIDTH),
		20375 => to_signed(30397, LUT_AMPL_WIDTH),
		20376 => to_signed(30396, LUT_AMPL_WIDTH),
		20377 => to_signed(30395, LUT_AMPL_WIDTH),
		20378 => to_signed(30394, LUT_AMPL_WIDTH),
		20379 => to_signed(30393, LUT_AMPL_WIDTH),
		20380 => to_signed(30392, LUT_AMPL_WIDTH),
		20381 => to_signed(30390, LUT_AMPL_WIDTH),
		20382 => to_signed(30389, LUT_AMPL_WIDTH),
		20383 => to_signed(30388, LUT_AMPL_WIDTH),
		20384 => to_signed(30387, LUT_AMPL_WIDTH),
		20385 => to_signed(30386, LUT_AMPL_WIDTH),
		20386 => to_signed(30385, LUT_AMPL_WIDTH),
		20387 => to_signed(30383, LUT_AMPL_WIDTH),
		20388 => to_signed(30382, LUT_AMPL_WIDTH),
		20389 => to_signed(30381, LUT_AMPL_WIDTH),
		20390 => to_signed(30380, LUT_AMPL_WIDTH),
		20391 => to_signed(30379, LUT_AMPL_WIDTH),
		20392 => to_signed(30377, LUT_AMPL_WIDTH),
		20393 => to_signed(30376, LUT_AMPL_WIDTH),
		20394 => to_signed(30375, LUT_AMPL_WIDTH),
		20395 => to_signed(30374, LUT_AMPL_WIDTH),
		20396 => to_signed(30373, LUT_AMPL_WIDTH),
		20397 => to_signed(30372, LUT_AMPL_WIDTH),
		20398 => to_signed(30370, LUT_AMPL_WIDTH),
		20399 => to_signed(30369, LUT_AMPL_WIDTH),
		20400 => to_signed(30368, LUT_AMPL_WIDTH),
		20401 => to_signed(30367, LUT_AMPL_WIDTH),
		20402 => to_signed(30366, LUT_AMPL_WIDTH),
		20403 => to_signed(30365, LUT_AMPL_WIDTH),
		20404 => to_signed(30363, LUT_AMPL_WIDTH),
		20405 => to_signed(30362, LUT_AMPL_WIDTH),
		20406 => to_signed(30361, LUT_AMPL_WIDTH),
		20407 => to_signed(30360, LUT_AMPL_WIDTH),
		20408 => to_signed(30359, LUT_AMPL_WIDTH),
		20409 => to_signed(30357, LUT_AMPL_WIDTH),
		20410 => to_signed(30356, LUT_AMPL_WIDTH),
		20411 => to_signed(30355, LUT_AMPL_WIDTH),
		20412 => to_signed(30354, LUT_AMPL_WIDTH),
		20413 => to_signed(30353, LUT_AMPL_WIDTH),
		20414 => to_signed(30351, LUT_AMPL_WIDTH),
		20415 => to_signed(30350, LUT_AMPL_WIDTH),
		20416 => to_signed(30349, LUT_AMPL_WIDTH),
		20417 => to_signed(30348, LUT_AMPL_WIDTH),
		20418 => to_signed(30347, LUT_AMPL_WIDTH),
		20419 => to_signed(30346, LUT_AMPL_WIDTH),
		20420 => to_signed(30344, LUT_AMPL_WIDTH),
		20421 => to_signed(30343, LUT_AMPL_WIDTH),
		20422 => to_signed(30342, LUT_AMPL_WIDTH),
		20423 => to_signed(30341, LUT_AMPL_WIDTH),
		20424 => to_signed(30340, LUT_AMPL_WIDTH),
		20425 => to_signed(30338, LUT_AMPL_WIDTH),
		20426 => to_signed(30337, LUT_AMPL_WIDTH),
		20427 => to_signed(30336, LUT_AMPL_WIDTH),
		20428 => to_signed(30335, LUT_AMPL_WIDTH),
		20429 => to_signed(30334, LUT_AMPL_WIDTH),
		20430 => to_signed(30333, LUT_AMPL_WIDTH),
		20431 => to_signed(30331, LUT_AMPL_WIDTH),
		20432 => to_signed(30330, LUT_AMPL_WIDTH),
		20433 => to_signed(30329, LUT_AMPL_WIDTH),
		20434 => to_signed(30328, LUT_AMPL_WIDTH),
		20435 => to_signed(30327, LUT_AMPL_WIDTH),
		20436 => to_signed(30325, LUT_AMPL_WIDTH),
		20437 => to_signed(30324, LUT_AMPL_WIDTH),
		20438 => to_signed(30323, LUT_AMPL_WIDTH),
		20439 => to_signed(30322, LUT_AMPL_WIDTH),
		20440 => to_signed(30321, LUT_AMPL_WIDTH),
		20441 => to_signed(30319, LUT_AMPL_WIDTH),
		20442 => to_signed(30318, LUT_AMPL_WIDTH),
		20443 => to_signed(30317, LUT_AMPL_WIDTH),
		20444 => to_signed(30316, LUT_AMPL_WIDTH),
		20445 => to_signed(30315, LUT_AMPL_WIDTH),
		20446 => to_signed(30313, LUT_AMPL_WIDTH),
		20447 => to_signed(30312, LUT_AMPL_WIDTH),
		20448 => to_signed(30311, LUT_AMPL_WIDTH),
		20449 => to_signed(30310, LUT_AMPL_WIDTH),
		20450 => to_signed(30309, LUT_AMPL_WIDTH),
		20451 => to_signed(30308, LUT_AMPL_WIDTH),
		20452 => to_signed(30306, LUT_AMPL_WIDTH),
		20453 => to_signed(30305, LUT_AMPL_WIDTH),
		20454 => to_signed(30304, LUT_AMPL_WIDTH),
		20455 => to_signed(30303, LUT_AMPL_WIDTH),
		20456 => to_signed(30302, LUT_AMPL_WIDTH),
		20457 => to_signed(30300, LUT_AMPL_WIDTH),
		20458 => to_signed(30299, LUT_AMPL_WIDTH),
		20459 => to_signed(30298, LUT_AMPL_WIDTH),
		20460 => to_signed(30297, LUT_AMPL_WIDTH),
		20461 => to_signed(30296, LUT_AMPL_WIDTH),
		20462 => to_signed(30294, LUT_AMPL_WIDTH),
		20463 => to_signed(30293, LUT_AMPL_WIDTH),
		20464 => to_signed(30292, LUT_AMPL_WIDTH),
		20465 => to_signed(30291, LUT_AMPL_WIDTH),
		20466 => to_signed(30290, LUT_AMPL_WIDTH),
		20467 => to_signed(30288, LUT_AMPL_WIDTH),
		20468 => to_signed(30287, LUT_AMPL_WIDTH),
		20469 => to_signed(30286, LUT_AMPL_WIDTH),
		20470 => to_signed(30285, LUT_AMPL_WIDTH),
		20471 => to_signed(30284, LUT_AMPL_WIDTH),
		20472 => to_signed(30282, LUT_AMPL_WIDTH),
		20473 => to_signed(30281, LUT_AMPL_WIDTH),
		20474 => to_signed(30280, LUT_AMPL_WIDTH),
		20475 => to_signed(30279, LUT_AMPL_WIDTH),
		20476 => to_signed(30278, LUT_AMPL_WIDTH),
		20477 => to_signed(30276, LUT_AMPL_WIDTH),
		20478 => to_signed(30275, LUT_AMPL_WIDTH),
		20479 => to_signed(30274, LUT_AMPL_WIDTH),
		20480 => to_signed(30273, LUT_AMPL_WIDTH),
		20481 => to_signed(30272, LUT_AMPL_WIDTH),
		20482 => to_signed(30270, LUT_AMPL_WIDTH),
		20483 => to_signed(30269, LUT_AMPL_WIDTH),
		20484 => to_signed(30268, LUT_AMPL_WIDTH),
		20485 => to_signed(30267, LUT_AMPL_WIDTH),
		20486 => to_signed(30266, LUT_AMPL_WIDTH),
		20487 => to_signed(30264, LUT_AMPL_WIDTH),
		20488 => to_signed(30263, LUT_AMPL_WIDTH),
		20489 => to_signed(30262, LUT_AMPL_WIDTH),
		20490 => to_signed(30261, LUT_AMPL_WIDTH),
		20491 => to_signed(30260, LUT_AMPL_WIDTH),
		20492 => to_signed(30258, LUT_AMPL_WIDTH),
		20493 => to_signed(30257, LUT_AMPL_WIDTH),
		20494 => to_signed(30256, LUT_AMPL_WIDTH),
		20495 => to_signed(30255, LUT_AMPL_WIDTH),
		20496 => to_signed(30253, LUT_AMPL_WIDTH),
		20497 => to_signed(30252, LUT_AMPL_WIDTH),
		20498 => to_signed(30251, LUT_AMPL_WIDTH),
		20499 => to_signed(30250, LUT_AMPL_WIDTH),
		20500 => to_signed(30249, LUT_AMPL_WIDTH),
		20501 => to_signed(30247, LUT_AMPL_WIDTH),
		20502 => to_signed(30246, LUT_AMPL_WIDTH),
		20503 => to_signed(30245, LUT_AMPL_WIDTH),
		20504 => to_signed(30244, LUT_AMPL_WIDTH),
		20505 => to_signed(30243, LUT_AMPL_WIDTH),
		20506 => to_signed(30241, LUT_AMPL_WIDTH),
		20507 => to_signed(30240, LUT_AMPL_WIDTH),
		20508 => to_signed(30239, LUT_AMPL_WIDTH),
		20509 => to_signed(30238, LUT_AMPL_WIDTH),
		20510 => to_signed(30237, LUT_AMPL_WIDTH),
		20511 => to_signed(30235, LUT_AMPL_WIDTH),
		20512 => to_signed(30234, LUT_AMPL_WIDTH),
		20513 => to_signed(30233, LUT_AMPL_WIDTH),
		20514 => to_signed(30232, LUT_AMPL_WIDTH),
		20515 => to_signed(30231, LUT_AMPL_WIDTH),
		20516 => to_signed(30229, LUT_AMPL_WIDTH),
		20517 => to_signed(30228, LUT_AMPL_WIDTH),
		20518 => to_signed(30227, LUT_AMPL_WIDTH),
		20519 => to_signed(30226, LUT_AMPL_WIDTH),
		20520 => to_signed(30224, LUT_AMPL_WIDTH),
		20521 => to_signed(30223, LUT_AMPL_WIDTH),
		20522 => to_signed(30222, LUT_AMPL_WIDTH),
		20523 => to_signed(30221, LUT_AMPL_WIDTH),
		20524 => to_signed(30220, LUT_AMPL_WIDTH),
		20525 => to_signed(30218, LUT_AMPL_WIDTH),
		20526 => to_signed(30217, LUT_AMPL_WIDTH),
		20527 => to_signed(30216, LUT_AMPL_WIDTH),
		20528 => to_signed(30215, LUT_AMPL_WIDTH),
		20529 => to_signed(30214, LUT_AMPL_WIDTH),
		20530 => to_signed(30212, LUT_AMPL_WIDTH),
		20531 => to_signed(30211, LUT_AMPL_WIDTH),
		20532 => to_signed(30210, LUT_AMPL_WIDTH),
		20533 => to_signed(30209, LUT_AMPL_WIDTH),
		20534 => to_signed(30207, LUT_AMPL_WIDTH),
		20535 => to_signed(30206, LUT_AMPL_WIDTH),
		20536 => to_signed(30205, LUT_AMPL_WIDTH),
		20537 => to_signed(30204, LUT_AMPL_WIDTH),
		20538 => to_signed(30203, LUT_AMPL_WIDTH),
		20539 => to_signed(30201, LUT_AMPL_WIDTH),
		20540 => to_signed(30200, LUT_AMPL_WIDTH),
		20541 => to_signed(30199, LUT_AMPL_WIDTH),
		20542 => to_signed(30198, LUT_AMPL_WIDTH),
		20543 => to_signed(30196, LUT_AMPL_WIDTH),
		20544 => to_signed(30195, LUT_AMPL_WIDTH),
		20545 => to_signed(30194, LUT_AMPL_WIDTH),
		20546 => to_signed(30193, LUT_AMPL_WIDTH),
		20547 => to_signed(30192, LUT_AMPL_WIDTH),
		20548 => to_signed(30190, LUT_AMPL_WIDTH),
		20549 => to_signed(30189, LUT_AMPL_WIDTH),
		20550 => to_signed(30188, LUT_AMPL_WIDTH),
		20551 => to_signed(30187, LUT_AMPL_WIDTH),
		20552 => to_signed(30185, LUT_AMPL_WIDTH),
		20553 => to_signed(30184, LUT_AMPL_WIDTH),
		20554 => to_signed(30183, LUT_AMPL_WIDTH),
		20555 => to_signed(30182, LUT_AMPL_WIDTH),
		20556 => to_signed(30181, LUT_AMPL_WIDTH),
		20557 => to_signed(30179, LUT_AMPL_WIDTH),
		20558 => to_signed(30178, LUT_AMPL_WIDTH),
		20559 => to_signed(30177, LUT_AMPL_WIDTH),
		20560 => to_signed(30176, LUT_AMPL_WIDTH),
		20561 => to_signed(30174, LUT_AMPL_WIDTH),
		20562 => to_signed(30173, LUT_AMPL_WIDTH),
		20563 => to_signed(30172, LUT_AMPL_WIDTH),
		20564 => to_signed(30171, LUT_AMPL_WIDTH),
		20565 => to_signed(30170, LUT_AMPL_WIDTH),
		20566 => to_signed(30168, LUT_AMPL_WIDTH),
		20567 => to_signed(30167, LUT_AMPL_WIDTH),
		20568 => to_signed(30166, LUT_AMPL_WIDTH),
		20569 => to_signed(30165, LUT_AMPL_WIDTH),
		20570 => to_signed(30163, LUT_AMPL_WIDTH),
		20571 => to_signed(30162, LUT_AMPL_WIDTH),
		20572 => to_signed(30161, LUT_AMPL_WIDTH),
		20573 => to_signed(30160, LUT_AMPL_WIDTH),
		20574 => to_signed(30159, LUT_AMPL_WIDTH),
		20575 => to_signed(30157, LUT_AMPL_WIDTH),
		20576 => to_signed(30156, LUT_AMPL_WIDTH),
		20577 => to_signed(30155, LUT_AMPL_WIDTH),
		20578 => to_signed(30154, LUT_AMPL_WIDTH),
		20579 => to_signed(30152, LUT_AMPL_WIDTH),
		20580 => to_signed(30151, LUT_AMPL_WIDTH),
		20581 => to_signed(30150, LUT_AMPL_WIDTH),
		20582 => to_signed(30149, LUT_AMPL_WIDTH),
		20583 => to_signed(30147, LUT_AMPL_WIDTH),
		20584 => to_signed(30146, LUT_AMPL_WIDTH),
		20585 => to_signed(30145, LUT_AMPL_WIDTH),
		20586 => to_signed(30144, LUT_AMPL_WIDTH),
		20587 => to_signed(30143, LUT_AMPL_WIDTH),
		20588 => to_signed(30141, LUT_AMPL_WIDTH),
		20589 => to_signed(30140, LUT_AMPL_WIDTH),
		20590 => to_signed(30139, LUT_AMPL_WIDTH),
		20591 => to_signed(30138, LUT_AMPL_WIDTH),
		20592 => to_signed(30136, LUT_AMPL_WIDTH),
		20593 => to_signed(30135, LUT_AMPL_WIDTH),
		20594 => to_signed(30134, LUT_AMPL_WIDTH),
		20595 => to_signed(30133, LUT_AMPL_WIDTH),
		20596 => to_signed(30131, LUT_AMPL_WIDTH),
		20597 => to_signed(30130, LUT_AMPL_WIDTH),
		20598 => to_signed(30129, LUT_AMPL_WIDTH),
		20599 => to_signed(30128, LUT_AMPL_WIDTH),
		20600 => to_signed(30126, LUT_AMPL_WIDTH),
		20601 => to_signed(30125, LUT_AMPL_WIDTH),
		20602 => to_signed(30124, LUT_AMPL_WIDTH),
		20603 => to_signed(30123, LUT_AMPL_WIDTH),
		20604 => to_signed(30122, LUT_AMPL_WIDTH),
		20605 => to_signed(30120, LUT_AMPL_WIDTH),
		20606 => to_signed(30119, LUT_AMPL_WIDTH),
		20607 => to_signed(30118, LUT_AMPL_WIDTH),
		20608 => to_signed(30117, LUT_AMPL_WIDTH),
		20609 => to_signed(30115, LUT_AMPL_WIDTH),
		20610 => to_signed(30114, LUT_AMPL_WIDTH),
		20611 => to_signed(30113, LUT_AMPL_WIDTH),
		20612 => to_signed(30112, LUT_AMPL_WIDTH),
		20613 => to_signed(30110, LUT_AMPL_WIDTH),
		20614 => to_signed(30109, LUT_AMPL_WIDTH),
		20615 => to_signed(30108, LUT_AMPL_WIDTH),
		20616 => to_signed(30107, LUT_AMPL_WIDTH),
		20617 => to_signed(30105, LUT_AMPL_WIDTH),
		20618 => to_signed(30104, LUT_AMPL_WIDTH),
		20619 => to_signed(30103, LUT_AMPL_WIDTH),
		20620 => to_signed(30102, LUT_AMPL_WIDTH),
		20621 => to_signed(30100, LUT_AMPL_WIDTH),
		20622 => to_signed(30099, LUT_AMPL_WIDTH),
		20623 => to_signed(30098, LUT_AMPL_WIDTH),
		20624 => to_signed(30097, LUT_AMPL_WIDTH),
		20625 => to_signed(30096, LUT_AMPL_WIDTH),
		20626 => to_signed(30094, LUT_AMPL_WIDTH),
		20627 => to_signed(30093, LUT_AMPL_WIDTH),
		20628 => to_signed(30092, LUT_AMPL_WIDTH),
		20629 => to_signed(30091, LUT_AMPL_WIDTH),
		20630 => to_signed(30089, LUT_AMPL_WIDTH),
		20631 => to_signed(30088, LUT_AMPL_WIDTH),
		20632 => to_signed(30087, LUT_AMPL_WIDTH),
		20633 => to_signed(30086, LUT_AMPL_WIDTH),
		20634 => to_signed(30084, LUT_AMPL_WIDTH),
		20635 => to_signed(30083, LUT_AMPL_WIDTH),
		20636 => to_signed(30082, LUT_AMPL_WIDTH),
		20637 => to_signed(30081, LUT_AMPL_WIDTH),
		20638 => to_signed(30079, LUT_AMPL_WIDTH),
		20639 => to_signed(30078, LUT_AMPL_WIDTH),
		20640 => to_signed(30077, LUT_AMPL_WIDTH),
		20641 => to_signed(30076, LUT_AMPL_WIDTH),
		20642 => to_signed(30074, LUT_AMPL_WIDTH),
		20643 => to_signed(30073, LUT_AMPL_WIDTH),
		20644 => to_signed(30072, LUT_AMPL_WIDTH),
		20645 => to_signed(30071, LUT_AMPL_WIDTH),
		20646 => to_signed(30069, LUT_AMPL_WIDTH),
		20647 => to_signed(30068, LUT_AMPL_WIDTH),
		20648 => to_signed(30067, LUT_AMPL_WIDTH),
		20649 => to_signed(30066, LUT_AMPL_WIDTH),
		20650 => to_signed(30064, LUT_AMPL_WIDTH),
		20651 => to_signed(30063, LUT_AMPL_WIDTH),
		20652 => to_signed(30062, LUT_AMPL_WIDTH),
		20653 => to_signed(30061, LUT_AMPL_WIDTH),
		20654 => to_signed(30059, LUT_AMPL_WIDTH),
		20655 => to_signed(30058, LUT_AMPL_WIDTH),
		20656 => to_signed(30057, LUT_AMPL_WIDTH),
		20657 => to_signed(30056, LUT_AMPL_WIDTH),
		20658 => to_signed(30054, LUT_AMPL_WIDTH),
		20659 => to_signed(30053, LUT_AMPL_WIDTH),
		20660 => to_signed(30052, LUT_AMPL_WIDTH),
		20661 => to_signed(30051, LUT_AMPL_WIDTH),
		20662 => to_signed(30049, LUT_AMPL_WIDTH),
		20663 => to_signed(30048, LUT_AMPL_WIDTH),
		20664 => to_signed(30047, LUT_AMPL_WIDTH),
		20665 => to_signed(30046, LUT_AMPL_WIDTH),
		20666 => to_signed(30044, LUT_AMPL_WIDTH),
		20667 => to_signed(30043, LUT_AMPL_WIDTH),
		20668 => to_signed(30042, LUT_AMPL_WIDTH),
		20669 => to_signed(30041, LUT_AMPL_WIDTH),
		20670 => to_signed(30039, LUT_AMPL_WIDTH),
		20671 => to_signed(30038, LUT_AMPL_WIDTH),
		20672 => to_signed(30037, LUT_AMPL_WIDTH),
		20673 => to_signed(30036, LUT_AMPL_WIDTH),
		20674 => to_signed(30034, LUT_AMPL_WIDTH),
		20675 => to_signed(30033, LUT_AMPL_WIDTH),
		20676 => to_signed(30032, LUT_AMPL_WIDTH),
		20677 => to_signed(30031, LUT_AMPL_WIDTH),
		20678 => to_signed(30029, LUT_AMPL_WIDTH),
		20679 => to_signed(30028, LUT_AMPL_WIDTH),
		20680 => to_signed(30027, LUT_AMPL_WIDTH),
		20681 => to_signed(30026, LUT_AMPL_WIDTH),
		20682 => to_signed(30024, LUT_AMPL_WIDTH),
		20683 => to_signed(30023, LUT_AMPL_WIDTH),
		20684 => to_signed(30022, LUT_AMPL_WIDTH),
		20685 => to_signed(30020, LUT_AMPL_WIDTH),
		20686 => to_signed(30019, LUT_AMPL_WIDTH),
		20687 => to_signed(30018, LUT_AMPL_WIDTH),
		20688 => to_signed(30017, LUT_AMPL_WIDTH),
		20689 => to_signed(30015, LUT_AMPL_WIDTH),
		20690 => to_signed(30014, LUT_AMPL_WIDTH),
		20691 => to_signed(30013, LUT_AMPL_WIDTH),
		20692 => to_signed(30012, LUT_AMPL_WIDTH),
		20693 => to_signed(30010, LUT_AMPL_WIDTH),
		20694 => to_signed(30009, LUT_AMPL_WIDTH),
		20695 => to_signed(30008, LUT_AMPL_WIDTH),
		20696 => to_signed(30007, LUT_AMPL_WIDTH),
		20697 => to_signed(30005, LUT_AMPL_WIDTH),
		20698 => to_signed(30004, LUT_AMPL_WIDTH),
		20699 => to_signed(30003, LUT_AMPL_WIDTH),
		20700 => to_signed(30002, LUT_AMPL_WIDTH),
		20701 => to_signed(30000, LUT_AMPL_WIDTH),
		20702 => to_signed(29999, LUT_AMPL_WIDTH),
		20703 => to_signed(29998, LUT_AMPL_WIDTH),
		20704 => to_signed(29997, LUT_AMPL_WIDTH),
		20705 => to_signed(29995, LUT_AMPL_WIDTH),
		20706 => to_signed(29994, LUT_AMPL_WIDTH),
		20707 => to_signed(29993, LUT_AMPL_WIDTH),
		20708 => to_signed(29991, LUT_AMPL_WIDTH),
		20709 => to_signed(29990, LUT_AMPL_WIDTH),
		20710 => to_signed(29989, LUT_AMPL_WIDTH),
		20711 => to_signed(29988, LUT_AMPL_WIDTH),
		20712 => to_signed(29986, LUT_AMPL_WIDTH),
		20713 => to_signed(29985, LUT_AMPL_WIDTH),
		20714 => to_signed(29984, LUT_AMPL_WIDTH),
		20715 => to_signed(29983, LUT_AMPL_WIDTH),
		20716 => to_signed(29981, LUT_AMPL_WIDTH),
		20717 => to_signed(29980, LUT_AMPL_WIDTH),
		20718 => to_signed(29979, LUT_AMPL_WIDTH),
		20719 => to_signed(29978, LUT_AMPL_WIDTH),
		20720 => to_signed(29976, LUT_AMPL_WIDTH),
		20721 => to_signed(29975, LUT_AMPL_WIDTH),
		20722 => to_signed(29974, LUT_AMPL_WIDTH),
		20723 => to_signed(29972, LUT_AMPL_WIDTH),
		20724 => to_signed(29971, LUT_AMPL_WIDTH),
		20725 => to_signed(29970, LUT_AMPL_WIDTH),
		20726 => to_signed(29969, LUT_AMPL_WIDTH),
		20727 => to_signed(29967, LUT_AMPL_WIDTH),
		20728 => to_signed(29966, LUT_AMPL_WIDTH),
		20729 => to_signed(29965, LUT_AMPL_WIDTH),
		20730 => to_signed(29964, LUT_AMPL_WIDTH),
		20731 => to_signed(29962, LUT_AMPL_WIDTH),
		20732 => to_signed(29961, LUT_AMPL_WIDTH),
		20733 => to_signed(29960, LUT_AMPL_WIDTH),
		20734 => to_signed(29958, LUT_AMPL_WIDTH),
		20735 => to_signed(29957, LUT_AMPL_WIDTH),
		20736 => to_signed(29956, LUT_AMPL_WIDTH),
		20737 => to_signed(29955, LUT_AMPL_WIDTH),
		20738 => to_signed(29953, LUT_AMPL_WIDTH),
		20739 => to_signed(29952, LUT_AMPL_WIDTH),
		20740 => to_signed(29951, LUT_AMPL_WIDTH),
		20741 => to_signed(29950, LUT_AMPL_WIDTH),
		20742 => to_signed(29948, LUT_AMPL_WIDTH),
		20743 => to_signed(29947, LUT_AMPL_WIDTH),
		20744 => to_signed(29946, LUT_AMPL_WIDTH),
		20745 => to_signed(29944, LUT_AMPL_WIDTH),
		20746 => to_signed(29943, LUT_AMPL_WIDTH),
		20747 => to_signed(29942, LUT_AMPL_WIDTH),
		20748 => to_signed(29941, LUT_AMPL_WIDTH),
		20749 => to_signed(29939, LUT_AMPL_WIDTH),
		20750 => to_signed(29938, LUT_AMPL_WIDTH),
		20751 => to_signed(29937, LUT_AMPL_WIDTH),
		20752 => to_signed(29936, LUT_AMPL_WIDTH),
		20753 => to_signed(29934, LUT_AMPL_WIDTH),
		20754 => to_signed(29933, LUT_AMPL_WIDTH),
		20755 => to_signed(29932, LUT_AMPL_WIDTH),
		20756 => to_signed(29930, LUT_AMPL_WIDTH),
		20757 => to_signed(29929, LUT_AMPL_WIDTH),
		20758 => to_signed(29928, LUT_AMPL_WIDTH),
		20759 => to_signed(29927, LUT_AMPL_WIDTH),
		20760 => to_signed(29925, LUT_AMPL_WIDTH),
		20761 => to_signed(29924, LUT_AMPL_WIDTH),
		20762 => to_signed(29923, LUT_AMPL_WIDTH),
		20763 => to_signed(29921, LUT_AMPL_WIDTH),
		20764 => to_signed(29920, LUT_AMPL_WIDTH),
		20765 => to_signed(29919, LUT_AMPL_WIDTH),
		20766 => to_signed(29918, LUT_AMPL_WIDTH),
		20767 => to_signed(29916, LUT_AMPL_WIDTH),
		20768 => to_signed(29915, LUT_AMPL_WIDTH),
		20769 => to_signed(29914, LUT_AMPL_WIDTH),
		20770 => to_signed(29912, LUT_AMPL_WIDTH),
		20771 => to_signed(29911, LUT_AMPL_WIDTH),
		20772 => to_signed(29910, LUT_AMPL_WIDTH),
		20773 => to_signed(29909, LUT_AMPL_WIDTH),
		20774 => to_signed(29907, LUT_AMPL_WIDTH),
		20775 => to_signed(29906, LUT_AMPL_WIDTH),
		20776 => to_signed(29905, LUT_AMPL_WIDTH),
		20777 => to_signed(29903, LUT_AMPL_WIDTH),
		20778 => to_signed(29902, LUT_AMPL_WIDTH),
		20779 => to_signed(29901, LUT_AMPL_WIDTH),
		20780 => to_signed(29900, LUT_AMPL_WIDTH),
		20781 => to_signed(29898, LUT_AMPL_WIDTH),
		20782 => to_signed(29897, LUT_AMPL_WIDTH),
		20783 => to_signed(29896, LUT_AMPL_WIDTH),
		20784 => to_signed(29894, LUT_AMPL_WIDTH),
		20785 => to_signed(29893, LUT_AMPL_WIDTH),
		20786 => to_signed(29892, LUT_AMPL_WIDTH),
		20787 => to_signed(29891, LUT_AMPL_WIDTH),
		20788 => to_signed(29889, LUT_AMPL_WIDTH),
		20789 => to_signed(29888, LUT_AMPL_WIDTH),
		20790 => to_signed(29887, LUT_AMPL_WIDTH),
		20791 => to_signed(29885, LUT_AMPL_WIDTH),
		20792 => to_signed(29884, LUT_AMPL_WIDTH),
		20793 => to_signed(29883, LUT_AMPL_WIDTH),
		20794 => to_signed(29882, LUT_AMPL_WIDTH),
		20795 => to_signed(29880, LUT_AMPL_WIDTH),
		20796 => to_signed(29879, LUT_AMPL_WIDTH),
		20797 => to_signed(29878, LUT_AMPL_WIDTH),
		20798 => to_signed(29876, LUT_AMPL_WIDTH),
		20799 => to_signed(29875, LUT_AMPL_WIDTH),
		20800 => to_signed(29874, LUT_AMPL_WIDTH),
		20801 => to_signed(29873, LUT_AMPL_WIDTH),
		20802 => to_signed(29871, LUT_AMPL_WIDTH),
		20803 => to_signed(29870, LUT_AMPL_WIDTH),
		20804 => to_signed(29869, LUT_AMPL_WIDTH),
		20805 => to_signed(29867, LUT_AMPL_WIDTH),
		20806 => to_signed(29866, LUT_AMPL_WIDTH),
		20807 => to_signed(29865, LUT_AMPL_WIDTH),
		20808 => to_signed(29864, LUT_AMPL_WIDTH),
		20809 => to_signed(29862, LUT_AMPL_WIDTH),
		20810 => to_signed(29861, LUT_AMPL_WIDTH),
		20811 => to_signed(29860, LUT_AMPL_WIDTH),
		20812 => to_signed(29858, LUT_AMPL_WIDTH),
		20813 => to_signed(29857, LUT_AMPL_WIDTH),
		20814 => to_signed(29856, LUT_AMPL_WIDTH),
		20815 => to_signed(29854, LUT_AMPL_WIDTH),
		20816 => to_signed(29853, LUT_AMPL_WIDTH),
		20817 => to_signed(29852, LUT_AMPL_WIDTH),
		20818 => to_signed(29851, LUT_AMPL_WIDTH),
		20819 => to_signed(29849, LUT_AMPL_WIDTH),
		20820 => to_signed(29848, LUT_AMPL_WIDTH),
		20821 => to_signed(29847, LUT_AMPL_WIDTH),
		20822 => to_signed(29845, LUT_AMPL_WIDTH),
		20823 => to_signed(29844, LUT_AMPL_WIDTH),
		20824 => to_signed(29843, LUT_AMPL_WIDTH),
		20825 => to_signed(29842, LUT_AMPL_WIDTH),
		20826 => to_signed(29840, LUT_AMPL_WIDTH),
		20827 => to_signed(29839, LUT_AMPL_WIDTH),
		20828 => to_signed(29838, LUT_AMPL_WIDTH),
		20829 => to_signed(29836, LUT_AMPL_WIDTH),
		20830 => to_signed(29835, LUT_AMPL_WIDTH),
		20831 => to_signed(29834, LUT_AMPL_WIDTH),
		20832 => to_signed(29832, LUT_AMPL_WIDTH),
		20833 => to_signed(29831, LUT_AMPL_WIDTH),
		20834 => to_signed(29830, LUT_AMPL_WIDTH),
		20835 => to_signed(29829, LUT_AMPL_WIDTH),
		20836 => to_signed(29827, LUT_AMPL_WIDTH),
		20837 => to_signed(29826, LUT_AMPL_WIDTH),
		20838 => to_signed(29825, LUT_AMPL_WIDTH),
		20839 => to_signed(29823, LUT_AMPL_WIDTH),
		20840 => to_signed(29822, LUT_AMPL_WIDTH),
		20841 => to_signed(29821, LUT_AMPL_WIDTH),
		20842 => to_signed(29819, LUT_AMPL_WIDTH),
		20843 => to_signed(29818, LUT_AMPL_WIDTH),
		20844 => to_signed(29817, LUT_AMPL_WIDTH),
		20845 => to_signed(29816, LUT_AMPL_WIDTH),
		20846 => to_signed(29814, LUT_AMPL_WIDTH),
		20847 => to_signed(29813, LUT_AMPL_WIDTH),
		20848 => to_signed(29812, LUT_AMPL_WIDTH),
		20849 => to_signed(29810, LUT_AMPL_WIDTH),
		20850 => to_signed(29809, LUT_AMPL_WIDTH),
		20851 => to_signed(29808, LUT_AMPL_WIDTH),
		20852 => to_signed(29806, LUT_AMPL_WIDTH),
		20853 => to_signed(29805, LUT_AMPL_WIDTH),
		20854 => to_signed(29804, LUT_AMPL_WIDTH),
		20855 => to_signed(29802, LUT_AMPL_WIDTH),
		20856 => to_signed(29801, LUT_AMPL_WIDTH),
		20857 => to_signed(29800, LUT_AMPL_WIDTH),
		20858 => to_signed(29799, LUT_AMPL_WIDTH),
		20859 => to_signed(29797, LUT_AMPL_WIDTH),
		20860 => to_signed(29796, LUT_AMPL_WIDTH),
		20861 => to_signed(29795, LUT_AMPL_WIDTH),
		20862 => to_signed(29793, LUT_AMPL_WIDTH),
		20863 => to_signed(29792, LUT_AMPL_WIDTH),
		20864 => to_signed(29791, LUT_AMPL_WIDTH),
		20865 => to_signed(29789, LUT_AMPL_WIDTH),
		20866 => to_signed(29788, LUT_AMPL_WIDTH),
		20867 => to_signed(29787, LUT_AMPL_WIDTH),
		20868 => to_signed(29785, LUT_AMPL_WIDTH),
		20869 => to_signed(29784, LUT_AMPL_WIDTH),
		20870 => to_signed(29783, LUT_AMPL_WIDTH),
		20871 => to_signed(29782, LUT_AMPL_WIDTH),
		20872 => to_signed(29780, LUT_AMPL_WIDTH),
		20873 => to_signed(29779, LUT_AMPL_WIDTH),
		20874 => to_signed(29778, LUT_AMPL_WIDTH),
		20875 => to_signed(29776, LUT_AMPL_WIDTH),
		20876 => to_signed(29775, LUT_AMPL_WIDTH),
		20877 => to_signed(29774, LUT_AMPL_WIDTH),
		20878 => to_signed(29772, LUT_AMPL_WIDTH),
		20879 => to_signed(29771, LUT_AMPL_WIDTH),
		20880 => to_signed(29770, LUT_AMPL_WIDTH),
		20881 => to_signed(29768, LUT_AMPL_WIDTH),
		20882 => to_signed(29767, LUT_AMPL_WIDTH),
		20883 => to_signed(29766, LUT_AMPL_WIDTH),
		20884 => to_signed(29764, LUT_AMPL_WIDTH),
		20885 => to_signed(29763, LUT_AMPL_WIDTH),
		20886 => to_signed(29762, LUT_AMPL_WIDTH),
		20887 => to_signed(29761, LUT_AMPL_WIDTH),
		20888 => to_signed(29759, LUT_AMPL_WIDTH),
		20889 => to_signed(29758, LUT_AMPL_WIDTH),
		20890 => to_signed(29757, LUT_AMPL_WIDTH),
		20891 => to_signed(29755, LUT_AMPL_WIDTH),
		20892 => to_signed(29754, LUT_AMPL_WIDTH),
		20893 => to_signed(29753, LUT_AMPL_WIDTH),
		20894 => to_signed(29751, LUT_AMPL_WIDTH),
		20895 => to_signed(29750, LUT_AMPL_WIDTH),
		20896 => to_signed(29749, LUT_AMPL_WIDTH),
		20897 => to_signed(29747, LUT_AMPL_WIDTH),
		20898 => to_signed(29746, LUT_AMPL_WIDTH),
		20899 => to_signed(29745, LUT_AMPL_WIDTH),
		20900 => to_signed(29743, LUT_AMPL_WIDTH),
		20901 => to_signed(29742, LUT_AMPL_WIDTH),
		20902 => to_signed(29741, LUT_AMPL_WIDTH),
		20903 => to_signed(29739, LUT_AMPL_WIDTH),
		20904 => to_signed(29738, LUT_AMPL_WIDTH),
		20905 => to_signed(29737, LUT_AMPL_WIDTH),
		20906 => to_signed(29736, LUT_AMPL_WIDTH),
		20907 => to_signed(29734, LUT_AMPL_WIDTH),
		20908 => to_signed(29733, LUT_AMPL_WIDTH),
		20909 => to_signed(29732, LUT_AMPL_WIDTH),
		20910 => to_signed(29730, LUT_AMPL_WIDTH),
		20911 => to_signed(29729, LUT_AMPL_WIDTH),
		20912 => to_signed(29728, LUT_AMPL_WIDTH),
		20913 => to_signed(29726, LUT_AMPL_WIDTH),
		20914 => to_signed(29725, LUT_AMPL_WIDTH),
		20915 => to_signed(29724, LUT_AMPL_WIDTH),
		20916 => to_signed(29722, LUT_AMPL_WIDTH),
		20917 => to_signed(29721, LUT_AMPL_WIDTH),
		20918 => to_signed(29720, LUT_AMPL_WIDTH),
		20919 => to_signed(29718, LUT_AMPL_WIDTH),
		20920 => to_signed(29717, LUT_AMPL_WIDTH),
		20921 => to_signed(29716, LUT_AMPL_WIDTH),
		20922 => to_signed(29714, LUT_AMPL_WIDTH),
		20923 => to_signed(29713, LUT_AMPL_WIDTH),
		20924 => to_signed(29712, LUT_AMPL_WIDTH),
		20925 => to_signed(29710, LUT_AMPL_WIDTH),
		20926 => to_signed(29709, LUT_AMPL_WIDTH),
		20927 => to_signed(29708, LUT_AMPL_WIDTH),
		20928 => to_signed(29706, LUT_AMPL_WIDTH),
		20929 => to_signed(29705, LUT_AMPL_WIDTH),
		20930 => to_signed(29704, LUT_AMPL_WIDTH),
		20931 => to_signed(29702, LUT_AMPL_WIDTH),
		20932 => to_signed(29701, LUT_AMPL_WIDTH),
		20933 => to_signed(29700, LUT_AMPL_WIDTH),
		20934 => to_signed(29698, LUT_AMPL_WIDTH),
		20935 => to_signed(29697, LUT_AMPL_WIDTH),
		20936 => to_signed(29696, LUT_AMPL_WIDTH),
		20937 => to_signed(29694, LUT_AMPL_WIDTH),
		20938 => to_signed(29693, LUT_AMPL_WIDTH),
		20939 => to_signed(29692, LUT_AMPL_WIDTH),
		20940 => to_signed(29690, LUT_AMPL_WIDTH),
		20941 => to_signed(29689, LUT_AMPL_WIDTH),
		20942 => to_signed(29688, LUT_AMPL_WIDTH),
		20943 => to_signed(29687, LUT_AMPL_WIDTH),
		20944 => to_signed(29685, LUT_AMPL_WIDTH),
		20945 => to_signed(29684, LUT_AMPL_WIDTH),
		20946 => to_signed(29683, LUT_AMPL_WIDTH),
		20947 => to_signed(29681, LUT_AMPL_WIDTH),
		20948 => to_signed(29680, LUT_AMPL_WIDTH),
		20949 => to_signed(29679, LUT_AMPL_WIDTH),
		20950 => to_signed(29677, LUT_AMPL_WIDTH),
		20951 => to_signed(29676, LUT_AMPL_WIDTH),
		20952 => to_signed(29675, LUT_AMPL_WIDTH),
		20953 => to_signed(29673, LUT_AMPL_WIDTH),
		20954 => to_signed(29672, LUT_AMPL_WIDTH),
		20955 => to_signed(29671, LUT_AMPL_WIDTH),
		20956 => to_signed(29669, LUT_AMPL_WIDTH),
		20957 => to_signed(29668, LUT_AMPL_WIDTH),
		20958 => to_signed(29667, LUT_AMPL_WIDTH),
		20959 => to_signed(29665, LUT_AMPL_WIDTH),
		20960 => to_signed(29664, LUT_AMPL_WIDTH),
		20961 => to_signed(29663, LUT_AMPL_WIDTH),
		20962 => to_signed(29661, LUT_AMPL_WIDTH),
		20963 => to_signed(29660, LUT_AMPL_WIDTH),
		20964 => to_signed(29659, LUT_AMPL_WIDTH),
		20965 => to_signed(29657, LUT_AMPL_WIDTH),
		20966 => to_signed(29656, LUT_AMPL_WIDTH),
		20967 => to_signed(29655, LUT_AMPL_WIDTH),
		20968 => to_signed(29653, LUT_AMPL_WIDTH),
		20969 => to_signed(29652, LUT_AMPL_WIDTH),
		20970 => to_signed(29651, LUT_AMPL_WIDTH),
		20971 => to_signed(29649, LUT_AMPL_WIDTH),
		20972 => to_signed(29648, LUT_AMPL_WIDTH),
		20973 => to_signed(29646, LUT_AMPL_WIDTH),
		20974 => to_signed(29645, LUT_AMPL_WIDTH),
		20975 => to_signed(29644, LUT_AMPL_WIDTH),
		20976 => to_signed(29642, LUT_AMPL_WIDTH),
		20977 => to_signed(29641, LUT_AMPL_WIDTH),
		20978 => to_signed(29640, LUT_AMPL_WIDTH),
		20979 => to_signed(29638, LUT_AMPL_WIDTH),
		20980 => to_signed(29637, LUT_AMPL_WIDTH),
		20981 => to_signed(29636, LUT_AMPL_WIDTH),
		20982 => to_signed(29634, LUT_AMPL_WIDTH),
		20983 => to_signed(29633, LUT_AMPL_WIDTH),
		20984 => to_signed(29632, LUT_AMPL_WIDTH),
		20985 => to_signed(29630, LUT_AMPL_WIDTH),
		20986 => to_signed(29629, LUT_AMPL_WIDTH),
		20987 => to_signed(29628, LUT_AMPL_WIDTH),
		20988 => to_signed(29626, LUT_AMPL_WIDTH),
		20989 => to_signed(29625, LUT_AMPL_WIDTH),
		20990 => to_signed(29624, LUT_AMPL_WIDTH),
		20991 => to_signed(29622, LUT_AMPL_WIDTH),
		20992 => to_signed(29621, LUT_AMPL_WIDTH),
		20993 => to_signed(29620, LUT_AMPL_WIDTH),
		20994 => to_signed(29618, LUT_AMPL_WIDTH),
		20995 => to_signed(29617, LUT_AMPL_WIDTH),
		20996 => to_signed(29616, LUT_AMPL_WIDTH),
		20997 => to_signed(29614, LUT_AMPL_WIDTH),
		20998 => to_signed(29613, LUT_AMPL_WIDTH),
		20999 => to_signed(29612, LUT_AMPL_WIDTH),
		21000 => to_signed(29610, LUT_AMPL_WIDTH),
		21001 => to_signed(29609, LUT_AMPL_WIDTH),
		21002 => to_signed(29608, LUT_AMPL_WIDTH),
		21003 => to_signed(29606, LUT_AMPL_WIDTH),
		21004 => to_signed(29605, LUT_AMPL_WIDTH),
		21005 => to_signed(29604, LUT_AMPL_WIDTH),
		21006 => to_signed(29602, LUT_AMPL_WIDTH),
		21007 => to_signed(29601, LUT_AMPL_WIDTH),
		21008 => to_signed(29599, LUT_AMPL_WIDTH),
		21009 => to_signed(29598, LUT_AMPL_WIDTH),
		21010 => to_signed(29597, LUT_AMPL_WIDTH),
		21011 => to_signed(29595, LUT_AMPL_WIDTH),
		21012 => to_signed(29594, LUT_AMPL_WIDTH),
		21013 => to_signed(29593, LUT_AMPL_WIDTH),
		21014 => to_signed(29591, LUT_AMPL_WIDTH),
		21015 => to_signed(29590, LUT_AMPL_WIDTH),
		21016 => to_signed(29589, LUT_AMPL_WIDTH),
		21017 => to_signed(29587, LUT_AMPL_WIDTH),
		21018 => to_signed(29586, LUT_AMPL_WIDTH),
		21019 => to_signed(29585, LUT_AMPL_WIDTH),
		21020 => to_signed(29583, LUT_AMPL_WIDTH),
		21021 => to_signed(29582, LUT_AMPL_WIDTH),
		21022 => to_signed(29581, LUT_AMPL_WIDTH),
		21023 => to_signed(29579, LUT_AMPL_WIDTH),
		21024 => to_signed(29578, LUT_AMPL_WIDTH),
		21025 => to_signed(29577, LUT_AMPL_WIDTH),
		21026 => to_signed(29575, LUT_AMPL_WIDTH),
		21027 => to_signed(29574, LUT_AMPL_WIDTH),
		21028 => to_signed(29572, LUT_AMPL_WIDTH),
		21029 => to_signed(29571, LUT_AMPL_WIDTH),
		21030 => to_signed(29570, LUT_AMPL_WIDTH),
		21031 => to_signed(29568, LUT_AMPL_WIDTH),
		21032 => to_signed(29567, LUT_AMPL_WIDTH),
		21033 => to_signed(29566, LUT_AMPL_WIDTH),
		21034 => to_signed(29564, LUT_AMPL_WIDTH),
		21035 => to_signed(29563, LUT_AMPL_WIDTH),
		21036 => to_signed(29562, LUT_AMPL_WIDTH),
		21037 => to_signed(29560, LUT_AMPL_WIDTH),
		21038 => to_signed(29559, LUT_AMPL_WIDTH),
		21039 => to_signed(29558, LUT_AMPL_WIDTH),
		21040 => to_signed(29556, LUT_AMPL_WIDTH),
		21041 => to_signed(29555, LUT_AMPL_WIDTH),
		21042 => to_signed(29554, LUT_AMPL_WIDTH),
		21043 => to_signed(29552, LUT_AMPL_WIDTH),
		21044 => to_signed(29551, LUT_AMPL_WIDTH),
		21045 => to_signed(29549, LUT_AMPL_WIDTH),
		21046 => to_signed(29548, LUT_AMPL_WIDTH),
		21047 => to_signed(29547, LUT_AMPL_WIDTH),
		21048 => to_signed(29545, LUT_AMPL_WIDTH),
		21049 => to_signed(29544, LUT_AMPL_WIDTH),
		21050 => to_signed(29543, LUT_AMPL_WIDTH),
		21051 => to_signed(29541, LUT_AMPL_WIDTH),
		21052 => to_signed(29540, LUT_AMPL_WIDTH),
		21053 => to_signed(29539, LUT_AMPL_WIDTH),
		21054 => to_signed(29537, LUT_AMPL_WIDTH),
		21055 => to_signed(29536, LUT_AMPL_WIDTH),
		21056 => to_signed(29534, LUT_AMPL_WIDTH),
		21057 => to_signed(29533, LUT_AMPL_WIDTH),
		21058 => to_signed(29532, LUT_AMPL_WIDTH),
		21059 => to_signed(29530, LUT_AMPL_WIDTH),
		21060 => to_signed(29529, LUT_AMPL_WIDTH),
		21061 => to_signed(29528, LUT_AMPL_WIDTH),
		21062 => to_signed(29526, LUT_AMPL_WIDTH),
		21063 => to_signed(29525, LUT_AMPL_WIDTH),
		21064 => to_signed(29524, LUT_AMPL_WIDTH),
		21065 => to_signed(29522, LUT_AMPL_WIDTH),
		21066 => to_signed(29521, LUT_AMPL_WIDTH),
		21067 => to_signed(29520, LUT_AMPL_WIDTH),
		21068 => to_signed(29518, LUT_AMPL_WIDTH),
		21069 => to_signed(29517, LUT_AMPL_WIDTH),
		21070 => to_signed(29515, LUT_AMPL_WIDTH),
		21071 => to_signed(29514, LUT_AMPL_WIDTH),
		21072 => to_signed(29513, LUT_AMPL_WIDTH),
		21073 => to_signed(29511, LUT_AMPL_WIDTH),
		21074 => to_signed(29510, LUT_AMPL_WIDTH),
		21075 => to_signed(29509, LUT_AMPL_WIDTH),
		21076 => to_signed(29507, LUT_AMPL_WIDTH),
		21077 => to_signed(29506, LUT_AMPL_WIDTH),
		21078 => to_signed(29504, LUT_AMPL_WIDTH),
		21079 => to_signed(29503, LUT_AMPL_WIDTH),
		21080 => to_signed(29502, LUT_AMPL_WIDTH),
		21081 => to_signed(29500, LUT_AMPL_WIDTH),
		21082 => to_signed(29499, LUT_AMPL_WIDTH),
		21083 => to_signed(29498, LUT_AMPL_WIDTH),
		21084 => to_signed(29496, LUT_AMPL_WIDTH),
		21085 => to_signed(29495, LUT_AMPL_WIDTH),
		21086 => to_signed(29494, LUT_AMPL_WIDTH),
		21087 => to_signed(29492, LUT_AMPL_WIDTH),
		21088 => to_signed(29491, LUT_AMPL_WIDTH),
		21089 => to_signed(29489, LUT_AMPL_WIDTH),
		21090 => to_signed(29488, LUT_AMPL_WIDTH),
		21091 => to_signed(29487, LUT_AMPL_WIDTH),
		21092 => to_signed(29485, LUT_AMPL_WIDTH),
		21093 => to_signed(29484, LUT_AMPL_WIDTH),
		21094 => to_signed(29483, LUT_AMPL_WIDTH),
		21095 => to_signed(29481, LUT_AMPL_WIDTH),
		21096 => to_signed(29480, LUT_AMPL_WIDTH),
		21097 => to_signed(29478, LUT_AMPL_WIDTH),
		21098 => to_signed(29477, LUT_AMPL_WIDTH),
		21099 => to_signed(29476, LUT_AMPL_WIDTH),
		21100 => to_signed(29474, LUT_AMPL_WIDTH),
		21101 => to_signed(29473, LUT_AMPL_WIDTH),
		21102 => to_signed(29472, LUT_AMPL_WIDTH),
		21103 => to_signed(29470, LUT_AMPL_WIDTH),
		21104 => to_signed(29469, LUT_AMPL_WIDTH),
		21105 => to_signed(29468, LUT_AMPL_WIDTH),
		21106 => to_signed(29466, LUT_AMPL_WIDTH),
		21107 => to_signed(29465, LUT_AMPL_WIDTH),
		21108 => to_signed(29463, LUT_AMPL_WIDTH),
		21109 => to_signed(29462, LUT_AMPL_WIDTH),
		21110 => to_signed(29461, LUT_AMPL_WIDTH),
		21111 => to_signed(29459, LUT_AMPL_WIDTH),
		21112 => to_signed(29458, LUT_AMPL_WIDTH),
		21113 => to_signed(29457, LUT_AMPL_WIDTH),
		21114 => to_signed(29455, LUT_AMPL_WIDTH),
		21115 => to_signed(29454, LUT_AMPL_WIDTH),
		21116 => to_signed(29452, LUT_AMPL_WIDTH),
		21117 => to_signed(29451, LUT_AMPL_WIDTH),
		21118 => to_signed(29450, LUT_AMPL_WIDTH),
		21119 => to_signed(29448, LUT_AMPL_WIDTH),
		21120 => to_signed(29447, LUT_AMPL_WIDTH),
		21121 => to_signed(29445, LUT_AMPL_WIDTH),
		21122 => to_signed(29444, LUT_AMPL_WIDTH),
		21123 => to_signed(29443, LUT_AMPL_WIDTH),
		21124 => to_signed(29441, LUT_AMPL_WIDTH),
		21125 => to_signed(29440, LUT_AMPL_WIDTH),
		21126 => to_signed(29439, LUT_AMPL_WIDTH),
		21127 => to_signed(29437, LUT_AMPL_WIDTH),
		21128 => to_signed(29436, LUT_AMPL_WIDTH),
		21129 => to_signed(29434, LUT_AMPL_WIDTH),
		21130 => to_signed(29433, LUT_AMPL_WIDTH),
		21131 => to_signed(29432, LUT_AMPL_WIDTH),
		21132 => to_signed(29430, LUT_AMPL_WIDTH),
		21133 => to_signed(29429, LUT_AMPL_WIDTH),
		21134 => to_signed(29428, LUT_AMPL_WIDTH),
		21135 => to_signed(29426, LUT_AMPL_WIDTH),
		21136 => to_signed(29425, LUT_AMPL_WIDTH),
		21137 => to_signed(29423, LUT_AMPL_WIDTH),
		21138 => to_signed(29422, LUT_AMPL_WIDTH),
		21139 => to_signed(29421, LUT_AMPL_WIDTH),
		21140 => to_signed(29419, LUT_AMPL_WIDTH),
		21141 => to_signed(29418, LUT_AMPL_WIDTH),
		21142 => to_signed(29416, LUT_AMPL_WIDTH),
		21143 => to_signed(29415, LUT_AMPL_WIDTH),
		21144 => to_signed(29414, LUT_AMPL_WIDTH),
		21145 => to_signed(29412, LUT_AMPL_WIDTH),
		21146 => to_signed(29411, LUT_AMPL_WIDTH),
		21147 => to_signed(29410, LUT_AMPL_WIDTH),
		21148 => to_signed(29408, LUT_AMPL_WIDTH),
		21149 => to_signed(29407, LUT_AMPL_WIDTH),
		21150 => to_signed(29405, LUT_AMPL_WIDTH),
		21151 => to_signed(29404, LUT_AMPL_WIDTH),
		21152 => to_signed(29403, LUT_AMPL_WIDTH),
		21153 => to_signed(29401, LUT_AMPL_WIDTH),
		21154 => to_signed(29400, LUT_AMPL_WIDTH),
		21155 => to_signed(29398, LUT_AMPL_WIDTH),
		21156 => to_signed(29397, LUT_AMPL_WIDTH),
		21157 => to_signed(29396, LUT_AMPL_WIDTH),
		21158 => to_signed(29394, LUT_AMPL_WIDTH),
		21159 => to_signed(29393, LUT_AMPL_WIDTH),
		21160 => to_signed(29392, LUT_AMPL_WIDTH),
		21161 => to_signed(29390, LUT_AMPL_WIDTH),
		21162 => to_signed(29389, LUT_AMPL_WIDTH),
		21163 => to_signed(29387, LUT_AMPL_WIDTH),
		21164 => to_signed(29386, LUT_AMPL_WIDTH),
		21165 => to_signed(29385, LUT_AMPL_WIDTH),
		21166 => to_signed(29383, LUT_AMPL_WIDTH),
		21167 => to_signed(29382, LUT_AMPL_WIDTH),
		21168 => to_signed(29380, LUT_AMPL_WIDTH),
		21169 => to_signed(29379, LUT_AMPL_WIDTH),
		21170 => to_signed(29378, LUT_AMPL_WIDTH),
		21171 => to_signed(29376, LUT_AMPL_WIDTH),
		21172 => to_signed(29375, LUT_AMPL_WIDTH),
		21173 => to_signed(29373, LUT_AMPL_WIDTH),
		21174 => to_signed(29372, LUT_AMPL_WIDTH),
		21175 => to_signed(29371, LUT_AMPL_WIDTH),
		21176 => to_signed(29369, LUT_AMPL_WIDTH),
		21177 => to_signed(29368, LUT_AMPL_WIDTH),
		21178 => to_signed(29366, LUT_AMPL_WIDTH),
		21179 => to_signed(29365, LUT_AMPL_WIDTH),
		21180 => to_signed(29364, LUT_AMPL_WIDTH),
		21181 => to_signed(29362, LUT_AMPL_WIDTH),
		21182 => to_signed(29361, LUT_AMPL_WIDTH),
		21183 => to_signed(29360, LUT_AMPL_WIDTH),
		21184 => to_signed(29358, LUT_AMPL_WIDTH),
		21185 => to_signed(29357, LUT_AMPL_WIDTH),
		21186 => to_signed(29355, LUT_AMPL_WIDTH),
		21187 => to_signed(29354, LUT_AMPL_WIDTH),
		21188 => to_signed(29353, LUT_AMPL_WIDTH),
		21189 => to_signed(29351, LUT_AMPL_WIDTH),
		21190 => to_signed(29350, LUT_AMPL_WIDTH),
		21191 => to_signed(29348, LUT_AMPL_WIDTH),
		21192 => to_signed(29347, LUT_AMPL_WIDTH),
		21193 => to_signed(29346, LUT_AMPL_WIDTH),
		21194 => to_signed(29344, LUT_AMPL_WIDTH),
		21195 => to_signed(29343, LUT_AMPL_WIDTH),
		21196 => to_signed(29341, LUT_AMPL_WIDTH),
		21197 => to_signed(29340, LUT_AMPL_WIDTH),
		21198 => to_signed(29339, LUT_AMPL_WIDTH),
		21199 => to_signed(29337, LUT_AMPL_WIDTH),
		21200 => to_signed(29336, LUT_AMPL_WIDTH),
		21201 => to_signed(29334, LUT_AMPL_WIDTH),
		21202 => to_signed(29333, LUT_AMPL_WIDTH),
		21203 => to_signed(29332, LUT_AMPL_WIDTH),
		21204 => to_signed(29330, LUT_AMPL_WIDTH),
		21205 => to_signed(29329, LUT_AMPL_WIDTH),
		21206 => to_signed(29327, LUT_AMPL_WIDTH),
		21207 => to_signed(29326, LUT_AMPL_WIDTH),
		21208 => to_signed(29325, LUT_AMPL_WIDTH),
		21209 => to_signed(29323, LUT_AMPL_WIDTH),
		21210 => to_signed(29322, LUT_AMPL_WIDTH),
		21211 => to_signed(29320, LUT_AMPL_WIDTH),
		21212 => to_signed(29319, LUT_AMPL_WIDTH),
		21213 => to_signed(29318, LUT_AMPL_WIDTH),
		21214 => to_signed(29316, LUT_AMPL_WIDTH),
		21215 => to_signed(29315, LUT_AMPL_WIDTH),
		21216 => to_signed(29313, LUT_AMPL_WIDTH),
		21217 => to_signed(29312, LUT_AMPL_WIDTH),
		21218 => to_signed(29311, LUT_AMPL_WIDTH),
		21219 => to_signed(29309, LUT_AMPL_WIDTH),
		21220 => to_signed(29308, LUT_AMPL_WIDTH),
		21221 => to_signed(29306, LUT_AMPL_WIDTH),
		21222 => to_signed(29305, LUT_AMPL_WIDTH),
		21223 => to_signed(29304, LUT_AMPL_WIDTH),
		21224 => to_signed(29302, LUT_AMPL_WIDTH),
		21225 => to_signed(29301, LUT_AMPL_WIDTH),
		21226 => to_signed(29299, LUT_AMPL_WIDTH),
		21227 => to_signed(29298, LUT_AMPL_WIDTH),
		21228 => to_signed(29296, LUT_AMPL_WIDTH),
		21229 => to_signed(29295, LUT_AMPL_WIDTH),
		21230 => to_signed(29294, LUT_AMPL_WIDTH),
		21231 => to_signed(29292, LUT_AMPL_WIDTH),
		21232 => to_signed(29291, LUT_AMPL_WIDTH),
		21233 => to_signed(29289, LUT_AMPL_WIDTH),
		21234 => to_signed(29288, LUT_AMPL_WIDTH),
		21235 => to_signed(29287, LUT_AMPL_WIDTH),
		21236 => to_signed(29285, LUT_AMPL_WIDTH),
		21237 => to_signed(29284, LUT_AMPL_WIDTH),
		21238 => to_signed(29282, LUT_AMPL_WIDTH),
		21239 => to_signed(29281, LUT_AMPL_WIDTH),
		21240 => to_signed(29280, LUT_AMPL_WIDTH),
		21241 => to_signed(29278, LUT_AMPL_WIDTH),
		21242 => to_signed(29277, LUT_AMPL_WIDTH),
		21243 => to_signed(29275, LUT_AMPL_WIDTH),
		21244 => to_signed(29274, LUT_AMPL_WIDTH),
		21245 => to_signed(29273, LUT_AMPL_WIDTH),
		21246 => to_signed(29271, LUT_AMPL_WIDTH),
		21247 => to_signed(29270, LUT_AMPL_WIDTH),
		21248 => to_signed(29268, LUT_AMPL_WIDTH),
		21249 => to_signed(29267, LUT_AMPL_WIDTH),
		21250 => to_signed(29265, LUT_AMPL_WIDTH),
		21251 => to_signed(29264, LUT_AMPL_WIDTH),
		21252 => to_signed(29263, LUT_AMPL_WIDTH),
		21253 => to_signed(29261, LUT_AMPL_WIDTH),
		21254 => to_signed(29260, LUT_AMPL_WIDTH),
		21255 => to_signed(29258, LUT_AMPL_WIDTH),
		21256 => to_signed(29257, LUT_AMPL_WIDTH),
		21257 => to_signed(29256, LUT_AMPL_WIDTH),
		21258 => to_signed(29254, LUT_AMPL_WIDTH),
		21259 => to_signed(29253, LUT_AMPL_WIDTH),
		21260 => to_signed(29251, LUT_AMPL_WIDTH),
		21261 => to_signed(29250, LUT_AMPL_WIDTH),
		21262 => to_signed(29248, LUT_AMPL_WIDTH),
		21263 => to_signed(29247, LUT_AMPL_WIDTH),
		21264 => to_signed(29246, LUT_AMPL_WIDTH),
		21265 => to_signed(29244, LUT_AMPL_WIDTH),
		21266 => to_signed(29243, LUT_AMPL_WIDTH),
		21267 => to_signed(29241, LUT_AMPL_WIDTH),
		21268 => to_signed(29240, LUT_AMPL_WIDTH),
		21269 => to_signed(29239, LUT_AMPL_WIDTH),
		21270 => to_signed(29237, LUT_AMPL_WIDTH),
		21271 => to_signed(29236, LUT_AMPL_WIDTH),
		21272 => to_signed(29234, LUT_AMPL_WIDTH),
		21273 => to_signed(29233, LUT_AMPL_WIDTH),
		21274 => to_signed(29231, LUT_AMPL_WIDTH),
		21275 => to_signed(29230, LUT_AMPL_WIDTH),
		21276 => to_signed(29229, LUT_AMPL_WIDTH),
		21277 => to_signed(29227, LUT_AMPL_WIDTH),
		21278 => to_signed(29226, LUT_AMPL_WIDTH),
		21279 => to_signed(29224, LUT_AMPL_WIDTH),
		21280 => to_signed(29223, LUT_AMPL_WIDTH),
		21281 => to_signed(29222, LUT_AMPL_WIDTH),
		21282 => to_signed(29220, LUT_AMPL_WIDTH),
		21283 => to_signed(29219, LUT_AMPL_WIDTH),
		21284 => to_signed(29217, LUT_AMPL_WIDTH),
		21285 => to_signed(29216, LUT_AMPL_WIDTH),
		21286 => to_signed(29214, LUT_AMPL_WIDTH),
		21287 => to_signed(29213, LUT_AMPL_WIDTH),
		21288 => to_signed(29212, LUT_AMPL_WIDTH),
		21289 => to_signed(29210, LUT_AMPL_WIDTH),
		21290 => to_signed(29209, LUT_AMPL_WIDTH),
		21291 => to_signed(29207, LUT_AMPL_WIDTH),
		21292 => to_signed(29206, LUT_AMPL_WIDTH),
		21293 => to_signed(29204, LUT_AMPL_WIDTH),
		21294 => to_signed(29203, LUT_AMPL_WIDTH),
		21295 => to_signed(29202, LUT_AMPL_WIDTH),
		21296 => to_signed(29200, LUT_AMPL_WIDTH),
		21297 => to_signed(29199, LUT_AMPL_WIDTH),
		21298 => to_signed(29197, LUT_AMPL_WIDTH),
		21299 => to_signed(29196, LUT_AMPL_WIDTH),
		21300 => to_signed(29194, LUT_AMPL_WIDTH),
		21301 => to_signed(29193, LUT_AMPL_WIDTH),
		21302 => to_signed(29192, LUT_AMPL_WIDTH),
		21303 => to_signed(29190, LUT_AMPL_WIDTH),
		21304 => to_signed(29189, LUT_AMPL_WIDTH),
		21305 => to_signed(29187, LUT_AMPL_WIDTH),
		21306 => to_signed(29186, LUT_AMPL_WIDTH),
		21307 => to_signed(29184, LUT_AMPL_WIDTH),
		21308 => to_signed(29183, LUT_AMPL_WIDTH),
		21309 => to_signed(29182, LUT_AMPL_WIDTH),
		21310 => to_signed(29180, LUT_AMPL_WIDTH),
		21311 => to_signed(29179, LUT_AMPL_WIDTH),
		21312 => to_signed(29177, LUT_AMPL_WIDTH),
		21313 => to_signed(29176, LUT_AMPL_WIDTH),
		21314 => to_signed(29174, LUT_AMPL_WIDTH),
		21315 => to_signed(29173, LUT_AMPL_WIDTH),
		21316 => to_signed(29172, LUT_AMPL_WIDTH),
		21317 => to_signed(29170, LUT_AMPL_WIDTH),
		21318 => to_signed(29169, LUT_AMPL_WIDTH),
		21319 => to_signed(29167, LUT_AMPL_WIDTH),
		21320 => to_signed(29166, LUT_AMPL_WIDTH),
		21321 => to_signed(29164, LUT_AMPL_WIDTH),
		21322 => to_signed(29163, LUT_AMPL_WIDTH),
		21323 => to_signed(29162, LUT_AMPL_WIDTH),
		21324 => to_signed(29160, LUT_AMPL_WIDTH),
		21325 => to_signed(29159, LUT_AMPL_WIDTH),
		21326 => to_signed(29157, LUT_AMPL_WIDTH),
		21327 => to_signed(29156, LUT_AMPL_WIDTH),
		21328 => to_signed(29154, LUT_AMPL_WIDTH),
		21329 => to_signed(29153, LUT_AMPL_WIDTH),
		21330 => to_signed(29152, LUT_AMPL_WIDTH),
		21331 => to_signed(29150, LUT_AMPL_WIDTH),
		21332 => to_signed(29149, LUT_AMPL_WIDTH),
		21333 => to_signed(29147, LUT_AMPL_WIDTH),
		21334 => to_signed(29146, LUT_AMPL_WIDTH),
		21335 => to_signed(29144, LUT_AMPL_WIDTH),
		21336 => to_signed(29143, LUT_AMPL_WIDTH),
		21337 => to_signed(29142, LUT_AMPL_WIDTH),
		21338 => to_signed(29140, LUT_AMPL_WIDTH),
		21339 => to_signed(29139, LUT_AMPL_WIDTH),
		21340 => to_signed(29137, LUT_AMPL_WIDTH),
		21341 => to_signed(29136, LUT_AMPL_WIDTH),
		21342 => to_signed(29134, LUT_AMPL_WIDTH),
		21343 => to_signed(29133, LUT_AMPL_WIDTH),
		21344 => to_signed(29131, LUT_AMPL_WIDTH),
		21345 => to_signed(29130, LUT_AMPL_WIDTH),
		21346 => to_signed(29129, LUT_AMPL_WIDTH),
		21347 => to_signed(29127, LUT_AMPL_WIDTH),
		21348 => to_signed(29126, LUT_AMPL_WIDTH),
		21349 => to_signed(29124, LUT_AMPL_WIDTH),
		21350 => to_signed(29123, LUT_AMPL_WIDTH),
		21351 => to_signed(29121, LUT_AMPL_WIDTH),
		21352 => to_signed(29120, LUT_AMPL_WIDTH),
		21353 => to_signed(29118, LUT_AMPL_WIDTH),
		21354 => to_signed(29117, LUT_AMPL_WIDTH),
		21355 => to_signed(29116, LUT_AMPL_WIDTH),
		21356 => to_signed(29114, LUT_AMPL_WIDTH),
		21357 => to_signed(29113, LUT_AMPL_WIDTH),
		21358 => to_signed(29111, LUT_AMPL_WIDTH),
		21359 => to_signed(29110, LUT_AMPL_WIDTH),
		21360 => to_signed(29108, LUT_AMPL_WIDTH),
		21361 => to_signed(29107, LUT_AMPL_WIDTH),
		21362 => to_signed(29106, LUT_AMPL_WIDTH),
		21363 => to_signed(29104, LUT_AMPL_WIDTH),
		21364 => to_signed(29103, LUT_AMPL_WIDTH),
		21365 => to_signed(29101, LUT_AMPL_WIDTH),
		21366 => to_signed(29100, LUT_AMPL_WIDTH),
		21367 => to_signed(29098, LUT_AMPL_WIDTH),
		21368 => to_signed(29097, LUT_AMPL_WIDTH),
		21369 => to_signed(29095, LUT_AMPL_WIDTH),
		21370 => to_signed(29094, LUT_AMPL_WIDTH),
		21371 => to_signed(29093, LUT_AMPL_WIDTH),
		21372 => to_signed(29091, LUT_AMPL_WIDTH),
		21373 => to_signed(29090, LUT_AMPL_WIDTH),
		21374 => to_signed(29088, LUT_AMPL_WIDTH),
		21375 => to_signed(29087, LUT_AMPL_WIDTH),
		21376 => to_signed(29085, LUT_AMPL_WIDTH),
		21377 => to_signed(29084, LUT_AMPL_WIDTH),
		21378 => to_signed(29082, LUT_AMPL_WIDTH),
		21379 => to_signed(29081, LUT_AMPL_WIDTH),
		21380 => to_signed(29079, LUT_AMPL_WIDTH),
		21381 => to_signed(29078, LUT_AMPL_WIDTH),
		21382 => to_signed(29077, LUT_AMPL_WIDTH),
		21383 => to_signed(29075, LUT_AMPL_WIDTH),
		21384 => to_signed(29074, LUT_AMPL_WIDTH),
		21385 => to_signed(29072, LUT_AMPL_WIDTH),
		21386 => to_signed(29071, LUT_AMPL_WIDTH),
		21387 => to_signed(29069, LUT_AMPL_WIDTH),
		21388 => to_signed(29068, LUT_AMPL_WIDTH),
		21389 => to_signed(29066, LUT_AMPL_WIDTH),
		21390 => to_signed(29065, LUT_AMPL_WIDTH),
		21391 => to_signed(29064, LUT_AMPL_WIDTH),
		21392 => to_signed(29062, LUT_AMPL_WIDTH),
		21393 => to_signed(29061, LUT_AMPL_WIDTH),
		21394 => to_signed(29059, LUT_AMPL_WIDTH),
		21395 => to_signed(29058, LUT_AMPL_WIDTH),
		21396 => to_signed(29056, LUT_AMPL_WIDTH),
		21397 => to_signed(29055, LUT_AMPL_WIDTH),
		21398 => to_signed(29053, LUT_AMPL_WIDTH),
		21399 => to_signed(29052, LUT_AMPL_WIDTH),
		21400 => to_signed(29050, LUT_AMPL_WIDTH),
		21401 => to_signed(29049, LUT_AMPL_WIDTH),
		21402 => to_signed(29048, LUT_AMPL_WIDTH),
		21403 => to_signed(29046, LUT_AMPL_WIDTH),
		21404 => to_signed(29045, LUT_AMPL_WIDTH),
		21405 => to_signed(29043, LUT_AMPL_WIDTH),
		21406 => to_signed(29042, LUT_AMPL_WIDTH),
		21407 => to_signed(29040, LUT_AMPL_WIDTH),
		21408 => to_signed(29039, LUT_AMPL_WIDTH),
		21409 => to_signed(29037, LUT_AMPL_WIDTH),
		21410 => to_signed(29036, LUT_AMPL_WIDTH),
		21411 => to_signed(29034, LUT_AMPL_WIDTH),
		21412 => to_signed(29033, LUT_AMPL_WIDTH),
		21413 => to_signed(29032, LUT_AMPL_WIDTH),
		21414 => to_signed(29030, LUT_AMPL_WIDTH),
		21415 => to_signed(29029, LUT_AMPL_WIDTH),
		21416 => to_signed(29027, LUT_AMPL_WIDTH),
		21417 => to_signed(29026, LUT_AMPL_WIDTH),
		21418 => to_signed(29024, LUT_AMPL_WIDTH),
		21419 => to_signed(29023, LUT_AMPL_WIDTH),
		21420 => to_signed(29021, LUT_AMPL_WIDTH),
		21421 => to_signed(29020, LUT_AMPL_WIDTH),
		21422 => to_signed(29018, LUT_AMPL_WIDTH),
		21423 => to_signed(29017, LUT_AMPL_WIDTH),
		21424 => to_signed(29016, LUT_AMPL_WIDTH),
		21425 => to_signed(29014, LUT_AMPL_WIDTH),
		21426 => to_signed(29013, LUT_AMPL_WIDTH),
		21427 => to_signed(29011, LUT_AMPL_WIDTH),
		21428 => to_signed(29010, LUT_AMPL_WIDTH),
		21429 => to_signed(29008, LUT_AMPL_WIDTH),
		21430 => to_signed(29007, LUT_AMPL_WIDTH),
		21431 => to_signed(29005, LUT_AMPL_WIDTH),
		21432 => to_signed(29004, LUT_AMPL_WIDTH),
		21433 => to_signed(29002, LUT_AMPL_WIDTH),
		21434 => to_signed(29001, LUT_AMPL_WIDTH),
		21435 => to_signed(28999, LUT_AMPL_WIDTH),
		21436 => to_signed(28998, LUT_AMPL_WIDTH),
		21437 => to_signed(28997, LUT_AMPL_WIDTH),
		21438 => to_signed(28995, LUT_AMPL_WIDTH),
		21439 => to_signed(28994, LUT_AMPL_WIDTH),
		21440 => to_signed(28992, LUT_AMPL_WIDTH),
		21441 => to_signed(28991, LUT_AMPL_WIDTH),
		21442 => to_signed(28989, LUT_AMPL_WIDTH),
		21443 => to_signed(28988, LUT_AMPL_WIDTH),
		21444 => to_signed(28986, LUT_AMPL_WIDTH),
		21445 => to_signed(28985, LUT_AMPL_WIDTH),
		21446 => to_signed(28983, LUT_AMPL_WIDTH),
		21447 => to_signed(28982, LUT_AMPL_WIDTH),
		21448 => to_signed(28980, LUT_AMPL_WIDTH),
		21449 => to_signed(28979, LUT_AMPL_WIDTH),
		21450 => to_signed(28977, LUT_AMPL_WIDTH),
		21451 => to_signed(28976, LUT_AMPL_WIDTH),
		21452 => to_signed(28975, LUT_AMPL_WIDTH),
		21453 => to_signed(28973, LUT_AMPL_WIDTH),
		21454 => to_signed(28972, LUT_AMPL_WIDTH),
		21455 => to_signed(28970, LUT_AMPL_WIDTH),
		21456 => to_signed(28969, LUT_AMPL_WIDTH),
		21457 => to_signed(28967, LUT_AMPL_WIDTH),
		21458 => to_signed(28966, LUT_AMPL_WIDTH),
		21459 => to_signed(28964, LUT_AMPL_WIDTH),
		21460 => to_signed(28963, LUT_AMPL_WIDTH),
		21461 => to_signed(28961, LUT_AMPL_WIDTH),
		21462 => to_signed(28960, LUT_AMPL_WIDTH),
		21463 => to_signed(28958, LUT_AMPL_WIDTH),
		21464 => to_signed(28957, LUT_AMPL_WIDTH),
		21465 => to_signed(28955, LUT_AMPL_WIDTH),
		21466 => to_signed(28954, LUT_AMPL_WIDTH),
		21467 => to_signed(28953, LUT_AMPL_WIDTH),
		21468 => to_signed(28951, LUT_AMPL_WIDTH),
		21469 => to_signed(28950, LUT_AMPL_WIDTH),
		21470 => to_signed(28948, LUT_AMPL_WIDTH),
		21471 => to_signed(28947, LUT_AMPL_WIDTH),
		21472 => to_signed(28945, LUT_AMPL_WIDTH),
		21473 => to_signed(28944, LUT_AMPL_WIDTH),
		21474 => to_signed(28942, LUT_AMPL_WIDTH),
		21475 => to_signed(28941, LUT_AMPL_WIDTH),
		21476 => to_signed(28939, LUT_AMPL_WIDTH),
		21477 => to_signed(28938, LUT_AMPL_WIDTH),
		21478 => to_signed(28936, LUT_AMPL_WIDTH),
		21479 => to_signed(28935, LUT_AMPL_WIDTH),
		21480 => to_signed(28933, LUT_AMPL_WIDTH),
		21481 => to_signed(28932, LUT_AMPL_WIDTH),
		21482 => to_signed(28930, LUT_AMPL_WIDTH),
		21483 => to_signed(28929, LUT_AMPL_WIDTH),
		21484 => to_signed(28927, LUT_AMPL_WIDTH),
		21485 => to_signed(28926, LUT_AMPL_WIDTH),
		21486 => to_signed(28925, LUT_AMPL_WIDTH),
		21487 => to_signed(28923, LUT_AMPL_WIDTH),
		21488 => to_signed(28922, LUT_AMPL_WIDTH),
		21489 => to_signed(28920, LUT_AMPL_WIDTH),
		21490 => to_signed(28919, LUT_AMPL_WIDTH),
		21491 => to_signed(28917, LUT_AMPL_WIDTH),
		21492 => to_signed(28916, LUT_AMPL_WIDTH),
		21493 => to_signed(28914, LUT_AMPL_WIDTH),
		21494 => to_signed(28913, LUT_AMPL_WIDTH),
		21495 => to_signed(28911, LUT_AMPL_WIDTH),
		21496 => to_signed(28910, LUT_AMPL_WIDTH),
		21497 => to_signed(28908, LUT_AMPL_WIDTH),
		21498 => to_signed(28907, LUT_AMPL_WIDTH),
		21499 => to_signed(28905, LUT_AMPL_WIDTH),
		21500 => to_signed(28904, LUT_AMPL_WIDTH),
		21501 => to_signed(28902, LUT_AMPL_WIDTH),
		21502 => to_signed(28901, LUT_AMPL_WIDTH),
		21503 => to_signed(28899, LUT_AMPL_WIDTH),
		21504 => to_signed(28898, LUT_AMPL_WIDTH),
		21505 => to_signed(28896, LUT_AMPL_WIDTH),
		21506 => to_signed(28895, LUT_AMPL_WIDTH),
		21507 => to_signed(28893, LUT_AMPL_WIDTH),
		21508 => to_signed(28892, LUT_AMPL_WIDTH),
		21509 => to_signed(28891, LUT_AMPL_WIDTH),
		21510 => to_signed(28889, LUT_AMPL_WIDTH),
		21511 => to_signed(28888, LUT_AMPL_WIDTH),
		21512 => to_signed(28886, LUT_AMPL_WIDTH),
		21513 => to_signed(28885, LUT_AMPL_WIDTH),
		21514 => to_signed(28883, LUT_AMPL_WIDTH),
		21515 => to_signed(28882, LUT_AMPL_WIDTH),
		21516 => to_signed(28880, LUT_AMPL_WIDTH),
		21517 => to_signed(28879, LUT_AMPL_WIDTH),
		21518 => to_signed(28877, LUT_AMPL_WIDTH),
		21519 => to_signed(28876, LUT_AMPL_WIDTH),
		21520 => to_signed(28874, LUT_AMPL_WIDTH),
		21521 => to_signed(28873, LUT_AMPL_WIDTH),
		21522 => to_signed(28871, LUT_AMPL_WIDTH),
		21523 => to_signed(28870, LUT_AMPL_WIDTH),
		21524 => to_signed(28868, LUT_AMPL_WIDTH),
		21525 => to_signed(28867, LUT_AMPL_WIDTH),
		21526 => to_signed(28865, LUT_AMPL_WIDTH),
		21527 => to_signed(28864, LUT_AMPL_WIDTH),
		21528 => to_signed(28862, LUT_AMPL_WIDTH),
		21529 => to_signed(28861, LUT_AMPL_WIDTH),
		21530 => to_signed(28859, LUT_AMPL_WIDTH),
		21531 => to_signed(28858, LUT_AMPL_WIDTH),
		21532 => to_signed(28856, LUT_AMPL_WIDTH),
		21533 => to_signed(28855, LUT_AMPL_WIDTH),
		21534 => to_signed(28853, LUT_AMPL_WIDTH),
		21535 => to_signed(28852, LUT_AMPL_WIDTH),
		21536 => to_signed(28850, LUT_AMPL_WIDTH),
		21537 => to_signed(28849, LUT_AMPL_WIDTH),
		21538 => to_signed(28847, LUT_AMPL_WIDTH),
		21539 => to_signed(28846, LUT_AMPL_WIDTH),
		21540 => to_signed(28844, LUT_AMPL_WIDTH),
		21541 => to_signed(28843, LUT_AMPL_WIDTH),
		21542 => to_signed(28841, LUT_AMPL_WIDTH),
		21543 => to_signed(28840, LUT_AMPL_WIDTH),
		21544 => to_signed(28838, LUT_AMPL_WIDTH),
		21545 => to_signed(28837, LUT_AMPL_WIDTH),
		21546 => to_signed(28835, LUT_AMPL_WIDTH),
		21547 => to_signed(28834, LUT_AMPL_WIDTH),
		21548 => to_signed(28832, LUT_AMPL_WIDTH),
		21549 => to_signed(28831, LUT_AMPL_WIDTH),
		21550 => to_signed(28830, LUT_AMPL_WIDTH),
		21551 => to_signed(28828, LUT_AMPL_WIDTH),
		21552 => to_signed(28827, LUT_AMPL_WIDTH),
		21553 => to_signed(28825, LUT_AMPL_WIDTH),
		21554 => to_signed(28824, LUT_AMPL_WIDTH),
		21555 => to_signed(28822, LUT_AMPL_WIDTH),
		21556 => to_signed(28821, LUT_AMPL_WIDTH),
		21557 => to_signed(28819, LUT_AMPL_WIDTH),
		21558 => to_signed(28818, LUT_AMPL_WIDTH),
		21559 => to_signed(28816, LUT_AMPL_WIDTH),
		21560 => to_signed(28815, LUT_AMPL_WIDTH),
		21561 => to_signed(28813, LUT_AMPL_WIDTH),
		21562 => to_signed(28812, LUT_AMPL_WIDTH),
		21563 => to_signed(28810, LUT_AMPL_WIDTH),
		21564 => to_signed(28809, LUT_AMPL_WIDTH),
		21565 => to_signed(28807, LUT_AMPL_WIDTH),
		21566 => to_signed(28806, LUT_AMPL_WIDTH),
		21567 => to_signed(28804, LUT_AMPL_WIDTH),
		21568 => to_signed(28803, LUT_AMPL_WIDTH),
		21569 => to_signed(28801, LUT_AMPL_WIDTH),
		21570 => to_signed(28800, LUT_AMPL_WIDTH),
		21571 => to_signed(28798, LUT_AMPL_WIDTH),
		21572 => to_signed(28797, LUT_AMPL_WIDTH),
		21573 => to_signed(28795, LUT_AMPL_WIDTH),
		21574 => to_signed(28794, LUT_AMPL_WIDTH),
		21575 => to_signed(28792, LUT_AMPL_WIDTH),
		21576 => to_signed(28791, LUT_AMPL_WIDTH),
		21577 => to_signed(28789, LUT_AMPL_WIDTH),
		21578 => to_signed(28788, LUT_AMPL_WIDTH),
		21579 => to_signed(28786, LUT_AMPL_WIDTH),
		21580 => to_signed(28785, LUT_AMPL_WIDTH),
		21581 => to_signed(28783, LUT_AMPL_WIDTH),
		21582 => to_signed(28782, LUT_AMPL_WIDTH),
		21583 => to_signed(28780, LUT_AMPL_WIDTH),
		21584 => to_signed(28779, LUT_AMPL_WIDTH),
		21585 => to_signed(28777, LUT_AMPL_WIDTH),
		21586 => to_signed(28776, LUT_AMPL_WIDTH),
		21587 => to_signed(28774, LUT_AMPL_WIDTH),
		21588 => to_signed(28773, LUT_AMPL_WIDTH),
		21589 => to_signed(28771, LUT_AMPL_WIDTH),
		21590 => to_signed(28770, LUT_AMPL_WIDTH),
		21591 => to_signed(28768, LUT_AMPL_WIDTH),
		21592 => to_signed(28767, LUT_AMPL_WIDTH),
		21593 => to_signed(28765, LUT_AMPL_WIDTH),
		21594 => to_signed(28764, LUT_AMPL_WIDTH),
		21595 => to_signed(28762, LUT_AMPL_WIDTH),
		21596 => to_signed(28761, LUT_AMPL_WIDTH),
		21597 => to_signed(28759, LUT_AMPL_WIDTH),
		21598 => to_signed(28758, LUT_AMPL_WIDTH),
		21599 => to_signed(28756, LUT_AMPL_WIDTH),
		21600 => to_signed(28755, LUT_AMPL_WIDTH),
		21601 => to_signed(28753, LUT_AMPL_WIDTH),
		21602 => to_signed(28752, LUT_AMPL_WIDTH),
		21603 => to_signed(28750, LUT_AMPL_WIDTH),
		21604 => to_signed(28748, LUT_AMPL_WIDTH),
		21605 => to_signed(28747, LUT_AMPL_WIDTH),
		21606 => to_signed(28745, LUT_AMPL_WIDTH),
		21607 => to_signed(28744, LUT_AMPL_WIDTH),
		21608 => to_signed(28742, LUT_AMPL_WIDTH),
		21609 => to_signed(28741, LUT_AMPL_WIDTH),
		21610 => to_signed(28739, LUT_AMPL_WIDTH),
		21611 => to_signed(28738, LUT_AMPL_WIDTH),
		21612 => to_signed(28736, LUT_AMPL_WIDTH),
		21613 => to_signed(28735, LUT_AMPL_WIDTH),
		21614 => to_signed(28733, LUT_AMPL_WIDTH),
		21615 => to_signed(28732, LUT_AMPL_WIDTH),
		21616 => to_signed(28730, LUT_AMPL_WIDTH),
		21617 => to_signed(28729, LUT_AMPL_WIDTH),
		21618 => to_signed(28727, LUT_AMPL_WIDTH),
		21619 => to_signed(28726, LUT_AMPL_WIDTH),
		21620 => to_signed(28724, LUT_AMPL_WIDTH),
		21621 => to_signed(28723, LUT_AMPL_WIDTH),
		21622 => to_signed(28721, LUT_AMPL_WIDTH),
		21623 => to_signed(28720, LUT_AMPL_WIDTH),
		21624 => to_signed(28718, LUT_AMPL_WIDTH),
		21625 => to_signed(28717, LUT_AMPL_WIDTH),
		21626 => to_signed(28715, LUT_AMPL_WIDTH),
		21627 => to_signed(28714, LUT_AMPL_WIDTH),
		21628 => to_signed(28712, LUT_AMPL_WIDTH),
		21629 => to_signed(28711, LUT_AMPL_WIDTH),
		21630 => to_signed(28709, LUT_AMPL_WIDTH),
		21631 => to_signed(28708, LUT_AMPL_WIDTH),
		21632 => to_signed(28706, LUT_AMPL_WIDTH),
		21633 => to_signed(28705, LUT_AMPL_WIDTH),
		21634 => to_signed(28703, LUT_AMPL_WIDTH),
		21635 => to_signed(28702, LUT_AMPL_WIDTH),
		21636 => to_signed(28700, LUT_AMPL_WIDTH),
		21637 => to_signed(28699, LUT_AMPL_WIDTH),
		21638 => to_signed(28697, LUT_AMPL_WIDTH),
		21639 => to_signed(28696, LUT_AMPL_WIDTH),
		21640 => to_signed(28694, LUT_AMPL_WIDTH),
		21641 => to_signed(28693, LUT_AMPL_WIDTH),
		21642 => to_signed(28691, LUT_AMPL_WIDTH),
		21643 => to_signed(28690, LUT_AMPL_WIDTH),
		21644 => to_signed(28688, LUT_AMPL_WIDTH),
		21645 => to_signed(28686, LUT_AMPL_WIDTH),
		21646 => to_signed(28685, LUT_AMPL_WIDTH),
		21647 => to_signed(28683, LUT_AMPL_WIDTH),
		21648 => to_signed(28682, LUT_AMPL_WIDTH),
		21649 => to_signed(28680, LUT_AMPL_WIDTH),
		21650 => to_signed(28679, LUT_AMPL_WIDTH),
		21651 => to_signed(28677, LUT_AMPL_WIDTH),
		21652 => to_signed(28676, LUT_AMPL_WIDTH),
		21653 => to_signed(28674, LUT_AMPL_WIDTH),
		21654 => to_signed(28673, LUT_AMPL_WIDTH),
		21655 => to_signed(28671, LUT_AMPL_WIDTH),
		21656 => to_signed(28670, LUT_AMPL_WIDTH),
		21657 => to_signed(28668, LUT_AMPL_WIDTH),
		21658 => to_signed(28667, LUT_AMPL_WIDTH),
		21659 => to_signed(28665, LUT_AMPL_WIDTH),
		21660 => to_signed(28664, LUT_AMPL_WIDTH),
		21661 => to_signed(28662, LUT_AMPL_WIDTH),
		21662 => to_signed(28661, LUT_AMPL_WIDTH),
		21663 => to_signed(28659, LUT_AMPL_WIDTH),
		21664 => to_signed(28658, LUT_AMPL_WIDTH),
		21665 => to_signed(28656, LUT_AMPL_WIDTH),
		21666 => to_signed(28655, LUT_AMPL_WIDTH),
		21667 => to_signed(28653, LUT_AMPL_WIDTH),
		21668 => to_signed(28651, LUT_AMPL_WIDTH),
		21669 => to_signed(28650, LUT_AMPL_WIDTH),
		21670 => to_signed(28648, LUT_AMPL_WIDTH),
		21671 => to_signed(28647, LUT_AMPL_WIDTH),
		21672 => to_signed(28645, LUT_AMPL_WIDTH),
		21673 => to_signed(28644, LUT_AMPL_WIDTH),
		21674 => to_signed(28642, LUT_AMPL_WIDTH),
		21675 => to_signed(28641, LUT_AMPL_WIDTH),
		21676 => to_signed(28639, LUT_AMPL_WIDTH),
		21677 => to_signed(28638, LUT_AMPL_WIDTH),
		21678 => to_signed(28636, LUT_AMPL_WIDTH),
		21679 => to_signed(28635, LUT_AMPL_WIDTH),
		21680 => to_signed(28633, LUT_AMPL_WIDTH),
		21681 => to_signed(28632, LUT_AMPL_WIDTH),
		21682 => to_signed(28630, LUT_AMPL_WIDTH),
		21683 => to_signed(28629, LUT_AMPL_WIDTH),
		21684 => to_signed(28627, LUT_AMPL_WIDTH),
		21685 => to_signed(28626, LUT_AMPL_WIDTH),
		21686 => to_signed(28624, LUT_AMPL_WIDTH),
		21687 => to_signed(28622, LUT_AMPL_WIDTH),
		21688 => to_signed(28621, LUT_AMPL_WIDTH),
		21689 => to_signed(28619, LUT_AMPL_WIDTH),
		21690 => to_signed(28618, LUT_AMPL_WIDTH),
		21691 => to_signed(28616, LUT_AMPL_WIDTH),
		21692 => to_signed(28615, LUT_AMPL_WIDTH),
		21693 => to_signed(28613, LUT_AMPL_WIDTH),
		21694 => to_signed(28612, LUT_AMPL_WIDTH),
		21695 => to_signed(28610, LUT_AMPL_WIDTH),
		21696 => to_signed(28609, LUT_AMPL_WIDTH),
		21697 => to_signed(28607, LUT_AMPL_WIDTH),
		21698 => to_signed(28606, LUT_AMPL_WIDTH),
		21699 => to_signed(28604, LUT_AMPL_WIDTH),
		21700 => to_signed(28603, LUT_AMPL_WIDTH),
		21701 => to_signed(28601, LUT_AMPL_WIDTH),
		21702 => to_signed(28600, LUT_AMPL_WIDTH),
		21703 => to_signed(28598, LUT_AMPL_WIDTH),
		21704 => to_signed(28596, LUT_AMPL_WIDTH),
		21705 => to_signed(28595, LUT_AMPL_WIDTH),
		21706 => to_signed(28593, LUT_AMPL_WIDTH),
		21707 => to_signed(28592, LUT_AMPL_WIDTH),
		21708 => to_signed(28590, LUT_AMPL_WIDTH),
		21709 => to_signed(28589, LUT_AMPL_WIDTH),
		21710 => to_signed(28587, LUT_AMPL_WIDTH),
		21711 => to_signed(28586, LUT_AMPL_WIDTH),
		21712 => to_signed(28584, LUT_AMPL_WIDTH),
		21713 => to_signed(28583, LUT_AMPL_WIDTH),
		21714 => to_signed(28581, LUT_AMPL_WIDTH),
		21715 => to_signed(28580, LUT_AMPL_WIDTH),
		21716 => to_signed(28578, LUT_AMPL_WIDTH),
		21717 => to_signed(28576, LUT_AMPL_WIDTH),
		21718 => to_signed(28575, LUT_AMPL_WIDTH),
		21719 => to_signed(28573, LUT_AMPL_WIDTH),
		21720 => to_signed(28572, LUT_AMPL_WIDTH),
		21721 => to_signed(28570, LUT_AMPL_WIDTH),
		21722 => to_signed(28569, LUT_AMPL_WIDTH),
		21723 => to_signed(28567, LUT_AMPL_WIDTH),
		21724 => to_signed(28566, LUT_AMPL_WIDTH),
		21725 => to_signed(28564, LUT_AMPL_WIDTH),
		21726 => to_signed(28563, LUT_AMPL_WIDTH),
		21727 => to_signed(28561, LUT_AMPL_WIDTH),
		21728 => to_signed(28560, LUT_AMPL_WIDTH),
		21729 => to_signed(28558, LUT_AMPL_WIDTH),
		21730 => to_signed(28556, LUT_AMPL_WIDTH),
		21731 => to_signed(28555, LUT_AMPL_WIDTH),
		21732 => to_signed(28553, LUT_AMPL_WIDTH),
		21733 => to_signed(28552, LUT_AMPL_WIDTH),
		21734 => to_signed(28550, LUT_AMPL_WIDTH),
		21735 => to_signed(28549, LUT_AMPL_WIDTH),
		21736 => to_signed(28547, LUT_AMPL_WIDTH),
		21737 => to_signed(28546, LUT_AMPL_WIDTH),
		21738 => to_signed(28544, LUT_AMPL_WIDTH),
		21739 => to_signed(28543, LUT_AMPL_WIDTH),
		21740 => to_signed(28541, LUT_AMPL_WIDTH),
		21741 => to_signed(28540, LUT_AMPL_WIDTH),
		21742 => to_signed(28538, LUT_AMPL_WIDTH),
		21743 => to_signed(28536, LUT_AMPL_WIDTH),
		21744 => to_signed(28535, LUT_AMPL_WIDTH),
		21745 => to_signed(28533, LUT_AMPL_WIDTH),
		21746 => to_signed(28532, LUT_AMPL_WIDTH),
		21747 => to_signed(28530, LUT_AMPL_WIDTH),
		21748 => to_signed(28529, LUT_AMPL_WIDTH),
		21749 => to_signed(28527, LUT_AMPL_WIDTH),
		21750 => to_signed(28526, LUT_AMPL_WIDTH),
		21751 => to_signed(28524, LUT_AMPL_WIDTH),
		21752 => to_signed(28523, LUT_AMPL_WIDTH),
		21753 => to_signed(28521, LUT_AMPL_WIDTH),
		21754 => to_signed(28519, LUT_AMPL_WIDTH),
		21755 => to_signed(28518, LUT_AMPL_WIDTH),
		21756 => to_signed(28516, LUT_AMPL_WIDTH),
		21757 => to_signed(28515, LUT_AMPL_WIDTH),
		21758 => to_signed(28513, LUT_AMPL_WIDTH),
		21759 => to_signed(28512, LUT_AMPL_WIDTH),
		21760 => to_signed(28510, LUT_AMPL_WIDTH),
		21761 => to_signed(28509, LUT_AMPL_WIDTH),
		21762 => to_signed(28507, LUT_AMPL_WIDTH),
		21763 => to_signed(28505, LUT_AMPL_WIDTH),
		21764 => to_signed(28504, LUT_AMPL_WIDTH),
		21765 => to_signed(28502, LUT_AMPL_WIDTH),
		21766 => to_signed(28501, LUT_AMPL_WIDTH),
		21767 => to_signed(28499, LUT_AMPL_WIDTH),
		21768 => to_signed(28498, LUT_AMPL_WIDTH),
		21769 => to_signed(28496, LUT_AMPL_WIDTH),
		21770 => to_signed(28495, LUT_AMPL_WIDTH),
		21771 => to_signed(28493, LUT_AMPL_WIDTH),
		21772 => to_signed(28492, LUT_AMPL_WIDTH),
		21773 => to_signed(28490, LUT_AMPL_WIDTH),
		21774 => to_signed(28488, LUT_AMPL_WIDTH),
		21775 => to_signed(28487, LUT_AMPL_WIDTH),
		21776 => to_signed(28485, LUT_AMPL_WIDTH),
		21777 => to_signed(28484, LUT_AMPL_WIDTH),
		21778 => to_signed(28482, LUT_AMPL_WIDTH),
		21779 => to_signed(28481, LUT_AMPL_WIDTH),
		21780 => to_signed(28479, LUT_AMPL_WIDTH),
		21781 => to_signed(28478, LUT_AMPL_WIDTH),
		21782 => to_signed(28476, LUT_AMPL_WIDTH),
		21783 => to_signed(28474, LUT_AMPL_WIDTH),
		21784 => to_signed(28473, LUT_AMPL_WIDTH),
		21785 => to_signed(28471, LUT_AMPL_WIDTH),
		21786 => to_signed(28470, LUT_AMPL_WIDTH),
		21787 => to_signed(28468, LUT_AMPL_WIDTH),
		21788 => to_signed(28467, LUT_AMPL_WIDTH),
		21789 => to_signed(28465, LUT_AMPL_WIDTH),
		21790 => to_signed(28464, LUT_AMPL_WIDTH),
		21791 => to_signed(28462, LUT_AMPL_WIDTH),
		21792 => to_signed(28460, LUT_AMPL_WIDTH),
		21793 => to_signed(28459, LUT_AMPL_WIDTH),
		21794 => to_signed(28457, LUT_AMPL_WIDTH),
		21795 => to_signed(28456, LUT_AMPL_WIDTH),
		21796 => to_signed(28454, LUT_AMPL_WIDTH),
		21797 => to_signed(28453, LUT_AMPL_WIDTH),
		21798 => to_signed(28451, LUT_AMPL_WIDTH),
		21799 => to_signed(28450, LUT_AMPL_WIDTH),
		21800 => to_signed(28448, LUT_AMPL_WIDTH),
		21801 => to_signed(28446, LUT_AMPL_WIDTH),
		21802 => to_signed(28445, LUT_AMPL_WIDTH),
		21803 => to_signed(28443, LUT_AMPL_WIDTH),
		21804 => to_signed(28442, LUT_AMPL_WIDTH),
		21805 => to_signed(28440, LUT_AMPL_WIDTH),
		21806 => to_signed(28439, LUT_AMPL_WIDTH),
		21807 => to_signed(28437, LUT_AMPL_WIDTH),
		21808 => to_signed(28436, LUT_AMPL_WIDTH),
		21809 => to_signed(28434, LUT_AMPL_WIDTH),
		21810 => to_signed(28432, LUT_AMPL_WIDTH),
		21811 => to_signed(28431, LUT_AMPL_WIDTH),
		21812 => to_signed(28429, LUT_AMPL_WIDTH),
		21813 => to_signed(28428, LUT_AMPL_WIDTH),
		21814 => to_signed(28426, LUT_AMPL_WIDTH),
		21815 => to_signed(28425, LUT_AMPL_WIDTH),
		21816 => to_signed(28423, LUT_AMPL_WIDTH),
		21817 => to_signed(28421, LUT_AMPL_WIDTH),
		21818 => to_signed(28420, LUT_AMPL_WIDTH),
		21819 => to_signed(28418, LUT_AMPL_WIDTH),
		21820 => to_signed(28417, LUT_AMPL_WIDTH),
		21821 => to_signed(28415, LUT_AMPL_WIDTH),
		21822 => to_signed(28414, LUT_AMPL_WIDTH),
		21823 => to_signed(28412, LUT_AMPL_WIDTH),
		21824 => to_signed(28411, LUT_AMPL_WIDTH),
		21825 => to_signed(28409, LUT_AMPL_WIDTH),
		21826 => to_signed(28407, LUT_AMPL_WIDTH),
		21827 => to_signed(28406, LUT_AMPL_WIDTH),
		21828 => to_signed(28404, LUT_AMPL_WIDTH),
		21829 => to_signed(28403, LUT_AMPL_WIDTH),
		21830 => to_signed(28401, LUT_AMPL_WIDTH),
		21831 => to_signed(28400, LUT_AMPL_WIDTH),
		21832 => to_signed(28398, LUT_AMPL_WIDTH),
		21833 => to_signed(28396, LUT_AMPL_WIDTH),
		21834 => to_signed(28395, LUT_AMPL_WIDTH),
		21835 => to_signed(28393, LUT_AMPL_WIDTH),
		21836 => to_signed(28392, LUT_AMPL_WIDTH),
		21837 => to_signed(28390, LUT_AMPL_WIDTH),
		21838 => to_signed(28389, LUT_AMPL_WIDTH),
		21839 => to_signed(28387, LUT_AMPL_WIDTH),
		21840 => to_signed(28385, LUT_AMPL_WIDTH),
		21841 => to_signed(28384, LUT_AMPL_WIDTH),
		21842 => to_signed(28382, LUT_AMPL_WIDTH),
		21843 => to_signed(28381, LUT_AMPL_WIDTH),
		21844 => to_signed(28379, LUT_AMPL_WIDTH),
		21845 => to_signed(28378, LUT_AMPL_WIDTH),
		21846 => to_signed(28376, LUT_AMPL_WIDTH),
		21847 => to_signed(28374, LUT_AMPL_WIDTH),
		21848 => to_signed(28373, LUT_AMPL_WIDTH),
		21849 => to_signed(28371, LUT_AMPL_WIDTH),
		21850 => to_signed(28370, LUT_AMPL_WIDTH),
		21851 => to_signed(28368, LUT_AMPL_WIDTH),
		21852 => to_signed(28367, LUT_AMPL_WIDTH),
		21853 => to_signed(28365, LUT_AMPL_WIDTH),
		21854 => to_signed(28363, LUT_AMPL_WIDTH),
		21855 => to_signed(28362, LUT_AMPL_WIDTH),
		21856 => to_signed(28360, LUT_AMPL_WIDTH),
		21857 => to_signed(28359, LUT_AMPL_WIDTH),
		21858 => to_signed(28357, LUT_AMPL_WIDTH),
		21859 => to_signed(28356, LUT_AMPL_WIDTH),
		21860 => to_signed(28354, LUT_AMPL_WIDTH),
		21861 => to_signed(28352, LUT_AMPL_WIDTH),
		21862 => to_signed(28351, LUT_AMPL_WIDTH),
		21863 => to_signed(28349, LUT_AMPL_WIDTH),
		21864 => to_signed(28348, LUT_AMPL_WIDTH),
		21865 => to_signed(28346, LUT_AMPL_WIDTH),
		21866 => to_signed(28345, LUT_AMPL_WIDTH),
		21867 => to_signed(28343, LUT_AMPL_WIDTH),
		21868 => to_signed(28341, LUT_AMPL_WIDTH),
		21869 => to_signed(28340, LUT_AMPL_WIDTH),
		21870 => to_signed(28338, LUT_AMPL_WIDTH),
		21871 => to_signed(28337, LUT_AMPL_WIDTH),
		21872 => to_signed(28335, LUT_AMPL_WIDTH),
		21873 => to_signed(28333, LUT_AMPL_WIDTH),
		21874 => to_signed(28332, LUT_AMPL_WIDTH),
		21875 => to_signed(28330, LUT_AMPL_WIDTH),
		21876 => to_signed(28329, LUT_AMPL_WIDTH),
		21877 => to_signed(28327, LUT_AMPL_WIDTH),
		21878 => to_signed(28326, LUT_AMPL_WIDTH),
		21879 => to_signed(28324, LUT_AMPL_WIDTH),
		21880 => to_signed(28322, LUT_AMPL_WIDTH),
		21881 => to_signed(28321, LUT_AMPL_WIDTH),
		21882 => to_signed(28319, LUT_AMPL_WIDTH),
		21883 => to_signed(28318, LUT_AMPL_WIDTH),
		21884 => to_signed(28316, LUT_AMPL_WIDTH),
		21885 => to_signed(28315, LUT_AMPL_WIDTH),
		21886 => to_signed(28313, LUT_AMPL_WIDTH),
		21887 => to_signed(28311, LUT_AMPL_WIDTH),
		21888 => to_signed(28310, LUT_AMPL_WIDTH),
		21889 => to_signed(28308, LUT_AMPL_WIDTH),
		21890 => to_signed(28307, LUT_AMPL_WIDTH),
		21891 => to_signed(28305, LUT_AMPL_WIDTH),
		21892 => to_signed(28303, LUT_AMPL_WIDTH),
		21893 => to_signed(28302, LUT_AMPL_WIDTH),
		21894 => to_signed(28300, LUT_AMPL_WIDTH),
		21895 => to_signed(28299, LUT_AMPL_WIDTH),
		21896 => to_signed(28297, LUT_AMPL_WIDTH),
		21897 => to_signed(28296, LUT_AMPL_WIDTH),
		21898 => to_signed(28294, LUT_AMPL_WIDTH),
		21899 => to_signed(28292, LUT_AMPL_WIDTH),
		21900 => to_signed(28291, LUT_AMPL_WIDTH),
		21901 => to_signed(28289, LUT_AMPL_WIDTH),
		21902 => to_signed(28288, LUT_AMPL_WIDTH),
		21903 => to_signed(28286, LUT_AMPL_WIDTH),
		21904 => to_signed(28284, LUT_AMPL_WIDTH),
		21905 => to_signed(28283, LUT_AMPL_WIDTH),
		21906 => to_signed(28281, LUT_AMPL_WIDTH),
		21907 => to_signed(28280, LUT_AMPL_WIDTH),
		21908 => to_signed(28278, LUT_AMPL_WIDTH),
		21909 => to_signed(28277, LUT_AMPL_WIDTH),
		21910 => to_signed(28275, LUT_AMPL_WIDTH),
		21911 => to_signed(28273, LUT_AMPL_WIDTH),
		21912 => to_signed(28272, LUT_AMPL_WIDTH),
		21913 => to_signed(28270, LUT_AMPL_WIDTH),
		21914 => to_signed(28269, LUT_AMPL_WIDTH),
		21915 => to_signed(28267, LUT_AMPL_WIDTH),
		21916 => to_signed(28265, LUT_AMPL_WIDTH),
		21917 => to_signed(28264, LUT_AMPL_WIDTH),
		21918 => to_signed(28262, LUT_AMPL_WIDTH),
		21919 => to_signed(28261, LUT_AMPL_WIDTH),
		21920 => to_signed(28259, LUT_AMPL_WIDTH),
		21921 => to_signed(28257, LUT_AMPL_WIDTH),
		21922 => to_signed(28256, LUT_AMPL_WIDTH),
		21923 => to_signed(28254, LUT_AMPL_WIDTH),
		21924 => to_signed(28253, LUT_AMPL_WIDTH),
		21925 => to_signed(28251, LUT_AMPL_WIDTH),
		21926 => to_signed(28249, LUT_AMPL_WIDTH),
		21927 => to_signed(28248, LUT_AMPL_WIDTH),
		21928 => to_signed(28246, LUT_AMPL_WIDTH),
		21929 => to_signed(28245, LUT_AMPL_WIDTH),
		21930 => to_signed(28243, LUT_AMPL_WIDTH),
		21931 => to_signed(28242, LUT_AMPL_WIDTH),
		21932 => to_signed(28240, LUT_AMPL_WIDTH),
		21933 => to_signed(28238, LUT_AMPL_WIDTH),
		21934 => to_signed(28237, LUT_AMPL_WIDTH),
		21935 => to_signed(28235, LUT_AMPL_WIDTH),
		21936 => to_signed(28234, LUT_AMPL_WIDTH),
		21937 => to_signed(28232, LUT_AMPL_WIDTH),
		21938 => to_signed(28230, LUT_AMPL_WIDTH),
		21939 => to_signed(28229, LUT_AMPL_WIDTH),
		21940 => to_signed(28227, LUT_AMPL_WIDTH),
		21941 => to_signed(28226, LUT_AMPL_WIDTH),
		21942 => to_signed(28224, LUT_AMPL_WIDTH),
		21943 => to_signed(28222, LUT_AMPL_WIDTH),
		21944 => to_signed(28221, LUT_AMPL_WIDTH),
		21945 => to_signed(28219, LUT_AMPL_WIDTH),
		21946 => to_signed(28218, LUT_AMPL_WIDTH),
		21947 => to_signed(28216, LUT_AMPL_WIDTH),
		21948 => to_signed(28214, LUT_AMPL_WIDTH),
		21949 => to_signed(28213, LUT_AMPL_WIDTH),
		21950 => to_signed(28211, LUT_AMPL_WIDTH),
		21951 => to_signed(28210, LUT_AMPL_WIDTH),
		21952 => to_signed(28208, LUT_AMPL_WIDTH),
		21953 => to_signed(28206, LUT_AMPL_WIDTH),
		21954 => to_signed(28205, LUT_AMPL_WIDTH),
		21955 => to_signed(28203, LUT_AMPL_WIDTH),
		21956 => to_signed(28202, LUT_AMPL_WIDTH),
		21957 => to_signed(28200, LUT_AMPL_WIDTH),
		21958 => to_signed(28198, LUT_AMPL_WIDTH),
		21959 => to_signed(28197, LUT_AMPL_WIDTH),
		21960 => to_signed(28195, LUT_AMPL_WIDTH),
		21961 => to_signed(28194, LUT_AMPL_WIDTH),
		21962 => to_signed(28192, LUT_AMPL_WIDTH),
		21963 => to_signed(28190, LUT_AMPL_WIDTH),
		21964 => to_signed(28189, LUT_AMPL_WIDTH),
		21965 => to_signed(28187, LUT_AMPL_WIDTH),
		21966 => to_signed(28186, LUT_AMPL_WIDTH),
		21967 => to_signed(28184, LUT_AMPL_WIDTH),
		21968 => to_signed(28182, LUT_AMPL_WIDTH),
		21969 => to_signed(28181, LUT_AMPL_WIDTH),
		21970 => to_signed(28179, LUT_AMPL_WIDTH),
		21971 => to_signed(28178, LUT_AMPL_WIDTH),
		21972 => to_signed(28176, LUT_AMPL_WIDTH),
		21973 => to_signed(28174, LUT_AMPL_WIDTH),
		21974 => to_signed(28173, LUT_AMPL_WIDTH),
		21975 => to_signed(28171, LUT_AMPL_WIDTH),
		21976 => to_signed(28170, LUT_AMPL_WIDTH),
		21977 => to_signed(28168, LUT_AMPL_WIDTH),
		21978 => to_signed(28166, LUT_AMPL_WIDTH),
		21979 => to_signed(28165, LUT_AMPL_WIDTH),
		21980 => to_signed(28163, LUT_AMPL_WIDTH),
		21981 => to_signed(28162, LUT_AMPL_WIDTH),
		21982 => to_signed(28160, LUT_AMPL_WIDTH),
		21983 => to_signed(28158, LUT_AMPL_WIDTH),
		21984 => to_signed(28157, LUT_AMPL_WIDTH),
		21985 => to_signed(28155, LUT_AMPL_WIDTH),
		21986 => to_signed(28154, LUT_AMPL_WIDTH),
		21987 => to_signed(28152, LUT_AMPL_WIDTH),
		21988 => to_signed(28150, LUT_AMPL_WIDTH),
		21989 => to_signed(28149, LUT_AMPL_WIDTH),
		21990 => to_signed(28147, LUT_AMPL_WIDTH),
		21991 => to_signed(28145, LUT_AMPL_WIDTH),
		21992 => to_signed(28144, LUT_AMPL_WIDTH),
		21993 => to_signed(28142, LUT_AMPL_WIDTH),
		21994 => to_signed(28141, LUT_AMPL_WIDTH),
		21995 => to_signed(28139, LUT_AMPL_WIDTH),
		21996 => to_signed(28137, LUT_AMPL_WIDTH),
		21997 => to_signed(28136, LUT_AMPL_WIDTH),
		21998 => to_signed(28134, LUT_AMPL_WIDTH),
		21999 => to_signed(28133, LUT_AMPL_WIDTH),
		22000 => to_signed(28131, LUT_AMPL_WIDTH),
		22001 => to_signed(28129, LUT_AMPL_WIDTH),
		22002 => to_signed(28128, LUT_AMPL_WIDTH),
		22003 => to_signed(28126, LUT_AMPL_WIDTH),
		22004 => to_signed(28125, LUT_AMPL_WIDTH),
		22005 => to_signed(28123, LUT_AMPL_WIDTH),
		22006 => to_signed(28121, LUT_AMPL_WIDTH),
		22007 => to_signed(28120, LUT_AMPL_WIDTH),
		22008 => to_signed(28118, LUT_AMPL_WIDTH),
		22009 => to_signed(28116, LUT_AMPL_WIDTH),
		22010 => to_signed(28115, LUT_AMPL_WIDTH),
		22011 => to_signed(28113, LUT_AMPL_WIDTH),
		22012 => to_signed(28112, LUT_AMPL_WIDTH),
		22013 => to_signed(28110, LUT_AMPL_WIDTH),
		22014 => to_signed(28108, LUT_AMPL_WIDTH),
		22015 => to_signed(28107, LUT_AMPL_WIDTH),
		22016 => to_signed(28105, LUT_AMPL_WIDTH),
		22017 => to_signed(28104, LUT_AMPL_WIDTH),
		22018 => to_signed(28102, LUT_AMPL_WIDTH),
		22019 => to_signed(28100, LUT_AMPL_WIDTH),
		22020 => to_signed(28099, LUT_AMPL_WIDTH),
		22021 => to_signed(28097, LUT_AMPL_WIDTH),
		22022 => to_signed(28095, LUT_AMPL_WIDTH),
		22023 => to_signed(28094, LUT_AMPL_WIDTH),
		22024 => to_signed(28092, LUT_AMPL_WIDTH),
		22025 => to_signed(28091, LUT_AMPL_WIDTH),
		22026 => to_signed(28089, LUT_AMPL_WIDTH),
		22027 => to_signed(28087, LUT_AMPL_WIDTH),
		22028 => to_signed(28086, LUT_AMPL_WIDTH),
		22029 => to_signed(28084, LUT_AMPL_WIDTH),
		22030 => to_signed(28083, LUT_AMPL_WIDTH),
		22031 => to_signed(28081, LUT_AMPL_WIDTH),
		22032 => to_signed(28079, LUT_AMPL_WIDTH),
		22033 => to_signed(28078, LUT_AMPL_WIDTH),
		22034 => to_signed(28076, LUT_AMPL_WIDTH),
		22035 => to_signed(28074, LUT_AMPL_WIDTH),
		22036 => to_signed(28073, LUT_AMPL_WIDTH),
		22037 => to_signed(28071, LUT_AMPL_WIDTH),
		22038 => to_signed(28070, LUT_AMPL_WIDTH),
		22039 => to_signed(28068, LUT_AMPL_WIDTH),
		22040 => to_signed(28066, LUT_AMPL_WIDTH),
		22041 => to_signed(28065, LUT_AMPL_WIDTH),
		22042 => to_signed(28063, LUT_AMPL_WIDTH),
		22043 => to_signed(28061, LUT_AMPL_WIDTH),
		22044 => to_signed(28060, LUT_AMPL_WIDTH),
		22045 => to_signed(28058, LUT_AMPL_WIDTH),
		22046 => to_signed(28057, LUT_AMPL_WIDTH),
		22047 => to_signed(28055, LUT_AMPL_WIDTH),
		22048 => to_signed(28053, LUT_AMPL_WIDTH),
		22049 => to_signed(28052, LUT_AMPL_WIDTH),
		22050 => to_signed(28050, LUT_AMPL_WIDTH),
		22051 => to_signed(28049, LUT_AMPL_WIDTH),
		22052 => to_signed(28047, LUT_AMPL_WIDTH),
		22053 => to_signed(28045, LUT_AMPL_WIDTH),
		22054 => to_signed(28044, LUT_AMPL_WIDTH),
		22055 => to_signed(28042, LUT_AMPL_WIDTH),
		22056 => to_signed(28040, LUT_AMPL_WIDTH),
		22057 => to_signed(28039, LUT_AMPL_WIDTH),
		22058 => to_signed(28037, LUT_AMPL_WIDTH),
		22059 => to_signed(28036, LUT_AMPL_WIDTH),
		22060 => to_signed(28034, LUT_AMPL_WIDTH),
		22061 => to_signed(28032, LUT_AMPL_WIDTH),
		22062 => to_signed(28031, LUT_AMPL_WIDTH),
		22063 => to_signed(28029, LUT_AMPL_WIDTH),
		22064 => to_signed(28027, LUT_AMPL_WIDTH),
		22065 => to_signed(28026, LUT_AMPL_WIDTH),
		22066 => to_signed(28024, LUT_AMPL_WIDTH),
		22067 => to_signed(28022, LUT_AMPL_WIDTH),
		22068 => to_signed(28021, LUT_AMPL_WIDTH),
		22069 => to_signed(28019, LUT_AMPL_WIDTH),
		22070 => to_signed(28018, LUT_AMPL_WIDTH),
		22071 => to_signed(28016, LUT_AMPL_WIDTH),
		22072 => to_signed(28014, LUT_AMPL_WIDTH),
		22073 => to_signed(28013, LUT_AMPL_WIDTH),
		22074 => to_signed(28011, LUT_AMPL_WIDTH),
		22075 => to_signed(28009, LUT_AMPL_WIDTH),
		22076 => to_signed(28008, LUT_AMPL_WIDTH),
		22077 => to_signed(28006, LUT_AMPL_WIDTH),
		22078 => to_signed(28005, LUT_AMPL_WIDTH),
		22079 => to_signed(28003, LUT_AMPL_WIDTH),
		22080 => to_signed(28001, LUT_AMPL_WIDTH),
		22081 => to_signed(28000, LUT_AMPL_WIDTH),
		22082 => to_signed(27998, LUT_AMPL_WIDTH),
		22083 => to_signed(27996, LUT_AMPL_WIDTH),
		22084 => to_signed(27995, LUT_AMPL_WIDTH),
		22085 => to_signed(27993, LUT_AMPL_WIDTH),
		22086 => to_signed(27992, LUT_AMPL_WIDTH),
		22087 => to_signed(27990, LUT_AMPL_WIDTH),
		22088 => to_signed(27988, LUT_AMPL_WIDTH),
		22089 => to_signed(27987, LUT_AMPL_WIDTH),
		22090 => to_signed(27985, LUT_AMPL_WIDTH),
		22091 => to_signed(27983, LUT_AMPL_WIDTH),
		22092 => to_signed(27982, LUT_AMPL_WIDTH),
		22093 => to_signed(27980, LUT_AMPL_WIDTH),
		22094 => to_signed(27978, LUT_AMPL_WIDTH),
		22095 => to_signed(27977, LUT_AMPL_WIDTH),
		22096 => to_signed(27975, LUT_AMPL_WIDTH),
		22097 => to_signed(27974, LUT_AMPL_WIDTH),
		22098 => to_signed(27972, LUT_AMPL_WIDTH),
		22099 => to_signed(27970, LUT_AMPL_WIDTH),
		22100 => to_signed(27969, LUT_AMPL_WIDTH),
		22101 => to_signed(27967, LUT_AMPL_WIDTH),
		22102 => to_signed(27965, LUT_AMPL_WIDTH),
		22103 => to_signed(27964, LUT_AMPL_WIDTH),
		22104 => to_signed(27962, LUT_AMPL_WIDTH),
		22105 => to_signed(27960, LUT_AMPL_WIDTH),
		22106 => to_signed(27959, LUT_AMPL_WIDTH),
		22107 => to_signed(27957, LUT_AMPL_WIDTH),
		22108 => to_signed(27956, LUT_AMPL_WIDTH),
		22109 => to_signed(27954, LUT_AMPL_WIDTH),
		22110 => to_signed(27952, LUT_AMPL_WIDTH),
		22111 => to_signed(27951, LUT_AMPL_WIDTH),
		22112 => to_signed(27949, LUT_AMPL_WIDTH),
		22113 => to_signed(27947, LUT_AMPL_WIDTH),
		22114 => to_signed(27946, LUT_AMPL_WIDTH),
		22115 => to_signed(27944, LUT_AMPL_WIDTH),
		22116 => to_signed(27942, LUT_AMPL_WIDTH),
		22117 => to_signed(27941, LUT_AMPL_WIDTH),
		22118 => to_signed(27939, LUT_AMPL_WIDTH),
		22119 => to_signed(27937, LUT_AMPL_WIDTH),
		22120 => to_signed(27936, LUT_AMPL_WIDTH),
		22121 => to_signed(27934, LUT_AMPL_WIDTH),
		22122 => to_signed(27933, LUT_AMPL_WIDTH),
		22123 => to_signed(27931, LUT_AMPL_WIDTH),
		22124 => to_signed(27929, LUT_AMPL_WIDTH),
		22125 => to_signed(27928, LUT_AMPL_WIDTH),
		22126 => to_signed(27926, LUT_AMPL_WIDTH),
		22127 => to_signed(27924, LUT_AMPL_WIDTH),
		22128 => to_signed(27923, LUT_AMPL_WIDTH),
		22129 => to_signed(27921, LUT_AMPL_WIDTH),
		22130 => to_signed(27919, LUT_AMPL_WIDTH),
		22131 => to_signed(27918, LUT_AMPL_WIDTH),
		22132 => to_signed(27916, LUT_AMPL_WIDTH),
		22133 => to_signed(27914, LUT_AMPL_WIDTH),
		22134 => to_signed(27913, LUT_AMPL_WIDTH),
		22135 => to_signed(27911, LUT_AMPL_WIDTH),
		22136 => to_signed(27910, LUT_AMPL_WIDTH),
		22137 => to_signed(27908, LUT_AMPL_WIDTH),
		22138 => to_signed(27906, LUT_AMPL_WIDTH),
		22139 => to_signed(27905, LUT_AMPL_WIDTH),
		22140 => to_signed(27903, LUT_AMPL_WIDTH),
		22141 => to_signed(27901, LUT_AMPL_WIDTH),
		22142 => to_signed(27900, LUT_AMPL_WIDTH),
		22143 => to_signed(27898, LUT_AMPL_WIDTH),
		22144 => to_signed(27896, LUT_AMPL_WIDTH),
		22145 => to_signed(27895, LUT_AMPL_WIDTH),
		22146 => to_signed(27893, LUT_AMPL_WIDTH),
		22147 => to_signed(27891, LUT_AMPL_WIDTH),
		22148 => to_signed(27890, LUT_AMPL_WIDTH),
		22149 => to_signed(27888, LUT_AMPL_WIDTH),
		22150 => to_signed(27886, LUT_AMPL_WIDTH),
		22151 => to_signed(27885, LUT_AMPL_WIDTH),
		22152 => to_signed(27883, LUT_AMPL_WIDTH),
		22153 => to_signed(27882, LUT_AMPL_WIDTH),
		22154 => to_signed(27880, LUT_AMPL_WIDTH),
		22155 => to_signed(27878, LUT_AMPL_WIDTH),
		22156 => to_signed(27877, LUT_AMPL_WIDTH),
		22157 => to_signed(27875, LUT_AMPL_WIDTH),
		22158 => to_signed(27873, LUT_AMPL_WIDTH),
		22159 => to_signed(27872, LUT_AMPL_WIDTH),
		22160 => to_signed(27870, LUT_AMPL_WIDTH),
		22161 => to_signed(27868, LUT_AMPL_WIDTH),
		22162 => to_signed(27867, LUT_AMPL_WIDTH),
		22163 => to_signed(27865, LUT_AMPL_WIDTH),
		22164 => to_signed(27863, LUT_AMPL_WIDTH),
		22165 => to_signed(27862, LUT_AMPL_WIDTH),
		22166 => to_signed(27860, LUT_AMPL_WIDTH),
		22167 => to_signed(27858, LUT_AMPL_WIDTH),
		22168 => to_signed(27857, LUT_AMPL_WIDTH),
		22169 => to_signed(27855, LUT_AMPL_WIDTH),
		22170 => to_signed(27853, LUT_AMPL_WIDTH),
		22171 => to_signed(27852, LUT_AMPL_WIDTH),
		22172 => to_signed(27850, LUT_AMPL_WIDTH),
		22173 => to_signed(27848, LUT_AMPL_WIDTH),
		22174 => to_signed(27847, LUT_AMPL_WIDTH),
		22175 => to_signed(27845, LUT_AMPL_WIDTH),
		22176 => to_signed(27843, LUT_AMPL_WIDTH),
		22177 => to_signed(27842, LUT_AMPL_WIDTH),
		22178 => to_signed(27840, LUT_AMPL_WIDTH),
		22179 => to_signed(27839, LUT_AMPL_WIDTH),
		22180 => to_signed(27837, LUT_AMPL_WIDTH),
		22181 => to_signed(27835, LUT_AMPL_WIDTH),
		22182 => to_signed(27834, LUT_AMPL_WIDTH),
		22183 => to_signed(27832, LUT_AMPL_WIDTH),
		22184 => to_signed(27830, LUT_AMPL_WIDTH),
		22185 => to_signed(27829, LUT_AMPL_WIDTH),
		22186 => to_signed(27827, LUT_AMPL_WIDTH),
		22187 => to_signed(27825, LUT_AMPL_WIDTH),
		22188 => to_signed(27824, LUT_AMPL_WIDTH),
		22189 => to_signed(27822, LUT_AMPL_WIDTH),
		22190 => to_signed(27820, LUT_AMPL_WIDTH),
		22191 => to_signed(27819, LUT_AMPL_WIDTH),
		22192 => to_signed(27817, LUT_AMPL_WIDTH),
		22193 => to_signed(27815, LUT_AMPL_WIDTH),
		22194 => to_signed(27814, LUT_AMPL_WIDTH),
		22195 => to_signed(27812, LUT_AMPL_WIDTH),
		22196 => to_signed(27810, LUT_AMPL_WIDTH),
		22197 => to_signed(27809, LUT_AMPL_WIDTH),
		22198 => to_signed(27807, LUT_AMPL_WIDTH),
		22199 => to_signed(27805, LUT_AMPL_WIDTH),
		22200 => to_signed(27804, LUT_AMPL_WIDTH),
		22201 => to_signed(27802, LUT_AMPL_WIDTH),
		22202 => to_signed(27800, LUT_AMPL_WIDTH),
		22203 => to_signed(27799, LUT_AMPL_WIDTH),
		22204 => to_signed(27797, LUT_AMPL_WIDTH),
		22205 => to_signed(27795, LUT_AMPL_WIDTH),
		22206 => to_signed(27794, LUT_AMPL_WIDTH),
		22207 => to_signed(27792, LUT_AMPL_WIDTH),
		22208 => to_signed(27790, LUT_AMPL_WIDTH),
		22209 => to_signed(27789, LUT_AMPL_WIDTH),
		22210 => to_signed(27787, LUT_AMPL_WIDTH),
		22211 => to_signed(27785, LUT_AMPL_WIDTH),
		22212 => to_signed(27784, LUT_AMPL_WIDTH),
		22213 => to_signed(27782, LUT_AMPL_WIDTH),
		22214 => to_signed(27780, LUT_AMPL_WIDTH),
		22215 => to_signed(27779, LUT_AMPL_WIDTH),
		22216 => to_signed(27777, LUT_AMPL_WIDTH),
		22217 => to_signed(27775, LUT_AMPL_WIDTH),
		22218 => to_signed(27774, LUT_AMPL_WIDTH),
		22219 => to_signed(27772, LUT_AMPL_WIDTH),
		22220 => to_signed(27770, LUT_AMPL_WIDTH),
		22221 => to_signed(27769, LUT_AMPL_WIDTH),
		22222 => to_signed(27767, LUT_AMPL_WIDTH),
		22223 => to_signed(27765, LUT_AMPL_WIDTH),
		22224 => to_signed(27764, LUT_AMPL_WIDTH),
		22225 => to_signed(27762, LUT_AMPL_WIDTH),
		22226 => to_signed(27760, LUT_AMPL_WIDTH),
		22227 => to_signed(27759, LUT_AMPL_WIDTH),
		22228 => to_signed(27757, LUT_AMPL_WIDTH),
		22229 => to_signed(27755, LUT_AMPL_WIDTH),
		22230 => to_signed(27754, LUT_AMPL_WIDTH),
		22231 => to_signed(27752, LUT_AMPL_WIDTH),
		22232 => to_signed(27750, LUT_AMPL_WIDTH),
		22233 => to_signed(27749, LUT_AMPL_WIDTH),
		22234 => to_signed(27747, LUT_AMPL_WIDTH),
		22235 => to_signed(27745, LUT_AMPL_WIDTH),
		22236 => to_signed(27744, LUT_AMPL_WIDTH),
		22237 => to_signed(27742, LUT_AMPL_WIDTH),
		22238 => to_signed(27740, LUT_AMPL_WIDTH),
		22239 => to_signed(27739, LUT_AMPL_WIDTH),
		22240 => to_signed(27737, LUT_AMPL_WIDTH),
		22241 => to_signed(27735, LUT_AMPL_WIDTH),
		22242 => to_signed(27734, LUT_AMPL_WIDTH),
		22243 => to_signed(27732, LUT_AMPL_WIDTH),
		22244 => to_signed(27730, LUT_AMPL_WIDTH),
		22245 => to_signed(27729, LUT_AMPL_WIDTH),
		22246 => to_signed(27727, LUT_AMPL_WIDTH),
		22247 => to_signed(27725, LUT_AMPL_WIDTH),
		22248 => to_signed(27724, LUT_AMPL_WIDTH),
		22249 => to_signed(27722, LUT_AMPL_WIDTH),
		22250 => to_signed(27720, LUT_AMPL_WIDTH),
		22251 => to_signed(27719, LUT_AMPL_WIDTH),
		22252 => to_signed(27717, LUT_AMPL_WIDTH),
		22253 => to_signed(27715, LUT_AMPL_WIDTH),
		22254 => to_signed(27714, LUT_AMPL_WIDTH),
		22255 => to_signed(27712, LUT_AMPL_WIDTH),
		22256 => to_signed(27710, LUT_AMPL_WIDTH),
		22257 => to_signed(27708, LUT_AMPL_WIDTH),
		22258 => to_signed(27707, LUT_AMPL_WIDTH),
		22259 => to_signed(27705, LUT_AMPL_WIDTH),
		22260 => to_signed(27703, LUT_AMPL_WIDTH),
		22261 => to_signed(27702, LUT_AMPL_WIDTH),
		22262 => to_signed(27700, LUT_AMPL_WIDTH),
		22263 => to_signed(27698, LUT_AMPL_WIDTH),
		22264 => to_signed(27697, LUT_AMPL_WIDTH),
		22265 => to_signed(27695, LUT_AMPL_WIDTH),
		22266 => to_signed(27693, LUT_AMPL_WIDTH),
		22267 => to_signed(27692, LUT_AMPL_WIDTH),
		22268 => to_signed(27690, LUT_AMPL_WIDTH),
		22269 => to_signed(27688, LUT_AMPL_WIDTH),
		22270 => to_signed(27687, LUT_AMPL_WIDTH),
		22271 => to_signed(27685, LUT_AMPL_WIDTH),
		22272 => to_signed(27683, LUT_AMPL_WIDTH),
		22273 => to_signed(27682, LUT_AMPL_WIDTH),
		22274 => to_signed(27680, LUT_AMPL_WIDTH),
		22275 => to_signed(27678, LUT_AMPL_WIDTH),
		22276 => to_signed(27677, LUT_AMPL_WIDTH),
		22277 => to_signed(27675, LUT_AMPL_WIDTH),
		22278 => to_signed(27673, LUT_AMPL_WIDTH),
		22279 => to_signed(27672, LUT_AMPL_WIDTH),
		22280 => to_signed(27670, LUT_AMPL_WIDTH),
		22281 => to_signed(27668, LUT_AMPL_WIDTH),
		22282 => to_signed(27666, LUT_AMPL_WIDTH),
		22283 => to_signed(27665, LUT_AMPL_WIDTH),
		22284 => to_signed(27663, LUT_AMPL_WIDTH),
		22285 => to_signed(27661, LUT_AMPL_WIDTH),
		22286 => to_signed(27660, LUT_AMPL_WIDTH),
		22287 => to_signed(27658, LUT_AMPL_WIDTH),
		22288 => to_signed(27656, LUT_AMPL_WIDTH),
		22289 => to_signed(27655, LUT_AMPL_WIDTH),
		22290 => to_signed(27653, LUT_AMPL_WIDTH),
		22291 => to_signed(27651, LUT_AMPL_WIDTH),
		22292 => to_signed(27650, LUT_AMPL_WIDTH),
		22293 => to_signed(27648, LUT_AMPL_WIDTH),
		22294 => to_signed(27646, LUT_AMPL_WIDTH),
		22295 => to_signed(27645, LUT_AMPL_WIDTH),
		22296 => to_signed(27643, LUT_AMPL_WIDTH),
		22297 => to_signed(27641, LUT_AMPL_WIDTH),
		22298 => to_signed(27640, LUT_AMPL_WIDTH),
		22299 => to_signed(27638, LUT_AMPL_WIDTH),
		22300 => to_signed(27636, LUT_AMPL_WIDTH),
		22301 => to_signed(27634, LUT_AMPL_WIDTH),
		22302 => to_signed(27633, LUT_AMPL_WIDTH),
		22303 => to_signed(27631, LUT_AMPL_WIDTH),
		22304 => to_signed(27629, LUT_AMPL_WIDTH),
		22305 => to_signed(27628, LUT_AMPL_WIDTH),
		22306 => to_signed(27626, LUT_AMPL_WIDTH),
		22307 => to_signed(27624, LUT_AMPL_WIDTH),
		22308 => to_signed(27623, LUT_AMPL_WIDTH),
		22309 => to_signed(27621, LUT_AMPL_WIDTH),
		22310 => to_signed(27619, LUT_AMPL_WIDTH),
		22311 => to_signed(27618, LUT_AMPL_WIDTH),
		22312 => to_signed(27616, LUT_AMPL_WIDTH),
		22313 => to_signed(27614, LUT_AMPL_WIDTH),
		22314 => to_signed(27613, LUT_AMPL_WIDTH),
		22315 => to_signed(27611, LUT_AMPL_WIDTH),
		22316 => to_signed(27609, LUT_AMPL_WIDTH),
		22317 => to_signed(27607, LUT_AMPL_WIDTH),
		22318 => to_signed(27606, LUT_AMPL_WIDTH),
		22319 => to_signed(27604, LUT_AMPL_WIDTH),
		22320 => to_signed(27602, LUT_AMPL_WIDTH),
		22321 => to_signed(27601, LUT_AMPL_WIDTH),
		22322 => to_signed(27599, LUT_AMPL_WIDTH),
		22323 => to_signed(27597, LUT_AMPL_WIDTH),
		22324 => to_signed(27596, LUT_AMPL_WIDTH),
		22325 => to_signed(27594, LUT_AMPL_WIDTH),
		22326 => to_signed(27592, LUT_AMPL_WIDTH),
		22327 => to_signed(27590, LUT_AMPL_WIDTH),
		22328 => to_signed(27589, LUT_AMPL_WIDTH),
		22329 => to_signed(27587, LUT_AMPL_WIDTH),
		22330 => to_signed(27585, LUT_AMPL_WIDTH),
		22331 => to_signed(27584, LUT_AMPL_WIDTH),
		22332 => to_signed(27582, LUT_AMPL_WIDTH),
		22333 => to_signed(27580, LUT_AMPL_WIDTH),
		22334 => to_signed(27579, LUT_AMPL_WIDTH),
		22335 => to_signed(27577, LUT_AMPL_WIDTH),
		22336 => to_signed(27575, LUT_AMPL_WIDTH),
		22337 => to_signed(27574, LUT_AMPL_WIDTH),
		22338 => to_signed(27572, LUT_AMPL_WIDTH),
		22339 => to_signed(27570, LUT_AMPL_WIDTH),
		22340 => to_signed(27568, LUT_AMPL_WIDTH),
		22341 => to_signed(27567, LUT_AMPL_WIDTH),
		22342 => to_signed(27565, LUT_AMPL_WIDTH),
		22343 => to_signed(27563, LUT_AMPL_WIDTH),
		22344 => to_signed(27562, LUT_AMPL_WIDTH),
		22345 => to_signed(27560, LUT_AMPL_WIDTH),
		22346 => to_signed(27558, LUT_AMPL_WIDTH),
		22347 => to_signed(27557, LUT_AMPL_WIDTH),
		22348 => to_signed(27555, LUT_AMPL_WIDTH),
		22349 => to_signed(27553, LUT_AMPL_WIDTH),
		22350 => to_signed(27551, LUT_AMPL_WIDTH),
		22351 => to_signed(27550, LUT_AMPL_WIDTH),
		22352 => to_signed(27548, LUT_AMPL_WIDTH),
		22353 => to_signed(27546, LUT_AMPL_WIDTH),
		22354 => to_signed(27545, LUT_AMPL_WIDTH),
		22355 => to_signed(27543, LUT_AMPL_WIDTH),
		22356 => to_signed(27541, LUT_AMPL_WIDTH),
		22357 => to_signed(27540, LUT_AMPL_WIDTH),
		22358 => to_signed(27538, LUT_AMPL_WIDTH),
		22359 => to_signed(27536, LUT_AMPL_WIDTH),
		22360 => to_signed(27534, LUT_AMPL_WIDTH),
		22361 => to_signed(27533, LUT_AMPL_WIDTH),
		22362 => to_signed(27531, LUT_AMPL_WIDTH),
		22363 => to_signed(27529, LUT_AMPL_WIDTH),
		22364 => to_signed(27528, LUT_AMPL_WIDTH),
		22365 => to_signed(27526, LUT_AMPL_WIDTH),
		22366 => to_signed(27524, LUT_AMPL_WIDTH),
		22367 => to_signed(27523, LUT_AMPL_WIDTH),
		22368 => to_signed(27521, LUT_AMPL_WIDTH),
		22369 => to_signed(27519, LUT_AMPL_WIDTH),
		22370 => to_signed(27517, LUT_AMPL_WIDTH),
		22371 => to_signed(27516, LUT_AMPL_WIDTH),
		22372 => to_signed(27514, LUT_AMPL_WIDTH),
		22373 => to_signed(27512, LUT_AMPL_WIDTH),
		22374 => to_signed(27511, LUT_AMPL_WIDTH),
		22375 => to_signed(27509, LUT_AMPL_WIDTH),
		22376 => to_signed(27507, LUT_AMPL_WIDTH),
		22377 => to_signed(27505, LUT_AMPL_WIDTH),
		22378 => to_signed(27504, LUT_AMPL_WIDTH),
		22379 => to_signed(27502, LUT_AMPL_WIDTH),
		22380 => to_signed(27500, LUT_AMPL_WIDTH),
		22381 => to_signed(27499, LUT_AMPL_WIDTH),
		22382 => to_signed(27497, LUT_AMPL_WIDTH),
		22383 => to_signed(27495, LUT_AMPL_WIDTH),
		22384 => to_signed(27493, LUT_AMPL_WIDTH),
		22385 => to_signed(27492, LUT_AMPL_WIDTH),
		22386 => to_signed(27490, LUT_AMPL_WIDTH),
		22387 => to_signed(27488, LUT_AMPL_WIDTH),
		22388 => to_signed(27487, LUT_AMPL_WIDTH),
		22389 => to_signed(27485, LUT_AMPL_WIDTH),
		22390 => to_signed(27483, LUT_AMPL_WIDTH),
		22391 => to_signed(27482, LUT_AMPL_WIDTH),
		22392 => to_signed(27480, LUT_AMPL_WIDTH),
		22393 => to_signed(27478, LUT_AMPL_WIDTH),
		22394 => to_signed(27476, LUT_AMPL_WIDTH),
		22395 => to_signed(27475, LUT_AMPL_WIDTH),
		22396 => to_signed(27473, LUT_AMPL_WIDTH),
		22397 => to_signed(27471, LUT_AMPL_WIDTH),
		22398 => to_signed(27470, LUT_AMPL_WIDTH),
		22399 => to_signed(27468, LUT_AMPL_WIDTH),
		22400 => to_signed(27466, LUT_AMPL_WIDTH),
		22401 => to_signed(27464, LUT_AMPL_WIDTH),
		22402 => to_signed(27463, LUT_AMPL_WIDTH),
		22403 => to_signed(27461, LUT_AMPL_WIDTH),
		22404 => to_signed(27459, LUT_AMPL_WIDTH),
		22405 => to_signed(27458, LUT_AMPL_WIDTH),
		22406 => to_signed(27456, LUT_AMPL_WIDTH),
		22407 => to_signed(27454, LUT_AMPL_WIDTH),
		22408 => to_signed(27452, LUT_AMPL_WIDTH),
		22409 => to_signed(27451, LUT_AMPL_WIDTH),
		22410 => to_signed(27449, LUT_AMPL_WIDTH),
		22411 => to_signed(27447, LUT_AMPL_WIDTH),
		22412 => to_signed(27446, LUT_AMPL_WIDTH),
		22413 => to_signed(27444, LUT_AMPL_WIDTH),
		22414 => to_signed(27442, LUT_AMPL_WIDTH),
		22415 => to_signed(27440, LUT_AMPL_WIDTH),
		22416 => to_signed(27439, LUT_AMPL_WIDTH),
		22417 => to_signed(27437, LUT_AMPL_WIDTH),
		22418 => to_signed(27435, LUT_AMPL_WIDTH),
		22419 => to_signed(27434, LUT_AMPL_WIDTH),
		22420 => to_signed(27432, LUT_AMPL_WIDTH),
		22421 => to_signed(27430, LUT_AMPL_WIDTH),
		22422 => to_signed(27428, LUT_AMPL_WIDTH),
		22423 => to_signed(27427, LUT_AMPL_WIDTH),
		22424 => to_signed(27425, LUT_AMPL_WIDTH),
		22425 => to_signed(27423, LUT_AMPL_WIDTH),
		22426 => to_signed(27421, LUT_AMPL_WIDTH),
		22427 => to_signed(27420, LUT_AMPL_WIDTH),
		22428 => to_signed(27418, LUT_AMPL_WIDTH),
		22429 => to_signed(27416, LUT_AMPL_WIDTH),
		22430 => to_signed(27415, LUT_AMPL_WIDTH),
		22431 => to_signed(27413, LUT_AMPL_WIDTH),
		22432 => to_signed(27411, LUT_AMPL_WIDTH),
		22433 => to_signed(27409, LUT_AMPL_WIDTH),
		22434 => to_signed(27408, LUT_AMPL_WIDTH),
		22435 => to_signed(27406, LUT_AMPL_WIDTH),
		22436 => to_signed(27404, LUT_AMPL_WIDTH),
		22437 => to_signed(27403, LUT_AMPL_WIDTH),
		22438 => to_signed(27401, LUT_AMPL_WIDTH),
		22439 => to_signed(27399, LUT_AMPL_WIDTH),
		22440 => to_signed(27397, LUT_AMPL_WIDTH),
		22441 => to_signed(27396, LUT_AMPL_WIDTH),
		22442 => to_signed(27394, LUT_AMPL_WIDTH),
		22443 => to_signed(27392, LUT_AMPL_WIDTH),
		22444 => to_signed(27390, LUT_AMPL_WIDTH),
		22445 => to_signed(27389, LUT_AMPL_WIDTH),
		22446 => to_signed(27387, LUT_AMPL_WIDTH),
		22447 => to_signed(27385, LUT_AMPL_WIDTH),
		22448 => to_signed(27384, LUT_AMPL_WIDTH),
		22449 => to_signed(27382, LUT_AMPL_WIDTH),
		22450 => to_signed(27380, LUT_AMPL_WIDTH),
		22451 => to_signed(27378, LUT_AMPL_WIDTH),
		22452 => to_signed(27377, LUT_AMPL_WIDTH),
		22453 => to_signed(27375, LUT_AMPL_WIDTH),
		22454 => to_signed(27373, LUT_AMPL_WIDTH),
		22455 => to_signed(27372, LUT_AMPL_WIDTH),
		22456 => to_signed(27370, LUT_AMPL_WIDTH),
		22457 => to_signed(27368, LUT_AMPL_WIDTH),
		22458 => to_signed(27366, LUT_AMPL_WIDTH),
		22459 => to_signed(27365, LUT_AMPL_WIDTH),
		22460 => to_signed(27363, LUT_AMPL_WIDTH),
		22461 => to_signed(27361, LUT_AMPL_WIDTH),
		22462 => to_signed(27359, LUT_AMPL_WIDTH),
		22463 => to_signed(27358, LUT_AMPL_WIDTH),
		22464 => to_signed(27356, LUT_AMPL_WIDTH),
		22465 => to_signed(27354, LUT_AMPL_WIDTH),
		22466 => to_signed(27352, LUT_AMPL_WIDTH),
		22467 => to_signed(27351, LUT_AMPL_WIDTH),
		22468 => to_signed(27349, LUT_AMPL_WIDTH),
		22469 => to_signed(27347, LUT_AMPL_WIDTH),
		22470 => to_signed(27346, LUT_AMPL_WIDTH),
		22471 => to_signed(27344, LUT_AMPL_WIDTH),
		22472 => to_signed(27342, LUT_AMPL_WIDTH),
		22473 => to_signed(27340, LUT_AMPL_WIDTH),
		22474 => to_signed(27339, LUT_AMPL_WIDTH),
		22475 => to_signed(27337, LUT_AMPL_WIDTH),
		22476 => to_signed(27335, LUT_AMPL_WIDTH),
		22477 => to_signed(27333, LUT_AMPL_WIDTH),
		22478 => to_signed(27332, LUT_AMPL_WIDTH),
		22479 => to_signed(27330, LUT_AMPL_WIDTH),
		22480 => to_signed(27328, LUT_AMPL_WIDTH),
		22481 => to_signed(27327, LUT_AMPL_WIDTH),
		22482 => to_signed(27325, LUT_AMPL_WIDTH),
		22483 => to_signed(27323, LUT_AMPL_WIDTH),
		22484 => to_signed(27321, LUT_AMPL_WIDTH),
		22485 => to_signed(27320, LUT_AMPL_WIDTH),
		22486 => to_signed(27318, LUT_AMPL_WIDTH),
		22487 => to_signed(27316, LUT_AMPL_WIDTH),
		22488 => to_signed(27314, LUT_AMPL_WIDTH),
		22489 => to_signed(27313, LUT_AMPL_WIDTH),
		22490 => to_signed(27311, LUT_AMPL_WIDTH),
		22491 => to_signed(27309, LUT_AMPL_WIDTH),
		22492 => to_signed(27307, LUT_AMPL_WIDTH),
		22493 => to_signed(27306, LUT_AMPL_WIDTH),
		22494 => to_signed(27304, LUT_AMPL_WIDTH),
		22495 => to_signed(27302, LUT_AMPL_WIDTH),
		22496 => to_signed(27300, LUT_AMPL_WIDTH),
		22497 => to_signed(27299, LUT_AMPL_WIDTH),
		22498 => to_signed(27297, LUT_AMPL_WIDTH),
		22499 => to_signed(27295, LUT_AMPL_WIDTH),
		22500 => to_signed(27294, LUT_AMPL_WIDTH),
		22501 => to_signed(27292, LUT_AMPL_WIDTH),
		22502 => to_signed(27290, LUT_AMPL_WIDTH),
		22503 => to_signed(27288, LUT_AMPL_WIDTH),
		22504 => to_signed(27287, LUT_AMPL_WIDTH),
		22505 => to_signed(27285, LUT_AMPL_WIDTH),
		22506 => to_signed(27283, LUT_AMPL_WIDTH),
		22507 => to_signed(27281, LUT_AMPL_WIDTH),
		22508 => to_signed(27280, LUT_AMPL_WIDTH),
		22509 => to_signed(27278, LUT_AMPL_WIDTH),
		22510 => to_signed(27276, LUT_AMPL_WIDTH),
		22511 => to_signed(27274, LUT_AMPL_WIDTH),
		22512 => to_signed(27273, LUT_AMPL_WIDTH),
		22513 => to_signed(27271, LUT_AMPL_WIDTH),
		22514 => to_signed(27269, LUT_AMPL_WIDTH),
		22515 => to_signed(27267, LUT_AMPL_WIDTH),
		22516 => to_signed(27266, LUT_AMPL_WIDTH),
		22517 => to_signed(27264, LUT_AMPL_WIDTH),
		22518 => to_signed(27262, LUT_AMPL_WIDTH),
		22519 => to_signed(27260, LUT_AMPL_WIDTH),
		22520 => to_signed(27259, LUT_AMPL_WIDTH),
		22521 => to_signed(27257, LUT_AMPL_WIDTH),
		22522 => to_signed(27255, LUT_AMPL_WIDTH),
		22523 => to_signed(27253, LUT_AMPL_WIDTH),
		22524 => to_signed(27252, LUT_AMPL_WIDTH),
		22525 => to_signed(27250, LUT_AMPL_WIDTH),
		22526 => to_signed(27248, LUT_AMPL_WIDTH),
		22527 => to_signed(27247, LUT_AMPL_WIDTH),
		22528 => to_signed(27245, LUT_AMPL_WIDTH),
		22529 => to_signed(27243, LUT_AMPL_WIDTH),
		22530 => to_signed(27241, LUT_AMPL_WIDTH),
		22531 => to_signed(27240, LUT_AMPL_WIDTH),
		22532 => to_signed(27238, LUT_AMPL_WIDTH),
		22533 => to_signed(27236, LUT_AMPL_WIDTH),
		22534 => to_signed(27234, LUT_AMPL_WIDTH),
		22535 => to_signed(27233, LUT_AMPL_WIDTH),
		22536 => to_signed(27231, LUT_AMPL_WIDTH),
		22537 => to_signed(27229, LUT_AMPL_WIDTH),
		22538 => to_signed(27227, LUT_AMPL_WIDTH),
		22539 => to_signed(27226, LUT_AMPL_WIDTH),
		22540 => to_signed(27224, LUT_AMPL_WIDTH),
		22541 => to_signed(27222, LUT_AMPL_WIDTH),
		22542 => to_signed(27220, LUT_AMPL_WIDTH),
		22543 => to_signed(27219, LUT_AMPL_WIDTH),
		22544 => to_signed(27217, LUT_AMPL_WIDTH),
		22545 => to_signed(27215, LUT_AMPL_WIDTH),
		22546 => to_signed(27213, LUT_AMPL_WIDTH),
		22547 => to_signed(27212, LUT_AMPL_WIDTH),
		22548 => to_signed(27210, LUT_AMPL_WIDTH),
		22549 => to_signed(27208, LUT_AMPL_WIDTH),
		22550 => to_signed(27206, LUT_AMPL_WIDTH),
		22551 => to_signed(27205, LUT_AMPL_WIDTH),
		22552 => to_signed(27203, LUT_AMPL_WIDTH),
		22553 => to_signed(27201, LUT_AMPL_WIDTH),
		22554 => to_signed(27199, LUT_AMPL_WIDTH),
		22555 => to_signed(27198, LUT_AMPL_WIDTH),
		22556 => to_signed(27196, LUT_AMPL_WIDTH),
		22557 => to_signed(27194, LUT_AMPL_WIDTH),
		22558 => to_signed(27192, LUT_AMPL_WIDTH),
		22559 => to_signed(27191, LUT_AMPL_WIDTH),
		22560 => to_signed(27189, LUT_AMPL_WIDTH),
		22561 => to_signed(27187, LUT_AMPL_WIDTH),
		22562 => to_signed(27185, LUT_AMPL_WIDTH),
		22563 => to_signed(27184, LUT_AMPL_WIDTH),
		22564 => to_signed(27182, LUT_AMPL_WIDTH),
		22565 => to_signed(27180, LUT_AMPL_WIDTH),
		22566 => to_signed(27178, LUT_AMPL_WIDTH),
		22567 => to_signed(27177, LUT_AMPL_WIDTH),
		22568 => to_signed(27175, LUT_AMPL_WIDTH),
		22569 => to_signed(27173, LUT_AMPL_WIDTH),
		22570 => to_signed(27171, LUT_AMPL_WIDTH),
		22571 => to_signed(27169, LUT_AMPL_WIDTH),
		22572 => to_signed(27168, LUT_AMPL_WIDTH),
		22573 => to_signed(27166, LUT_AMPL_WIDTH),
		22574 => to_signed(27164, LUT_AMPL_WIDTH),
		22575 => to_signed(27162, LUT_AMPL_WIDTH),
		22576 => to_signed(27161, LUT_AMPL_WIDTH),
		22577 => to_signed(27159, LUT_AMPL_WIDTH),
		22578 => to_signed(27157, LUT_AMPL_WIDTH),
		22579 => to_signed(27155, LUT_AMPL_WIDTH),
		22580 => to_signed(27154, LUT_AMPL_WIDTH),
		22581 => to_signed(27152, LUT_AMPL_WIDTH),
		22582 => to_signed(27150, LUT_AMPL_WIDTH),
		22583 => to_signed(27148, LUT_AMPL_WIDTH),
		22584 => to_signed(27147, LUT_AMPL_WIDTH),
		22585 => to_signed(27145, LUT_AMPL_WIDTH),
		22586 => to_signed(27143, LUT_AMPL_WIDTH),
		22587 => to_signed(27141, LUT_AMPL_WIDTH),
		22588 => to_signed(27140, LUT_AMPL_WIDTH),
		22589 => to_signed(27138, LUT_AMPL_WIDTH),
		22590 => to_signed(27136, LUT_AMPL_WIDTH),
		22591 => to_signed(27134, LUT_AMPL_WIDTH),
		22592 => to_signed(27133, LUT_AMPL_WIDTH),
		22593 => to_signed(27131, LUT_AMPL_WIDTH),
		22594 => to_signed(27129, LUT_AMPL_WIDTH),
		22595 => to_signed(27127, LUT_AMPL_WIDTH),
		22596 => to_signed(27126, LUT_AMPL_WIDTH),
		22597 => to_signed(27124, LUT_AMPL_WIDTH),
		22598 => to_signed(27122, LUT_AMPL_WIDTH),
		22599 => to_signed(27120, LUT_AMPL_WIDTH),
		22600 => to_signed(27118, LUT_AMPL_WIDTH),
		22601 => to_signed(27117, LUT_AMPL_WIDTH),
		22602 => to_signed(27115, LUT_AMPL_WIDTH),
		22603 => to_signed(27113, LUT_AMPL_WIDTH),
		22604 => to_signed(27111, LUT_AMPL_WIDTH),
		22605 => to_signed(27110, LUT_AMPL_WIDTH),
		22606 => to_signed(27108, LUT_AMPL_WIDTH),
		22607 => to_signed(27106, LUT_AMPL_WIDTH),
		22608 => to_signed(27104, LUT_AMPL_WIDTH),
		22609 => to_signed(27103, LUT_AMPL_WIDTH),
		22610 => to_signed(27101, LUT_AMPL_WIDTH),
		22611 => to_signed(27099, LUT_AMPL_WIDTH),
		22612 => to_signed(27097, LUT_AMPL_WIDTH),
		22613 => to_signed(27096, LUT_AMPL_WIDTH),
		22614 => to_signed(27094, LUT_AMPL_WIDTH),
		22615 => to_signed(27092, LUT_AMPL_WIDTH),
		22616 => to_signed(27090, LUT_AMPL_WIDTH),
		22617 => to_signed(27088, LUT_AMPL_WIDTH),
		22618 => to_signed(27087, LUT_AMPL_WIDTH),
		22619 => to_signed(27085, LUT_AMPL_WIDTH),
		22620 => to_signed(27083, LUT_AMPL_WIDTH),
		22621 => to_signed(27081, LUT_AMPL_WIDTH),
		22622 => to_signed(27080, LUT_AMPL_WIDTH),
		22623 => to_signed(27078, LUT_AMPL_WIDTH),
		22624 => to_signed(27076, LUT_AMPL_WIDTH),
		22625 => to_signed(27074, LUT_AMPL_WIDTH),
		22626 => to_signed(27073, LUT_AMPL_WIDTH),
		22627 => to_signed(27071, LUT_AMPL_WIDTH),
		22628 => to_signed(27069, LUT_AMPL_WIDTH),
		22629 => to_signed(27067, LUT_AMPL_WIDTH),
		22630 => to_signed(27065, LUT_AMPL_WIDTH),
		22631 => to_signed(27064, LUT_AMPL_WIDTH),
		22632 => to_signed(27062, LUT_AMPL_WIDTH),
		22633 => to_signed(27060, LUT_AMPL_WIDTH),
		22634 => to_signed(27058, LUT_AMPL_WIDTH),
		22635 => to_signed(27057, LUT_AMPL_WIDTH),
		22636 => to_signed(27055, LUT_AMPL_WIDTH),
		22637 => to_signed(27053, LUT_AMPL_WIDTH),
		22638 => to_signed(27051, LUT_AMPL_WIDTH),
		22639 => to_signed(27049, LUT_AMPL_WIDTH),
		22640 => to_signed(27048, LUT_AMPL_WIDTH),
		22641 => to_signed(27046, LUT_AMPL_WIDTH),
		22642 => to_signed(27044, LUT_AMPL_WIDTH),
		22643 => to_signed(27042, LUT_AMPL_WIDTH),
		22644 => to_signed(27041, LUT_AMPL_WIDTH),
		22645 => to_signed(27039, LUT_AMPL_WIDTH),
		22646 => to_signed(27037, LUT_AMPL_WIDTH),
		22647 => to_signed(27035, LUT_AMPL_WIDTH),
		22648 => to_signed(27034, LUT_AMPL_WIDTH),
		22649 => to_signed(27032, LUT_AMPL_WIDTH),
		22650 => to_signed(27030, LUT_AMPL_WIDTH),
		22651 => to_signed(27028, LUT_AMPL_WIDTH),
		22652 => to_signed(27026, LUT_AMPL_WIDTH),
		22653 => to_signed(27025, LUT_AMPL_WIDTH),
		22654 => to_signed(27023, LUT_AMPL_WIDTH),
		22655 => to_signed(27021, LUT_AMPL_WIDTH),
		22656 => to_signed(27019, LUT_AMPL_WIDTH),
		22657 => to_signed(27018, LUT_AMPL_WIDTH),
		22658 => to_signed(27016, LUT_AMPL_WIDTH),
		22659 => to_signed(27014, LUT_AMPL_WIDTH),
		22660 => to_signed(27012, LUT_AMPL_WIDTH),
		22661 => to_signed(27010, LUT_AMPL_WIDTH),
		22662 => to_signed(27009, LUT_AMPL_WIDTH),
		22663 => to_signed(27007, LUT_AMPL_WIDTH),
		22664 => to_signed(27005, LUT_AMPL_WIDTH),
		22665 => to_signed(27003, LUT_AMPL_WIDTH),
		22666 => to_signed(27002, LUT_AMPL_WIDTH),
		22667 => to_signed(27000, LUT_AMPL_WIDTH),
		22668 => to_signed(26998, LUT_AMPL_WIDTH),
		22669 => to_signed(26996, LUT_AMPL_WIDTH),
		22670 => to_signed(26994, LUT_AMPL_WIDTH),
		22671 => to_signed(26993, LUT_AMPL_WIDTH),
		22672 => to_signed(26991, LUT_AMPL_WIDTH),
		22673 => to_signed(26989, LUT_AMPL_WIDTH),
		22674 => to_signed(26987, LUT_AMPL_WIDTH),
		22675 => to_signed(26986, LUT_AMPL_WIDTH),
		22676 => to_signed(26984, LUT_AMPL_WIDTH),
		22677 => to_signed(26982, LUT_AMPL_WIDTH),
		22678 => to_signed(26980, LUT_AMPL_WIDTH),
		22679 => to_signed(26978, LUT_AMPL_WIDTH),
		22680 => to_signed(26977, LUT_AMPL_WIDTH),
		22681 => to_signed(26975, LUT_AMPL_WIDTH),
		22682 => to_signed(26973, LUT_AMPL_WIDTH),
		22683 => to_signed(26971, LUT_AMPL_WIDTH),
		22684 => to_signed(26969, LUT_AMPL_WIDTH),
		22685 => to_signed(26968, LUT_AMPL_WIDTH),
		22686 => to_signed(26966, LUT_AMPL_WIDTH),
		22687 => to_signed(26964, LUT_AMPL_WIDTH),
		22688 => to_signed(26962, LUT_AMPL_WIDTH),
		22689 => to_signed(26961, LUT_AMPL_WIDTH),
		22690 => to_signed(26959, LUT_AMPL_WIDTH),
		22691 => to_signed(26957, LUT_AMPL_WIDTH),
		22692 => to_signed(26955, LUT_AMPL_WIDTH),
		22693 => to_signed(26953, LUT_AMPL_WIDTH),
		22694 => to_signed(26952, LUT_AMPL_WIDTH),
		22695 => to_signed(26950, LUT_AMPL_WIDTH),
		22696 => to_signed(26948, LUT_AMPL_WIDTH),
		22697 => to_signed(26946, LUT_AMPL_WIDTH),
		22698 => to_signed(26944, LUT_AMPL_WIDTH),
		22699 => to_signed(26943, LUT_AMPL_WIDTH),
		22700 => to_signed(26941, LUT_AMPL_WIDTH),
		22701 => to_signed(26939, LUT_AMPL_WIDTH),
		22702 => to_signed(26937, LUT_AMPL_WIDTH),
		22703 => to_signed(26936, LUT_AMPL_WIDTH),
		22704 => to_signed(26934, LUT_AMPL_WIDTH),
		22705 => to_signed(26932, LUT_AMPL_WIDTH),
		22706 => to_signed(26930, LUT_AMPL_WIDTH),
		22707 => to_signed(26928, LUT_AMPL_WIDTH),
		22708 => to_signed(26927, LUT_AMPL_WIDTH),
		22709 => to_signed(26925, LUT_AMPL_WIDTH),
		22710 => to_signed(26923, LUT_AMPL_WIDTH),
		22711 => to_signed(26921, LUT_AMPL_WIDTH),
		22712 => to_signed(26919, LUT_AMPL_WIDTH),
		22713 => to_signed(26918, LUT_AMPL_WIDTH),
		22714 => to_signed(26916, LUT_AMPL_WIDTH),
		22715 => to_signed(26914, LUT_AMPL_WIDTH),
		22716 => to_signed(26912, LUT_AMPL_WIDTH),
		22717 => to_signed(26910, LUT_AMPL_WIDTH),
		22718 => to_signed(26909, LUT_AMPL_WIDTH),
		22719 => to_signed(26907, LUT_AMPL_WIDTH),
		22720 => to_signed(26905, LUT_AMPL_WIDTH),
		22721 => to_signed(26903, LUT_AMPL_WIDTH),
		22722 => to_signed(26901, LUT_AMPL_WIDTH),
		22723 => to_signed(26900, LUT_AMPL_WIDTH),
		22724 => to_signed(26898, LUT_AMPL_WIDTH),
		22725 => to_signed(26896, LUT_AMPL_WIDTH),
		22726 => to_signed(26894, LUT_AMPL_WIDTH),
		22727 => to_signed(26893, LUT_AMPL_WIDTH),
		22728 => to_signed(26891, LUT_AMPL_WIDTH),
		22729 => to_signed(26889, LUT_AMPL_WIDTH),
		22730 => to_signed(26887, LUT_AMPL_WIDTH),
		22731 => to_signed(26885, LUT_AMPL_WIDTH),
		22732 => to_signed(26884, LUT_AMPL_WIDTH),
		22733 => to_signed(26882, LUT_AMPL_WIDTH),
		22734 => to_signed(26880, LUT_AMPL_WIDTH),
		22735 => to_signed(26878, LUT_AMPL_WIDTH),
		22736 => to_signed(26876, LUT_AMPL_WIDTH),
		22737 => to_signed(26875, LUT_AMPL_WIDTH),
		22738 => to_signed(26873, LUT_AMPL_WIDTH),
		22739 => to_signed(26871, LUT_AMPL_WIDTH),
		22740 => to_signed(26869, LUT_AMPL_WIDTH),
		22741 => to_signed(26867, LUT_AMPL_WIDTH),
		22742 => to_signed(26866, LUT_AMPL_WIDTH),
		22743 => to_signed(26864, LUT_AMPL_WIDTH),
		22744 => to_signed(26862, LUT_AMPL_WIDTH),
		22745 => to_signed(26860, LUT_AMPL_WIDTH),
		22746 => to_signed(26858, LUT_AMPL_WIDTH),
		22747 => to_signed(26857, LUT_AMPL_WIDTH),
		22748 => to_signed(26855, LUT_AMPL_WIDTH),
		22749 => to_signed(26853, LUT_AMPL_WIDTH),
		22750 => to_signed(26851, LUT_AMPL_WIDTH),
		22751 => to_signed(26849, LUT_AMPL_WIDTH),
		22752 => to_signed(26848, LUT_AMPL_WIDTH),
		22753 => to_signed(26846, LUT_AMPL_WIDTH),
		22754 => to_signed(26844, LUT_AMPL_WIDTH),
		22755 => to_signed(26842, LUT_AMPL_WIDTH),
		22756 => to_signed(26840, LUT_AMPL_WIDTH),
		22757 => to_signed(26839, LUT_AMPL_WIDTH),
		22758 => to_signed(26837, LUT_AMPL_WIDTH),
		22759 => to_signed(26835, LUT_AMPL_WIDTH),
		22760 => to_signed(26833, LUT_AMPL_WIDTH),
		22761 => to_signed(26831, LUT_AMPL_WIDTH),
		22762 => to_signed(26830, LUT_AMPL_WIDTH),
		22763 => to_signed(26828, LUT_AMPL_WIDTH),
		22764 => to_signed(26826, LUT_AMPL_WIDTH),
		22765 => to_signed(26824, LUT_AMPL_WIDTH),
		22766 => to_signed(26822, LUT_AMPL_WIDTH),
		22767 => to_signed(26821, LUT_AMPL_WIDTH),
		22768 => to_signed(26819, LUT_AMPL_WIDTH),
		22769 => to_signed(26817, LUT_AMPL_WIDTH),
		22770 => to_signed(26815, LUT_AMPL_WIDTH),
		22771 => to_signed(26813, LUT_AMPL_WIDTH),
		22772 => to_signed(26811, LUT_AMPL_WIDTH),
		22773 => to_signed(26810, LUT_AMPL_WIDTH),
		22774 => to_signed(26808, LUT_AMPL_WIDTH),
		22775 => to_signed(26806, LUT_AMPL_WIDTH),
		22776 => to_signed(26804, LUT_AMPL_WIDTH),
		22777 => to_signed(26802, LUT_AMPL_WIDTH),
		22778 => to_signed(26801, LUT_AMPL_WIDTH),
		22779 => to_signed(26799, LUT_AMPL_WIDTH),
		22780 => to_signed(26797, LUT_AMPL_WIDTH),
		22781 => to_signed(26795, LUT_AMPL_WIDTH),
		22782 => to_signed(26793, LUT_AMPL_WIDTH),
		22783 => to_signed(26792, LUT_AMPL_WIDTH),
		22784 => to_signed(26790, LUT_AMPL_WIDTH),
		22785 => to_signed(26788, LUT_AMPL_WIDTH),
		22786 => to_signed(26786, LUT_AMPL_WIDTH),
		22787 => to_signed(26784, LUT_AMPL_WIDTH),
		22788 => to_signed(26783, LUT_AMPL_WIDTH),
		22789 => to_signed(26781, LUT_AMPL_WIDTH),
		22790 => to_signed(26779, LUT_AMPL_WIDTH),
		22791 => to_signed(26777, LUT_AMPL_WIDTH),
		22792 => to_signed(26775, LUT_AMPL_WIDTH),
		22793 => to_signed(26774, LUT_AMPL_WIDTH),
		22794 => to_signed(26772, LUT_AMPL_WIDTH),
		22795 => to_signed(26770, LUT_AMPL_WIDTH),
		22796 => to_signed(26768, LUT_AMPL_WIDTH),
		22797 => to_signed(26766, LUT_AMPL_WIDTH),
		22798 => to_signed(26764, LUT_AMPL_WIDTH),
		22799 => to_signed(26763, LUT_AMPL_WIDTH),
		22800 => to_signed(26761, LUT_AMPL_WIDTH),
		22801 => to_signed(26759, LUT_AMPL_WIDTH),
		22802 => to_signed(26757, LUT_AMPL_WIDTH),
		22803 => to_signed(26755, LUT_AMPL_WIDTH),
		22804 => to_signed(26754, LUT_AMPL_WIDTH),
		22805 => to_signed(26752, LUT_AMPL_WIDTH),
		22806 => to_signed(26750, LUT_AMPL_WIDTH),
		22807 => to_signed(26748, LUT_AMPL_WIDTH),
		22808 => to_signed(26746, LUT_AMPL_WIDTH),
		22809 => to_signed(26745, LUT_AMPL_WIDTH),
		22810 => to_signed(26743, LUT_AMPL_WIDTH),
		22811 => to_signed(26741, LUT_AMPL_WIDTH),
		22812 => to_signed(26739, LUT_AMPL_WIDTH),
		22813 => to_signed(26737, LUT_AMPL_WIDTH),
		22814 => to_signed(26735, LUT_AMPL_WIDTH),
		22815 => to_signed(26734, LUT_AMPL_WIDTH),
		22816 => to_signed(26732, LUT_AMPL_WIDTH),
		22817 => to_signed(26730, LUT_AMPL_WIDTH),
		22818 => to_signed(26728, LUT_AMPL_WIDTH),
		22819 => to_signed(26726, LUT_AMPL_WIDTH),
		22820 => to_signed(26725, LUT_AMPL_WIDTH),
		22821 => to_signed(26723, LUT_AMPL_WIDTH),
		22822 => to_signed(26721, LUT_AMPL_WIDTH),
		22823 => to_signed(26719, LUT_AMPL_WIDTH),
		22824 => to_signed(26717, LUT_AMPL_WIDTH),
		22825 => to_signed(26715, LUT_AMPL_WIDTH),
		22826 => to_signed(26714, LUT_AMPL_WIDTH),
		22827 => to_signed(26712, LUT_AMPL_WIDTH),
		22828 => to_signed(26710, LUT_AMPL_WIDTH),
		22829 => to_signed(26708, LUT_AMPL_WIDTH),
		22830 => to_signed(26706, LUT_AMPL_WIDTH),
		22831 => to_signed(26705, LUT_AMPL_WIDTH),
		22832 => to_signed(26703, LUT_AMPL_WIDTH),
		22833 => to_signed(26701, LUT_AMPL_WIDTH),
		22834 => to_signed(26699, LUT_AMPL_WIDTH),
		22835 => to_signed(26697, LUT_AMPL_WIDTH),
		22836 => to_signed(26695, LUT_AMPL_WIDTH),
		22837 => to_signed(26694, LUT_AMPL_WIDTH),
		22838 => to_signed(26692, LUT_AMPL_WIDTH),
		22839 => to_signed(26690, LUT_AMPL_WIDTH),
		22840 => to_signed(26688, LUT_AMPL_WIDTH),
		22841 => to_signed(26686, LUT_AMPL_WIDTH),
		22842 => to_signed(26684, LUT_AMPL_WIDTH),
		22843 => to_signed(26683, LUT_AMPL_WIDTH),
		22844 => to_signed(26681, LUT_AMPL_WIDTH),
		22845 => to_signed(26679, LUT_AMPL_WIDTH),
		22846 => to_signed(26677, LUT_AMPL_WIDTH),
		22847 => to_signed(26675, LUT_AMPL_WIDTH),
		22848 => to_signed(26674, LUT_AMPL_WIDTH),
		22849 => to_signed(26672, LUT_AMPL_WIDTH),
		22850 => to_signed(26670, LUT_AMPL_WIDTH),
		22851 => to_signed(26668, LUT_AMPL_WIDTH),
		22852 => to_signed(26666, LUT_AMPL_WIDTH),
		22853 => to_signed(26664, LUT_AMPL_WIDTH),
		22854 => to_signed(26663, LUT_AMPL_WIDTH),
		22855 => to_signed(26661, LUT_AMPL_WIDTH),
		22856 => to_signed(26659, LUT_AMPL_WIDTH),
		22857 => to_signed(26657, LUT_AMPL_WIDTH),
		22858 => to_signed(26655, LUT_AMPL_WIDTH),
		22859 => to_signed(26653, LUT_AMPL_WIDTH),
		22860 => to_signed(26652, LUT_AMPL_WIDTH),
		22861 => to_signed(26650, LUT_AMPL_WIDTH),
		22862 => to_signed(26648, LUT_AMPL_WIDTH),
		22863 => to_signed(26646, LUT_AMPL_WIDTH),
		22864 => to_signed(26644, LUT_AMPL_WIDTH),
		22865 => to_signed(26642, LUT_AMPL_WIDTH),
		22866 => to_signed(26641, LUT_AMPL_WIDTH),
		22867 => to_signed(26639, LUT_AMPL_WIDTH),
		22868 => to_signed(26637, LUT_AMPL_WIDTH),
		22869 => to_signed(26635, LUT_AMPL_WIDTH),
		22870 => to_signed(26633, LUT_AMPL_WIDTH),
		22871 => to_signed(26631, LUT_AMPL_WIDTH),
		22872 => to_signed(26630, LUT_AMPL_WIDTH),
		22873 => to_signed(26628, LUT_AMPL_WIDTH),
		22874 => to_signed(26626, LUT_AMPL_WIDTH),
		22875 => to_signed(26624, LUT_AMPL_WIDTH),
		22876 => to_signed(26622, LUT_AMPL_WIDTH),
		22877 => to_signed(26621, LUT_AMPL_WIDTH),
		22878 => to_signed(26619, LUT_AMPL_WIDTH),
		22879 => to_signed(26617, LUT_AMPL_WIDTH),
		22880 => to_signed(26615, LUT_AMPL_WIDTH),
		22881 => to_signed(26613, LUT_AMPL_WIDTH),
		22882 => to_signed(26611, LUT_AMPL_WIDTH),
		22883 => to_signed(26610, LUT_AMPL_WIDTH),
		22884 => to_signed(26608, LUT_AMPL_WIDTH),
		22885 => to_signed(26606, LUT_AMPL_WIDTH),
		22886 => to_signed(26604, LUT_AMPL_WIDTH),
		22887 => to_signed(26602, LUT_AMPL_WIDTH),
		22888 => to_signed(26600, LUT_AMPL_WIDTH),
		22889 => to_signed(26599, LUT_AMPL_WIDTH),
		22890 => to_signed(26597, LUT_AMPL_WIDTH),
		22891 => to_signed(26595, LUT_AMPL_WIDTH),
		22892 => to_signed(26593, LUT_AMPL_WIDTH),
		22893 => to_signed(26591, LUT_AMPL_WIDTH),
		22894 => to_signed(26589, LUT_AMPL_WIDTH),
		22895 => to_signed(26588, LUT_AMPL_WIDTH),
		22896 => to_signed(26586, LUT_AMPL_WIDTH),
		22897 => to_signed(26584, LUT_AMPL_WIDTH),
		22898 => to_signed(26582, LUT_AMPL_WIDTH),
		22899 => to_signed(26580, LUT_AMPL_WIDTH),
		22900 => to_signed(26578, LUT_AMPL_WIDTH),
		22901 => to_signed(26576, LUT_AMPL_WIDTH),
		22902 => to_signed(26575, LUT_AMPL_WIDTH),
		22903 => to_signed(26573, LUT_AMPL_WIDTH),
		22904 => to_signed(26571, LUT_AMPL_WIDTH),
		22905 => to_signed(26569, LUT_AMPL_WIDTH),
		22906 => to_signed(26567, LUT_AMPL_WIDTH),
		22907 => to_signed(26565, LUT_AMPL_WIDTH),
		22908 => to_signed(26564, LUT_AMPL_WIDTH),
		22909 => to_signed(26562, LUT_AMPL_WIDTH),
		22910 => to_signed(26560, LUT_AMPL_WIDTH),
		22911 => to_signed(26558, LUT_AMPL_WIDTH),
		22912 => to_signed(26556, LUT_AMPL_WIDTH),
		22913 => to_signed(26554, LUT_AMPL_WIDTH),
		22914 => to_signed(26553, LUT_AMPL_WIDTH),
		22915 => to_signed(26551, LUT_AMPL_WIDTH),
		22916 => to_signed(26549, LUT_AMPL_WIDTH),
		22917 => to_signed(26547, LUT_AMPL_WIDTH),
		22918 => to_signed(26545, LUT_AMPL_WIDTH),
		22919 => to_signed(26543, LUT_AMPL_WIDTH),
		22920 => to_signed(26542, LUT_AMPL_WIDTH),
		22921 => to_signed(26540, LUT_AMPL_WIDTH),
		22922 => to_signed(26538, LUT_AMPL_WIDTH),
		22923 => to_signed(26536, LUT_AMPL_WIDTH),
		22924 => to_signed(26534, LUT_AMPL_WIDTH),
		22925 => to_signed(26532, LUT_AMPL_WIDTH),
		22926 => to_signed(26530, LUT_AMPL_WIDTH),
		22927 => to_signed(26529, LUT_AMPL_WIDTH),
		22928 => to_signed(26527, LUT_AMPL_WIDTH),
		22929 => to_signed(26525, LUT_AMPL_WIDTH),
		22930 => to_signed(26523, LUT_AMPL_WIDTH),
		22931 => to_signed(26521, LUT_AMPL_WIDTH),
		22932 => to_signed(26519, LUT_AMPL_WIDTH),
		22933 => to_signed(26518, LUT_AMPL_WIDTH),
		22934 => to_signed(26516, LUT_AMPL_WIDTH),
		22935 => to_signed(26514, LUT_AMPL_WIDTH),
		22936 => to_signed(26512, LUT_AMPL_WIDTH),
		22937 => to_signed(26510, LUT_AMPL_WIDTH),
		22938 => to_signed(26508, LUT_AMPL_WIDTH),
		22939 => to_signed(26506, LUT_AMPL_WIDTH),
		22940 => to_signed(26505, LUT_AMPL_WIDTH),
		22941 => to_signed(26503, LUT_AMPL_WIDTH),
		22942 => to_signed(26501, LUT_AMPL_WIDTH),
		22943 => to_signed(26499, LUT_AMPL_WIDTH),
		22944 => to_signed(26497, LUT_AMPL_WIDTH),
		22945 => to_signed(26495, LUT_AMPL_WIDTH),
		22946 => to_signed(26494, LUT_AMPL_WIDTH),
		22947 => to_signed(26492, LUT_AMPL_WIDTH),
		22948 => to_signed(26490, LUT_AMPL_WIDTH),
		22949 => to_signed(26488, LUT_AMPL_WIDTH),
		22950 => to_signed(26486, LUT_AMPL_WIDTH),
		22951 => to_signed(26484, LUT_AMPL_WIDTH),
		22952 => to_signed(26482, LUT_AMPL_WIDTH),
		22953 => to_signed(26481, LUT_AMPL_WIDTH),
		22954 => to_signed(26479, LUT_AMPL_WIDTH),
		22955 => to_signed(26477, LUT_AMPL_WIDTH),
		22956 => to_signed(26475, LUT_AMPL_WIDTH),
		22957 => to_signed(26473, LUT_AMPL_WIDTH),
		22958 => to_signed(26471, LUT_AMPL_WIDTH),
		22959 => to_signed(26469, LUT_AMPL_WIDTH),
		22960 => to_signed(26468, LUT_AMPL_WIDTH),
		22961 => to_signed(26466, LUT_AMPL_WIDTH),
		22962 => to_signed(26464, LUT_AMPL_WIDTH),
		22963 => to_signed(26462, LUT_AMPL_WIDTH),
		22964 => to_signed(26460, LUT_AMPL_WIDTH),
		22965 => to_signed(26458, LUT_AMPL_WIDTH),
		22966 => to_signed(26457, LUT_AMPL_WIDTH),
		22967 => to_signed(26455, LUT_AMPL_WIDTH),
		22968 => to_signed(26453, LUT_AMPL_WIDTH),
		22969 => to_signed(26451, LUT_AMPL_WIDTH),
		22970 => to_signed(26449, LUT_AMPL_WIDTH),
		22971 => to_signed(26447, LUT_AMPL_WIDTH),
		22972 => to_signed(26445, LUT_AMPL_WIDTH),
		22973 => to_signed(26444, LUT_AMPL_WIDTH),
		22974 => to_signed(26442, LUT_AMPL_WIDTH),
		22975 => to_signed(26440, LUT_AMPL_WIDTH),
		22976 => to_signed(26438, LUT_AMPL_WIDTH),
		22977 => to_signed(26436, LUT_AMPL_WIDTH),
		22978 => to_signed(26434, LUT_AMPL_WIDTH),
		22979 => to_signed(26432, LUT_AMPL_WIDTH),
		22980 => to_signed(26431, LUT_AMPL_WIDTH),
		22981 => to_signed(26429, LUT_AMPL_WIDTH),
		22982 => to_signed(26427, LUT_AMPL_WIDTH),
		22983 => to_signed(26425, LUT_AMPL_WIDTH),
		22984 => to_signed(26423, LUT_AMPL_WIDTH),
		22985 => to_signed(26421, LUT_AMPL_WIDTH),
		22986 => to_signed(26419, LUT_AMPL_WIDTH),
		22987 => to_signed(26418, LUT_AMPL_WIDTH),
		22988 => to_signed(26416, LUT_AMPL_WIDTH),
		22989 => to_signed(26414, LUT_AMPL_WIDTH),
		22990 => to_signed(26412, LUT_AMPL_WIDTH),
		22991 => to_signed(26410, LUT_AMPL_WIDTH),
		22992 => to_signed(26408, LUT_AMPL_WIDTH),
		22993 => to_signed(26406, LUT_AMPL_WIDTH),
		22994 => to_signed(26405, LUT_AMPL_WIDTH),
		22995 => to_signed(26403, LUT_AMPL_WIDTH),
		22996 => to_signed(26401, LUT_AMPL_WIDTH),
		22997 => to_signed(26399, LUT_AMPL_WIDTH),
		22998 => to_signed(26397, LUT_AMPL_WIDTH),
		22999 => to_signed(26395, LUT_AMPL_WIDTH),
		23000 => to_signed(26393, LUT_AMPL_WIDTH),
		23001 => to_signed(26392, LUT_AMPL_WIDTH),
		23002 => to_signed(26390, LUT_AMPL_WIDTH),
		23003 => to_signed(26388, LUT_AMPL_WIDTH),
		23004 => to_signed(26386, LUT_AMPL_WIDTH),
		23005 => to_signed(26384, LUT_AMPL_WIDTH),
		23006 => to_signed(26382, LUT_AMPL_WIDTH),
		23007 => to_signed(26380, LUT_AMPL_WIDTH),
		23008 => to_signed(26378, LUT_AMPL_WIDTH),
		23009 => to_signed(26377, LUT_AMPL_WIDTH),
		23010 => to_signed(26375, LUT_AMPL_WIDTH),
		23011 => to_signed(26373, LUT_AMPL_WIDTH),
		23012 => to_signed(26371, LUT_AMPL_WIDTH),
		23013 => to_signed(26369, LUT_AMPL_WIDTH),
		23014 => to_signed(26367, LUT_AMPL_WIDTH),
		23015 => to_signed(26365, LUT_AMPL_WIDTH),
		23016 => to_signed(26364, LUT_AMPL_WIDTH),
		23017 => to_signed(26362, LUT_AMPL_WIDTH),
		23018 => to_signed(26360, LUT_AMPL_WIDTH),
		23019 => to_signed(26358, LUT_AMPL_WIDTH),
		23020 => to_signed(26356, LUT_AMPL_WIDTH),
		23021 => to_signed(26354, LUT_AMPL_WIDTH),
		23022 => to_signed(26352, LUT_AMPL_WIDTH),
		23023 => to_signed(26350, LUT_AMPL_WIDTH),
		23024 => to_signed(26349, LUT_AMPL_WIDTH),
		23025 => to_signed(26347, LUT_AMPL_WIDTH),
		23026 => to_signed(26345, LUT_AMPL_WIDTH),
		23027 => to_signed(26343, LUT_AMPL_WIDTH),
		23028 => to_signed(26341, LUT_AMPL_WIDTH),
		23029 => to_signed(26339, LUT_AMPL_WIDTH),
		23030 => to_signed(26337, LUT_AMPL_WIDTH),
		23031 => to_signed(26336, LUT_AMPL_WIDTH),
		23032 => to_signed(26334, LUT_AMPL_WIDTH),
		23033 => to_signed(26332, LUT_AMPL_WIDTH),
		23034 => to_signed(26330, LUT_AMPL_WIDTH),
		23035 => to_signed(26328, LUT_AMPL_WIDTH),
		23036 => to_signed(26326, LUT_AMPL_WIDTH),
		23037 => to_signed(26324, LUT_AMPL_WIDTH),
		23038 => to_signed(26322, LUT_AMPL_WIDTH),
		23039 => to_signed(26321, LUT_AMPL_WIDTH),
		23040 => to_signed(26319, LUT_AMPL_WIDTH),
		23041 => to_signed(26317, LUT_AMPL_WIDTH),
		23042 => to_signed(26315, LUT_AMPL_WIDTH),
		23043 => to_signed(26313, LUT_AMPL_WIDTH),
		23044 => to_signed(26311, LUT_AMPL_WIDTH),
		23045 => to_signed(26309, LUT_AMPL_WIDTH),
		23046 => to_signed(26307, LUT_AMPL_WIDTH),
		23047 => to_signed(26306, LUT_AMPL_WIDTH),
		23048 => to_signed(26304, LUT_AMPL_WIDTH),
		23049 => to_signed(26302, LUT_AMPL_WIDTH),
		23050 => to_signed(26300, LUT_AMPL_WIDTH),
		23051 => to_signed(26298, LUT_AMPL_WIDTH),
		23052 => to_signed(26296, LUT_AMPL_WIDTH),
		23053 => to_signed(26294, LUT_AMPL_WIDTH),
		23054 => to_signed(26292, LUT_AMPL_WIDTH),
		23055 => to_signed(26291, LUT_AMPL_WIDTH),
		23056 => to_signed(26289, LUT_AMPL_WIDTH),
		23057 => to_signed(26287, LUT_AMPL_WIDTH),
		23058 => to_signed(26285, LUT_AMPL_WIDTH),
		23059 => to_signed(26283, LUT_AMPL_WIDTH),
		23060 => to_signed(26281, LUT_AMPL_WIDTH),
		23061 => to_signed(26279, LUT_AMPL_WIDTH),
		23062 => to_signed(26277, LUT_AMPL_WIDTH),
		23063 => to_signed(26276, LUT_AMPL_WIDTH),
		23064 => to_signed(26274, LUT_AMPL_WIDTH),
		23065 => to_signed(26272, LUT_AMPL_WIDTH),
		23066 => to_signed(26270, LUT_AMPL_WIDTH),
		23067 => to_signed(26268, LUT_AMPL_WIDTH),
		23068 => to_signed(26266, LUT_AMPL_WIDTH),
		23069 => to_signed(26264, LUT_AMPL_WIDTH),
		23070 => to_signed(26262, LUT_AMPL_WIDTH),
		23071 => to_signed(26261, LUT_AMPL_WIDTH),
		23072 => to_signed(26259, LUT_AMPL_WIDTH),
		23073 => to_signed(26257, LUT_AMPL_WIDTH),
		23074 => to_signed(26255, LUT_AMPL_WIDTH),
		23075 => to_signed(26253, LUT_AMPL_WIDTH),
		23076 => to_signed(26251, LUT_AMPL_WIDTH),
		23077 => to_signed(26249, LUT_AMPL_WIDTH),
		23078 => to_signed(26247, LUT_AMPL_WIDTH),
		23079 => to_signed(26246, LUT_AMPL_WIDTH),
		23080 => to_signed(26244, LUT_AMPL_WIDTH),
		23081 => to_signed(26242, LUT_AMPL_WIDTH),
		23082 => to_signed(26240, LUT_AMPL_WIDTH),
		23083 => to_signed(26238, LUT_AMPL_WIDTH),
		23084 => to_signed(26236, LUT_AMPL_WIDTH),
		23085 => to_signed(26234, LUT_AMPL_WIDTH),
		23086 => to_signed(26232, LUT_AMPL_WIDTH),
		23087 => to_signed(26230, LUT_AMPL_WIDTH),
		23088 => to_signed(26229, LUT_AMPL_WIDTH),
		23089 => to_signed(26227, LUT_AMPL_WIDTH),
		23090 => to_signed(26225, LUT_AMPL_WIDTH),
		23091 => to_signed(26223, LUT_AMPL_WIDTH),
		23092 => to_signed(26221, LUT_AMPL_WIDTH),
		23093 => to_signed(26219, LUT_AMPL_WIDTH),
		23094 => to_signed(26217, LUT_AMPL_WIDTH),
		23095 => to_signed(26215, LUT_AMPL_WIDTH),
		23096 => to_signed(26214, LUT_AMPL_WIDTH),
		23097 => to_signed(26212, LUT_AMPL_WIDTH),
		23098 => to_signed(26210, LUT_AMPL_WIDTH),
		23099 => to_signed(26208, LUT_AMPL_WIDTH),
		23100 => to_signed(26206, LUT_AMPL_WIDTH),
		23101 => to_signed(26204, LUT_AMPL_WIDTH),
		23102 => to_signed(26202, LUT_AMPL_WIDTH),
		23103 => to_signed(26200, LUT_AMPL_WIDTH),
		23104 => to_signed(26198, LUT_AMPL_WIDTH),
		23105 => to_signed(26197, LUT_AMPL_WIDTH),
		23106 => to_signed(26195, LUT_AMPL_WIDTH),
		23107 => to_signed(26193, LUT_AMPL_WIDTH),
		23108 => to_signed(26191, LUT_AMPL_WIDTH),
		23109 => to_signed(26189, LUT_AMPL_WIDTH),
		23110 => to_signed(26187, LUT_AMPL_WIDTH),
		23111 => to_signed(26185, LUT_AMPL_WIDTH),
		23112 => to_signed(26183, LUT_AMPL_WIDTH),
		23113 => to_signed(26181, LUT_AMPL_WIDTH),
		23114 => to_signed(26180, LUT_AMPL_WIDTH),
		23115 => to_signed(26178, LUT_AMPL_WIDTH),
		23116 => to_signed(26176, LUT_AMPL_WIDTH),
		23117 => to_signed(26174, LUT_AMPL_WIDTH),
		23118 => to_signed(26172, LUT_AMPL_WIDTH),
		23119 => to_signed(26170, LUT_AMPL_WIDTH),
		23120 => to_signed(26168, LUT_AMPL_WIDTH),
		23121 => to_signed(26166, LUT_AMPL_WIDTH),
		23122 => to_signed(26164, LUT_AMPL_WIDTH),
		23123 => to_signed(26163, LUT_AMPL_WIDTH),
		23124 => to_signed(26161, LUT_AMPL_WIDTH),
		23125 => to_signed(26159, LUT_AMPL_WIDTH),
		23126 => to_signed(26157, LUT_AMPL_WIDTH),
		23127 => to_signed(26155, LUT_AMPL_WIDTH),
		23128 => to_signed(26153, LUT_AMPL_WIDTH),
		23129 => to_signed(26151, LUT_AMPL_WIDTH),
		23130 => to_signed(26149, LUT_AMPL_WIDTH),
		23131 => to_signed(26147, LUT_AMPL_WIDTH),
		23132 => to_signed(26146, LUT_AMPL_WIDTH),
		23133 => to_signed(26144, LUT_AMPL_WIDTH),
		23134 => to_signed(26142, LUT_AMPL_WIDTH),
		23135 => to_signed(26140, LUT_AMPL_WIDTH),
		23136 => to_signed(26138, LUT_AMPL_WIDTH),
		23137 => to_signed(26136, LUT_AMPL_WIDTH),
		23138 => to_signed(26134, LUT_AMPL_WIDTH),
		23139 => to_signed(26132, LUT_AMPL_WIDTH),
		23140 => to_signed(26130, LUT_AMPL_WIDTH),
		23141 => to_signed(26128, LUT_AMPL_WIDTH),
		23142 => to_signed(26127, LUT_AMPL_WIDTH),
		23143 => to_signed(26125, LUT_AMPL_WIDTH),
		23144 => to_signed(26123, LUT_AMPL_WIDTH),
		23145 => to_signed(26121, LUT_AMPL_WIDTH),
		23146 => to_signed(26119, LUT_AMPL_WIDTH),
		23147 => to_signed(26117, LUT_AMPL_WIDTH),
		23148 => to_signed(26115, LUT_AMPL_WIDTH),
		23149 => to_signed(26113, LUT_AMPL_WIDTH),
		23150 => to_signed(26111, LUT_AMPL_WIDTH),
		23151 => to_signed(26109, LUT_AMPL_WIDTH),
		23152 => to_signed(26108, LUT_AMPL_WIDTH),
		23153 => to_signed(26106, LUT_AMPL_WIDTH),
		23154 => to_signed(26104, LUT_AMPL_WIDTH),
		23155 => to_signed(26102, LUT_AMPL_WIDTH),
		23156 => to_signed(26100, LUT_AMPL_WIDTH),
		23157 => to_signed(26098, LUT_AMPL_WIDTH),
		23158 => to_signed(26096, LUT_AMPL_WIDTH),
		23159 => to_signed(26094, LUT_AMPL_WIDTH),
		23160 => to_signed(26092, LUT_AMPL_WIDTH),
		23161 => to_signed(26090, LUT_AMPL_WIDTH),
		23162 => to_signed(26089, LUT_AMPL_WIDTH),
		23163 => to_signed(26087, LUT_AMPL_WIDTH),
		23164 => to_signed(26085, LUT_AMPL_WIDTH),
		23165 => to_signed(26083, LUT_AMPL_WIDTH),
		23166 => to_signed(26081, LUT_AMPL_WIDTH),
		23167 => to_signed(26079, LUT_AMPL_WIDTH),
		23168 => to_signed(26077, LUT_AMPL_WIDTH),
		23169 => to_signed(26075, LUT_AMPL_WIDTH),
		23170 => to_signed(26073, LUT_AMPL_WIDTH),
		23171 => to_signed(26071, LUT_AMPL_WIDTH),
		23172 => to_signed(26070, LUT_AMPL_WIDTH),
		23173 => to_signed(26068, LUT_AMPL_WIDTH),
		23174 => to_signed(26066, LUT_AMPL_WIDTH),
		23175 => to_signed(26064, LUT_AMPL_WIDTH),
		23176 => to_signed(26062, LUT_AMPL_WIDTH),
		23177 => to_signed(26060, LUT_AMPL_WIDTH),
		23178 => to_signed(26058, LUT_AMPL_WIDTH),
		23179 => to_signed(26056, LUT_AMPL_WIDTH),
		23180 => to_signed(26054, LUT_AMPL_WIDTH),
		23181 => to_signed(26052, LUT_AMPL_WIDTH),
		23182 => to_signed(26051, LUT_AMPL_WIDTH),
		23183 => to_signed(26049, LUT_AMPL_WIDTH),
		23184 => to_signed(26047, LUT_AMPL_WIDTH),
		23185 => to_signed(26045, LUT_AMPL_WIDTH),
		23186 => to_signed(26043, LUT_AMPL_WIDTH),
		23187 => to_signed(26041, LUT_AMPL_WIDTH),
		23188 => to_signed(26039, LUT_AMPL_WIDTH),
		23189 => to_signed(26037, LUT_AMPL_WIDTH),
		23190 => to_signed(26035, LUT_AMPL_WIDTH),
		23191 => to_signed(26033, LUT_AMPL_WIDTH),
		23192 => to_signed(26031, LUT_AMPL_WIDTH),
		23193 => to_signed(26030, LUT_AMPL_WIDTH),
		23194 => to_signed(26028, LUT_AMPL_WIDTH),
		23195 => to_signed(26026, LUT_AMPL_WIDTH),
		23196 => to_signed(26024, LUT_AMPL_WIDTH),
		23197 => to_signed(26022, LUT_AMPL_WIDTH),
		23198 => to_signed(26020, LUT_AMPL_WIDTH),
		23199 => to_signed(26018, LUT_AMPL_WIDTH),
		23200 => to_signed(26016, LUT_AMPL_WIDTH),
		23201 => to_signed(26014, LUT_AMPL_WIDTH),
		23202 => to_signed(26012, LUT_AMPL_WIDTH),
		23203 => to_signed(26010, LUT_AMPL_WIDTH),
		23204 => to_signed(26009, LUT_AMPL_WIDTH),
		23205 => to_signed(26007, LUT_AMPL_WIDTH),
		23206 => to_signed(26005, LUT_AMPL_WIDTH),
		23207 => to_signed(26003, LUT_AMPL_WIDTH),
		23208 => to_signed(26001, LUT_AMPL_WIDTH),
		23209 => to_signed(25999, LUT_AMPL_WIDTH),
		23210 => to_signed(25997, LUT_AMPL_WIDTH),
		23211 => to_signed(25995, LUT_AMPL_WIDTH),
		23212 => to_signed(25993, LUT_AMPL_WIDTH),
		23213 => to_signed(25991, LUT_AMPL_WIDTH),
		23214 => to_signed(25989, LUT_AMPL_WIDTH),
		23215 => to_signed(25988, LUT_AMPL_WIDTH),
		23216 => to_signed(25986, LUT_AMPL_WIDTH),
		23217 => to_signed(25984, LUT_AMPL_WIDTH),
		23218 => to_signed(25982, LUT_AMPL_WIDTH),
		23219 => to_signed(25980, LUT_AMPL_WIDTH),
		23220 => to_signed(25978, LUT_AMPL_WIDTH),
		23221 => to_signed(25976, LUT_AMPL_WIDTH),
		23222 => to_signed(25974, LUT_AMPL_WIDTH),
		23223 => to_signed(25972, LUT_AMPL_WIDTH),
		23224 => to_signed(25970, LUT_AMPL_WIDTH),
		23225 => to_signed(25968, LUT_AMPL_WIDTH),
		23226 => to_signed(25966, LUT_AMPL_WIDTH),
		23227 => to_signed(25965, LUT_AMPL_WIDTH),
		23228 => to_signed(25963, LUT_AMPL_WIDTH),
		23229 => to_signed(25961, LUT_AMPL_WIDTH),
		23230 => to_signed(25959, LUT_AMPL_WIDTH),
		23231 => to_signed(25957, LUT_AMPL_WIDTH),
		23232 => to_signed(25955, LUT_AMPL_WIDTH),
		23233 => to_signed(25953, LUT_AMPL_WIDTH),
		23234 => to_signed(25951, LUT_AMPL_WIDTH),
		23235 => to_signed(25949, LUT_AMPL_WIDTH),
		23236 => to_signed(25947, LUT_AMPL_WIDTH),
		23237 => to_signed(25945, LUT_AMPL_WIDTH),
		23238 => to_signed(25943, LUT_AMPL_WIDTH),
		23239 => to_signed(25942, LUT_AMPL_WIDTH),
		23240 => to_signed(25940, LUT_AMPL_WIDTH),
		23241 => to_signed(25938, LUT_AMPL_WIDTH),
		23242 => to_signed(25936, LUT_AMPL_WIDTH),
		23243 => to_signed(25934, LUT_AMPL_WIDTH),
		23244 => to_signed(25932, LUT_AMPL_WIDTH),
		23245 => to_signed(25930, LUT_AMPL_WIDTH),
		23246 => to_signed(25928, LUT_AMPL_WIDTH),
		23247 => to_signed(25926, LUT_AMPL_WIDTH),
		23248 => to_signed(25924, LUT_AMPL_WIDTH),
		23249 => to_signed(25922, LUT_AMPL_WIDTH),
		23250 => to_signed(25920, LUT_AMPL_WIDTH),
		23251 => to_signed(25918, LUT_AMPL_WIDTH),
		23252 => to_signed(25917, LUT_AMPL_WIDTH),
		23253 => to_signed(25915, LUT_AMPL_WIDTH),
		23254 => to_signed(25913, LUT_AMPL_WIDTH),
		23255 => to_signed(25911, LUT_AMPL_WIDTH),
		23256 => to_signed(25909, LUT_AMPL_WIDTH),
		23257 => to_signed(25907, LUT_AMPL_WIDTH),
		23258 => to_signed(25905, LUT_AMPL_WIDTH),
		23259 => to_signed(25903, LUT_AMPL_WIDTH),
		23260 => to_signed(25901, LUT_AMPL_WIDTH),
		23261 => to_signed(25899, LUT_AMPL_WIDTH),
		23262 => to_signed(25897, LUT_AMPL_WIDTH),
		23263 => to_signed(25895, LUT_AMPL_WIDTH),
		23264 => to_signed(25893, LUT_AMPL_WIDTH),
		23265 => to_signed(25892, LUT_AMPL_WIDTH),
		23266 => to_signed(25890, LUT_AMPL_WIDTH),
		23267 => to_signed(25888, LUT_AMPL_WIDTH),
		23268 => to_signed(25886, LUT_AMPL_WIDTH),
		23269 => to_signed(25884, LUT_AMPL_WIDTH),
		23270 => to_signed(25882, LUT_AMPL_WIDTH),
		23271 => to_signed(25880, LUT_AMPL_WIDTH),
		23272 => to_signed(25878, LUT_AMPL_WIDTH),
		23273 => to_signed(25876, LUT_AMPL_WIDTH),
		23274 => to_signed(25874, LUT_AMPL_WIDTH),
		23275 => to_signed(25872, LUT_AMPL_WIDTH),
		23276 => to_signed(25870, LUT_AMPL_WIDTH),
		23277 => to_signed(25868, LUT_AMPL_WIDTH),
		23278 => to_signed(25866, LUT_AMPL_WIDTH),
		23279 => to_signed(25865, LUT_AMPL_WIDTH),
		23280 => to_signed(25863, LUT_AMPL_WIDTH),
		23281 => to_signed(25861, LUT_AMPL_WIDTH),
		23282 => to_signed(25859, LUT_AMPL_WIDTH),
		23283 => to_signed(25857, LUT_AMPL_WIDTH),
		23284 => to_signed(25855, LUT_AMPL_WIDTH),
		23285 => to_signed(25853, LUT_AMPL_WIDTH),
		23286 => to_signed(25851, LUT_AMPL_WIDTH),
		23287 => to_signed(25849, LUT_AMPL_WIDTH),
		23288 => to_signed(25847, LUT_AMPL_WIDTH),
		23289 => to_signed(25845, LUT_AMPL_WIDTH),
		23290 => to_signed(25843, LUT_AMPL_WIDTH),
		23291 => to_signed(25841, LUT_AMPL_WIDTH),
		23292 => to_signed(25839, LUT_AMPL_WIDTH),
		23293 => to_signed(25838, LUT_AMPL_WIDTH),
		23294 => to_signed(25836, LUT_AMPL_WIDTH),
		23295 => to_signed(25834, LUT_AMPL_WIDTH),
		23296 => to_signed(25832, LUT_AMPL_WIDTH),
		23297 => to_signed(25830, LUT_AMPL_WIDTH),
		23298 => to_signed(25828, LUT_AMPL_WIDTH),
		23299 => to_signed(25826, LUT_AMPL_WIDTH),
		23300 => to_signed(25824, LUT_AMPL_WIDTH),
		23301 => to_signed(25822, LUT_AMPL_WIDTH),
		23302 => to_signed(25820, LUT_AMPL_WIDTH),
		23303 => to_signed(25818, LUT_AMPL_WIDTH),
		23304 => to_signed(25816, LUT_AMPL_WIDTH),
		23305 => to_signed(25814, LUT_AMPL_WIDTH),
		23306 => to_signed(25812, LUT_AMPL_WIDTH),
		23307 => to_signed(25810, LUT_AMPL_WIDTH),
		23308 => to_signed(25809, LUT_AMPL_WIDTH),
		23309 => to_signed(25807, LUT_AMPL_WIDTH),
		23310 => to_signed(25805, LUT_AMPL_WIDTH),
		23311 => to_signed(25803, LUT_AMPL_WIDTH),
		23312 => to_signed(25801, LUT_AMPL_WIDTH),
		23313 => to_signed(25799, LUT_AMPL_WIDTH),
		23314 => to_signed(25797, LUT_AMPL_WIDTH),
		23315 => to_signed(25795, LUT_AMPL_WIDTH),
		23316 => to_signed(25793, LUT_AMPL_WIDTH),
		23317 => to_signed(25791, LUT_AMPL_WIDTH),
		23318 => to_signed(25789, LUT_AMPL_WIDTH),
		23319 => to_signed(25787, LUT_AMPL_WIDTH),
		23320 => to_signed(25785, LUT_AMPL_WIDTH),
		23321 => to_signed(25783, LUT_AMPL_WIDTH),
		23322 => to_signed(25781, LUT_AMPL_WIDTH),
		23323 => to_signed(25779, LUT_AMPL_WIDTH),
		23324 => to_signed(25778, LUT_AMPL_WIDTH),
		23325 => to_signed(25776, LUT_AMPL_WIDTH),
		23326 => to_signed(25774, LUT_AMPL_WIDTH),
		23327 => to_signed(25772, LUT_AMPL_WIDTH),
		23328 => to_signed(25770, LUT_AMPL_WIDTH),
		23329 => to_signed(25768, LUT_AMPL_WIDTH),
		23330 => to_signed(25766, LUT_AMPL_WIDTH),
		23331 => to_signed(25764, LUT_AMPL_WIDTH),
		23332 => to_signed(25762, LUT_AMPL_WIDTH),
		23333 => to_signed(25760, LUT_AMPL_WIDTH),
		23334 => to_signed(25758, LUT_AMPL_WIDTH),
		23335 => to_signed(25756, LUT_AMPL_WIDTH),
		23336 => to_signed(25754, LUT_AMPL_WIDTH),
		23337 => to_signed(25752, LUT_AMPL_WIDTH),
		23338 => to_signed(25750, LUT_AMPL_WIDTH),
		23339 => to_signed(25748, LUT_AMPL_WIDTH),
		23340 => to_signed(25746, LUT_AMPL_WIDTH),
		23341 => to_signed(25745, LUT_AMPL_WIDTH),
		23342 => to_signed(25743, LUT_AMPL_WIDTH),
		23343 => to_signed(25741, LUT_AMPL_WIDTH),
		23344 => to_signed(25739, LUT_AMPL_WIDTH),
		23345 => to_signed(25737, LUT_AMPL_WIDTH),
		23346 => to_signed(25735, LUT_AMPL_WIDTH),
		23347 => to_signed(25733, LUT_AMPL_WIDTH),
		23348 => to_signed(25731, LUT_AMPL_WIDTH),
		23349 => to_signed(25729, LUT_AMPL_WIDTH),
		23350 => to_signed(25727, LUT_AMPL_WIDTH),
		23351 => to_signed(25725, LUT_AMPL_WIDTH),
		23352 => to_signed(25723, LUT_AMPL_WIDTH),
		23353 => to_signed(25721, LUT_AMPL_WIDTH),
		23354 => to_signed(25719, LUT_AMPL_WIDTH),
		23355 => to_signed(25717, LUT_AMPL_WIDTH),
		23356 => to_signed(25715, LUT_AMPL_WIDTH),
		23357 => to_signed(25713, LUT_AMPL_WIDTH),
		23358 => to_signed(25711, LUT_AMPL_WIDTH),
		23359 => to_signed(25710, LUT_AMPL_WIDTH),
		23360 => to_signed(25708, LUT_AMPL_WIDTH),
		23361 => to_signed(25706, LUT_AMPL_WIDTH),
		23362 => to_signed(25704, LUT_AMPL_WIDTH),
		23363 => to_signed(25702, LUT_AMPL_WIDTH),
		23364 => to_signed(25700, LUT_AMPL_WIDTH),
		23365 => to_signed(25698, LUT_AMPL_WIDTH),
		23366 => to_signed(25696, LUT_AMPL_WIDTH),
		23367 => to_signed(25694, LUT_AMPL_WIDTH),
		23368 => to_signed(25692, LUT_AMPL_WIDTH),
		23369 => to_signed(25690, LUT_AMPL_WIDTH),
		23370 => to_signed(25688, LUT_AMPL_WIDTH),
		23371 => to_signed(25686, LUT_AMPL_WIDTH),
		23372 => to_signed(25684, LUT_AMPL_WIDTH),
		23373 => to_signed(25682, LUT_AMPL_WIDTH),
		23374 => to_signed(25680, LUT_AMPL_WIDTH),
		23375 => to_signed(25678, LUT_AMPL_WIDTH),
		23376 => to_signed(25676, LUT_AMPL_WIDTH),
		23377 => to_signed(25674, LUT_AMPL_WIDTH),
		23378 => to_signed(25672, LUT_AMPL_WIDTH),
		23379 => to_signed(25671, LUT_AMPL_WIDTH),
		23380 => to_signed(25669, LUT_AMPL_WIDTH),
		23381 => to_signed(25667, LUT_AMPL_WIDTH),
		23382 => to_signed(25665, LUT_AMPL_WIDTH),
		23383 => to_signed(25663, LUT_AMPL_WIDTH),
		23384 => to_signed(25661, LUT_AMPL_WIDTH),
		23385 => to_signed(25659, LUT_AMPL_WIDTH),
		23386 => to_signed(25657, LUT_AMPL_WIDTH),
		23387 => to_signed(25655, LUT_AMPL_WIDTH),
		23388 => to_signed(25653, LUT_AMPL_WIDTH),
		23389 => to_signed(25651, LUT_AMPL_WIDTH),
		23390 => to_signed(25649, LUT_AMPL_WIDTH),
		23391 => to_signed(25647, LUT_AMPL_WIDTH),
		23392 => to_signed(25645, LUT_AMPL_WIDTH),
		23393 => to_signed(25643, LUT_AMPL_WIDTH),
		23394 => to_signed(25641, LUT_AMPL_WIDTH),
		23395 => to_signed(25639, LUT_AMPL_WIDTH),
		23396 => to_signed(25637, LUT_AMPL_WIDTH),
		23397 => to_signed(25635, LUT_AMPL_WIDTH),
		23398 => to_signed(25633, LUT_AMPL_WIDTH),
		23399 => to_signed(25631, LUT_AMPL_WIDTH),
		23400 => to_signed(25629, LUT_AMPL_WIDTH),
		23401 => to_signed(25628, LUT_AMPL_WIDTH),
		23402 => to_signed(25626, LUT_AMPL_WIDTH),
		23403 => to_signed(25624, LUT_AMPL_WIDTH),
		23404 => to_signed(25622, LUT_AMPL_WIDTH),
		23405 => to_signed(25620, LUT_AMPL_WIDTH),
		23406 => to_signed(25618, LUT_AMPL_WIDTH),
		23407 => to_signed(25616, LUT_AMPL_WIDTH),
		23408 => to_signed(25614, LUT_AMPL_WIDTH),
		23409 => to_signed(25612, LUT_AMPL_WIDTH),
		23410 => to_signed(25610, LUT_AMPL_WIDTH),
		23411 => to_signed(25608, LUT_AMPL_WIDTH),
		23412 => to_signed(25606, LUT_AMPL_WIDTH),
		23413 => to_signed(25604, LUT_AMPL_WIDTH),
		23414 => to_signed(25602, LUT_AMPL_WIDTH),
		23415 => to_signed(25600, LUT_AMPL_WIDTH),
		23416 => to_signed(25598, LUT_AMPL_WIDTH),
		23417 => to_signed(25596, LUT_AMPL_WIDTH),
		23418 => to_signed(25594, LUT_AMPL_WIDTH),
		23419 => to_signed(25592, LUT_AMPL_WIDTH),
		23420 => to_signed(25590, LUT_AMPL_WIDTH),
		23421 => to_signed(25588, LUT_AMPL_WIDTH),
		23422 => to_signed(25586, LUT_AMPL_WIDTH),
		23423 => to_signed(25584, LUT_AMPL_WIDTH),
		23424 => to_signed(25582, LUT_AMPL_WIDTH),
		23425 => to_signed(25580, LUT_AMPL_WIDTH),
		23426 => to_signed(25578, LUT_AMPL_WIDTH),
		23427 => to_signed(25577, LUT_AMPL_WIDTH),
		23428 => to_signed(25575, LUT_AMPL_WIDTH),
		23429 => to_signed(25573, LUT_AMPL_WIDTH),
		23430 => to_signed(25571, LUT_AMPL_WIDTH),
		23431 => to_signed(25569, LUT_AMPL_WIDTH),
		23432 => to_signed(25567, LUT_AMPL_WIDTH),
		23433 => to_signed(25565, LUT_AMPL_WIDTH),
		23434 => to_signed(25563, LUT_AMPL_WIDTH),
		23435 => to_signed(25561, LUT_AMPL_WIDTH),
		23436 => to_signed(25559, LUT_AMPL_WIDTH),
		23437 => to_signed(25557, LUT_AMPL_WIDTH),
		23438 => to_signed(25555, LUT_AMPL_WIDTH),
		23439 => to_signed(25553, LUT_AMPL_WIDTH),
		23440 => to_signed(25551, LUT_AMPL_WIDTH),
		23441 => to_signed(25549, LUT_AMPL_WIDTH),
		23442 => to_signed(25547, LUT_AMPL_WIDTH),
		23443 => to_signed(25545, LUT_AMPL_WIDTH),
		23444 => to_signed(25543, LUT_AMPL_WIDTH),
		23445 => to_signed(25541, LUT_AMPL_WIDTH),
		23446 => to_signed(25539, LUT_AMPL_WIDTH),
		23447 => to_signed(25537, LUT_AMPL_WIDTH),
		23448 => to_signed(25535, LUT_AMPL_WIDTH),
		23449 => to_signed(25533, LUT_AMPL_WIDTH),
		23450 => to_signed(25531, LUT_AMPL_WIDTH),
		23451 => to_signed(25529, LUT_AMPL_WIDTH),
		23452 => to_signed(25527, LUT_AMPL_WIDTH),
		23453 => to_signed(25525, LUT_AMPL_WIDTH),
		23454 => to_signed(25523, LUT_AMPL_WIDTH),
		23455 => to_signed(25521, LUT_AMPL_WIDTH),
		23456 => to_signed(25519, LUT_AMPL_WIDTH),
		23457 => to_signed(25518, LUT_AMPL_WIDTH),
		23458 => to_signed(25516, LUT_AMPL_WIDTH),
		23459 => to_signed(25514, LUT_AMPL_WIDTH),
		23460 => to_signed(25512, LUT_AMPL_WIDTH),
		23461 => to_signed(25510, LUT_AMPL_WIDTH),
		23462 => to_signed(25508, LUT_AMPL_WIDTH),
		23463 => to_signed(25506, LUT_AMPL_WIDTH),
		23464 => to_signed(25504, LUT_AMPL_WIDTH),
		23465 => to_signed(25502, LUT_AMPL_WIDTH),
		23466 => to_signed(25500, LUT_AMPL_WIDTH),
		23467 => to_signed(25498, LUT_AMPL_WIDTH),
		23468 => to_signed(25496, LUT_AMPL_WIDTH),
		23469 => to_signed(25494, LUT_AMPL_WIDTH),
		23470 => to_signed(25492, LUT_AMPL_WIDTH),
		23471 => to_signed(25490, LUT_AMPL_WIDTH),
		23472 => to_signed(25488, LUT_AMPL_WIDTH),
		23473 => to_signed(25486, LUT_AMPL_WIDTH),
		23474 => to_signed(25484, LUT_AMPL_WIDTH),
		23475 => to_signed(25482, LUT_AMPL_WIDTH),
		23476 => to_signed(25480, LUT_AMPL_WIDTH),
		23477 => to_signed(25478, LUT_AMPL_WIDTH),
		23478 => to_signed(25476, LUT_AMPL_WIDTH),
		23479 => to_signed(25474, LUT_AMPL_WIDTH),
		23480 => to_signed(25472, LUT_AMPL_WIDTH),
		23481 => to_signed(25470, LUT_AMPL_WIDTH),
		23482 => to_signed(25468, LUT_AMPL_WIDTH),
		23483 => to_signed(25466, LUT_AMPL_WIDTH),
		23484 => to_signed(25464, LUT_AMPL_WIDTH),
		23485 => to_signed(25462, LUT_AMPL_WIDTH),
		23486 => to_signed(25460, LUT_AMPL_WIDTH),
		23487 => to_signed(25458, LUT_AMPL_WIDTH),
		23488 => to_signed(25456, LUT_AMPL_WIDTH),
		23489 => to_signed(25454, LUT_AMPL_WIDTH),
		23490 => to_signed(25452, LUT_AMPL_WIDTH),
		23491 => to_signed(25450, LUT_AMPL_WIDTH),
		23492 => to_signed(25448, LUT_AMPL_WIDTH),
		23493 => to_signed(25446, LUT_AMPL_WIDTH),
		23494 => to_signed(25444, LUT_AMPL_WIDTH),
		23495 => to_signed(25442, LUT_AMPL_WIDTH),
		23496 => to_signed(25440, LUT_AMPL_WIDTH),
		23497 => to_signed(25438, LUT_AMPL_WIDTH),
		23498 => to_signed(25437, LUT_AMPL_WIDTH),
		23499 => to_signed(25435, LUT_AMPL_WIDTH),
		23500 => to_signed(25433, LUT_AMPL_WIDTH),
		23501 => to_signed(25431, LUT_AMPL_WIDTH),
		23502 => to_signed(25429, LUT_AMPL_WIDTH),
		23503 => to_signed(25427, LUT_AMPL_WIDTH),
		23504 => to_signed(25425, LUT_AMPL_WIDTH),
		23505 => to_signed(25423, LUT_AMPL_WIDTH),
		23506 => to_signed(25421, LUT_AMPL_WIDTH),
		23507 => to_signed(25419, LUT_AMPL_WIDTH),
		23508 => to_signed(25417, LUT_AMPL_WIDTH),
		23509 => to_signed(25415, LUT_AMPL_WIDTH),
		23510 => to_signed(25413, LUT_AMPL_WIDTH),
		23511 => to_signed(25411, LUT_AMPL_WIDTH),
		23512 => to_signed(25409, LUT_AMPL_WIDTH),
		23513 => to_signed(25407, LUT_AMPL_WIDTH),
		23514 => to_signed(25405, LUT_AMPL_WIDTH),
		23515 => to_signed(25403, LUT_AMPL_WIDTH),
		23516 => to_signed(25401, LUT_AMPL_WIDTH),
		23517 => to_signed(25399, LUT_AMPL_WIDTH),
		23518 => to_signed(25397, LUT_AMPL_WIDTH),
		23519 => to_signed(25395, LUT_AMPL_WIDTH),
		23520 => to_signed(25393, LUT_AMPL_WIDTH),
		23521 => to_signed(25391, LUT_AMPL_WIDTH),
		23522 => to_signed(25389, LUT_AMPL_WIDTH),
		23523 => to_signed(25387, LUT_AMPL_WIDTH),
		23524 => to_signed(25385, LUT_AMPL_WIDTH),
		23525 => to_signed(25383, LUT_AMPL_WIDTH),
		23526 => to_signed(25381, LUT_AMPL_WIDTH),
		23527 => to_signed(25379, LUT_AMPL_WIDTH),
		23528 => to_signed(25377, LUT_AMPL_WIDTH),
		23529 => to_signed(25375, LUT_AMPL_WIDTH),
		23530 => to_signed(25373, LUT_AMPL_WIDTH),
		23531 => to_signed(25371, LUT_AMPL_WIDTH),
		23532 => to_signed(25369, LUT_AMPL_WIDTH),
		23533 => to_signed(25367, LUT_AMPL_WIDTH),
		23534 => to_signed(25365, LUT_AMPL_WIDTH),
		23535 => to_signed(25363, LUT_AMPL_WIDTH),
		23536 => to_signed(25361, LUT_AMPL_WIDTH),
		23537 => to_signed(25359, LUT_AMPL_WIDTH),
		23538 => to_signed(25357, LUT_AMPL_WIDTH),
		23539 => to_signed(25355, LUT_AMPL_WIDTH),
		23540 => to_signed(25353, LUT_AMPL_WIDTH),
		23541 => to_signed(25351, LUT_AMPL_WIDTH),
		23542 => to_signed(25349, LUT_AMPL_WIDTH),
		23543 => to_signed(25347, LUT_AMPL_WIDTH),
		23544 => to_signed(25345, LUT_AMPL_WIDTH),
		23545 => to_signed(25343, LUT_AMPL_WIDTH),
		23546 => to_signed(25341, LUT_AMPL_WIDTH),
		23547 => to_signed(25339, LUT_AMPL_WIDTH),
		23548 => to_signed(25337, LUT_AMPL_WIDTH),
		23549 => to_signed(25335, LUT_AMPL_WIDTH),
		23550 => to_signed(25333, LUT_AMPL_WIDTH),
		23551 => to_signed(25331, LUT_AMPL_WIDTH),
		23552 => to_signed(25329, LUT_AMPL_WIDTH),
		23553 => to_signed(25327, LUT_AMPL_WIDTH),
		23554 => to_signed(25325, LUT_AMPL_WIDTH),
		23555 => to_signed(25323, LUT_AMPL_WIDTH),
		23556 => to_signed(25321, LUT_AMPL_WIDTH),
		23557 => to_signed(25319, LUT_AMPL_WIDTH),
		23558 => to_signed(25317, LUT_AMPL_WIDTH),
		23559 => to_signed(25315, LUT_AMPL_WIDTH),
		23560 => to_signed(25313, LUT_AMPL_WIDTH),
		23561 => to_signed(25311, LUT_AMPL_WIDTH),
		23562 => to_signed(25309, LUT_AMPL_WIDTH),
		23563 => to_signed(25307, LUT_AMPL_WIDTH),
		23564 => to_signed(25305, LUT_AMPL_WIDTH),
		23565 => to_signed(25303, LUT_AMPL_WIDTH),
		23566 => to_signed(25301, LUT_AMPL_WIDTH),
		23567 => to_signed(25299, LUT_AMPL_WIDTH),
		23568 => to_signed(25297, LUT_AMPL_WIDTH),
		23569 => to_signed(25295, LUT_AMPL_WIDTH),
		23570 => to_signed(25293, LUT_AMPL_WIDTH),
		23571 => to_signed(25291, LUT_AMPL_WIDTH),
		23572 => to_signed(25289, LUT_AMPL_WIDTH),
		23573 => to_signed(25287, LUT_AMPL_WIDTH),
		23574 => to_signed(25285, LUT_AMPL_WIDTH),
		23575 => to_signed(25283, LUT_AMPL_WIDTH),
		23576 => to_signed(25281, LUT_AMPL_WIDTH),
		23577 => to_signed(25279, LUT_AMPL_WIDTH),
		23578 => to_signed(25277, LUT_AMPL_WIDTH),
		23579 => to_signed(25275, LUT_AMPL_WIDTH),
		23580 => to_signed(25273, LUT_AMPL_WIDTH),
		23581 => to_signed(25271, LUT_AMPL_WIDTH),
		23582 => to_signed(25269, LUT_AMPL_WIDTH),
		23583 => to_signed(25267, LUT_AMPL_WIDTH),
		23584 => to_signed(25265, LUT_AMPL_WIDTH),
		23585 => to_signed(25263, LUT_AMPL_WIDTH),
		23586 => to_signed(25261, LUT_AMPL_WIDTH),
		23587 => to_signed(25259, LUT_AMPL_WIDTH),
		23588 => to_signed(25257, LUT_AMPL_WIDTH),
		23589 => to_signed(25255, LUT_AMPL_WIDTH),
		23590 => to_signed(25253, LUT_AMPL_WIDTH),
		23591 => to_signed(25251, LUT_AMPL_WIDTH),
		23592 => to_signed(25249, LUT_AMPL_WIDTH),
		23593 => to_signed(25247, LUT_AMPL_WIDTH),
		23594 => to_signed(25245, LUT_AMPL_WIDTH),
		23595 => to_signed(25243, LUT_AMPL_WIDTH),
		23596 => to_signed(25241, LUT_AMPL_WIDTH),
		23597 => to_signed(25239, LUT_AMPL_WIDTH),
		23598 => to_signed(25237, LUT_AMPL_WIDTH),
		23599 => to_signed(25235, LUT_AMPL_WIDTH),
		23600 => to_signed(25233, LUT_AMPL_WIDTH),
		23601 => to_signed(25231, LUT_AMPL_WIDTH),
		23602 => to_signed(25229, LUT_AMPL_WIDTH),
		23603 => to_signed(25227, LUT_AMPL_WIDTH),
		23604 => to_signed(25225, LUT_AMPL_WIDTH),
		23605 => to_signed(25223, LUT_AMPL_WIDTH),
		23606 => to_signed(25221, LUT_AMPL_WIDTH),
		23607 => to_signed(25219, LUT_AMPL_WIDTH),
		23608 => to_signed(25217, LUT_AMPL_WIDTH),
		23609 => to_signed(25215, LUT_AMPL_WIDTH),
		23610 => to_signed(25213, LUT_AMPL_WIDTH),
		23611 => to_signed(25211, LUT_AMPL_WIDTH),
		23612 => to_signed(25209, LUT_AMPL_WIDTH),
		23613 => to_signed(25207, LUT_AMPL_WIDTH),
		23614 => to_signed(25205, LUT_AMPL_WIDTH),
		23615 => to_signed(25203, LUT_AMPL_WIDTH),
		23616 => to_signed(25201, LUT_AMPL_WIDTH),
		23617 => to_signed(25199, LUT_AMPL_WIDTH),
		23618 => to_signed(25197, LUT_AMPL_WIDTH),
		23619 => to_signed(25195, LUT_AMPL_WIDTH),
		23620 => to_signed(25193, LUT_AMPL_WIDTH),
		23621 => to_signed(25191, LUT_AMPL_WIDTH),
		23622 => to_signed(25189, LUT_AMPL_WIDTH),
		23623 => to_signed(25187, LUT_AMPL_WIDTH),
		23624 => to_signed(25185, LUT_AMPL_WIDTH),
		23625 => to_signed(25183, LUT_AMPL_WIDTH),
		23626 => to_signed(25181, LUT_AMPL_WIDTH),
		23627 => to_signed(25179, LUT_AMPL_WIDTH),
		23628 => to_signed(25177, LUT_AMPL_WIDTH),
		23629 => to_signed(25175, LUT_AMPL_WIDTH),
		23630 => to_signed(25173, LUT_AMPL_WIDTH),
		23631 => to_signed(25171, LUT_AMPL_WIDTH),
		23632 => to_signed(25169, LUT_AMPL_WIDTH),
		23633 => to_signed(25167, LUT_AMPL_WIDTH),
		23634 => to_signed(25165, LUT_AMPL_WIDTH),
		23635 => to_signed(25163, LUT_AMPL_WIDTH),
		23636 => to_signed(25161, LUT_AMPL_WIDTH),
		23637 => to_signed(25159, LUT_AMPL_WIDTH),
		23638 => to_signed(25157, LUT_AMPL_WIDTH),
		23639 => to_signed(25155, LUT_AMPL_WIDTH),
		23640 => to_signed(25153, LUT_AMPL_WIDTH),
		23641 => to_signed(25151, LUT_AMPL_WIDTH),
		23642 => to_signed(25149, LUT_AMPL_WIDTH),
		23643 => to_signed(25147, LUT_AMPL_WIDTH),
		23644 => to_signed(25145, LUT_AMPL_WIDTH),
		23645 => to_signed(25143, LUT_AMPL_WIDTH),
		23646 => to_signed(25141, LUT_AMPL_WIDTH),
		23647 => to_signed(25139, LUT_AMPL_WIDTH),
		23648 => to_signed(25137, LUT_AMPL_WIDTH),
		23649 => to_signed(25135, LUT_AMPL_WIDTH),
		23650 => to_signed(25133, LUT_AMPL_WIDTH),
		23651 => to_signed(25131, LUT_AMPL_WIDTH),
		23652 => to_signed(25129, LUT_AMPL_WIDTH),
		23653 => to_signed(25127, LUT_AMPL_WIDTH),
		23654 => to_signed(25125, LUT_AMPL_WIDTH),
		23655 => to_signed(25123, LUT_AMPL_WIDTH),
		23656 => to_signed(25121, LUT_AMPL_WIDTH),
		23657 => to_signed(25119, LUT_AMPL_WIDTH),
		23658 => to_signed(25117, LUT_AMPL_WIDTH),
		23659 => to_signed(25115, LUT_AMPL_WIDTH),
		23660 => to_signed(25113, LUT_AMPL_WIDTH),
		23661 => to_signed(25111, LUT_AMPL_WIDTH),
		23662 => to_signed(25109, LUT_AMPL_WIDTH),
		23663 => to_signed(25107, LUT_AMPL_WIDTH),
		23664 => to_signed(25105, LUT_AMPL_WIDTH),
		23665 => to_signed(25103, LUT_AMPL_WIDTH),
		23666 => to_signed(25101, LUT_AMPL_WIDTH),
		23667 => to_signed(25099, LUT_AMPL_WIDTH),
		23668 => to_signed(25096, LUT_AMPL_WIDTH),
		23669 => to_signed(25094, LUT_AMPL_WIDTH),
		23670 => to_signed(25092, LUT_AMPL_WIDTH),
		23671 => to_signed(25090, LUT_AMPL_WIDTH),
		23672 => to_signed(25088, LUT_AMPL_WIDTH),
		23673 => to_signed(25086, LUT_AMPL_WIDTH),
		23674 => to_signed(25084, LUT_AMPL_WIDTH),
		23675 => to_signed(25082, LUT_AMPL_WIDTH),
		23676 => to_signed(25080, LUT_AMPL_WIDTH),
		23677 => to_signed(25078, LUT_AMPL_WIDTH),
		23678 => to_signed(25076, LUT_AMPL_WIDTH),
		23679 => to_signed(25074, LUT_AMPL_WIDTH),
		23680 => to_signed(25072, LUT_AMPL_WIDTH),
		23681 => to_signed(25070, LUT_AMPL_WIDTH),
		23682 => to_signed(25068, LUT_AMPL_WIDTH),
		23683 => to_signed(25066, LUT_AMPL_WIDTH),
		23684 => to_signed(25064, LUT_AMPL_WIDTH),
		23685 => to_signed(25062, LUT_AMPL_WIDTH),
		23686 => to_signed(25060, LUT_AMPL_WIDTH),
		23687 => to_signed(25058, LUT_AMPL_WIDTH),
		23688 => to_signed(25056, LUT_AMPL_WIDTH),
		23689 => to_signed(25054, LUT_AMPL_WIDTH),
		23690 => to_signed(25052, LUT_AMPL_WIDTH),
		23691 => to_signed(25050, LUT_AMPL_WIDTH),
		23692 => to_signed(25048, LUT_AMPL_WIDTH),
		23693 => to_signed(25046, LUT_AMPL_WIDTH),
		23694 => to_signed(25044, LUT_AMPL_WIDTH),
		23695 => to_signed(25042, LUT_AMPL_WIDTH),
		23696 => to_signed(25040, LUT_AMPL_WIDTH),
		23697 => to_signed(25038, LUT_AMPL_WIDTH),
		23698 => to_signed(25036, LUT_AMPL_WIDTH),
		23699 => to_signed(25034, LUT_AMPL_WIDTH),
		23700 => to_signed(25032, LUT_AMPL_WIDTH),
		23701 => to_signed(25030, LUT_AMPL_WIDTH),
		23702 => to_signed(25028, LUT_AMPL_WIDTH),
		23703 => to_signed(25026, LUT_AMPL_WIDTH),
		23704 => to_signed(25024, LUT_AMPL_WIDTH),
		23705 => to_signed(25022, LUT_AMPL_WIDTH),
		23706 => to_signed(25020, LUT_AMPL_WIDTH),
		23707 => to_signed(25018, LUT_AMPL_WIDTH),
		23708 => to_signed(25016, LUT_AMPL_WIDTH),
		23709 => to_signed(25013, LUT_AMPL_WIDTH),
		23710 => to_signed(25011, LUT_AMPL_WIDTH),
		23711 => to_signed(25009, LUT_AMPL_WIDTH),
		23712 => to_signed(25007, LUT_AMPL_WIDTH),
		23713 => to_signed(25005, LUT_AMPL_WIDTH),
		23714 => to_signed(25003, LUT_AMPL_WIDTH),
		23715 => to_signed(25001, LUT_AMPL_WIDTH),
		23716 => to_signed(24999, LUT_AMPL_WIDTH),
		23717 => to_signed(24997, LUT_AMPL_WIDTH),
		23718 => to_signed(24995, LUT_AMPL_WIDTH),
		23719 => to_signed(24993, LUT_AMPL_WIDTH),
		23720 => to_signed(24991, LUT_AMPL_WIDTH),
		23721 => to_signed(24989, LUT_AMPL_WIDTH),
		23722 => to_signed(24987, LUT_AMPL_WIDTH),
		23723 => to_signed(24985, LUT_AMPL_WIDTH),
		23724 => to_signed(24983, LUT_AMPL_WIDTH),
		23725 => to_signed(24981, LUT_AMPL_WIDTH),
		23726 => to_signed(24979, LUT_AMPL_WIDTH),
		23727 => to_signed(24977, LUT_AMPL_WIDTH),
		23728 => to_signed(24975, LUT_AMPL_WIDTH),
		23729 => to_signed(24973, LUT_AMPL_WIDTH),
		23730 => to_signed(24971, LUT_AMPL_WIDTH),
		23731 => to_signed(24969, LUT_AMPL_WIDTH),
		23732 => to_signed(24967, LUT_AMPL_WIDTH),
		23733 => to_signed(24965, LUT_AMPL_WIDTH),
		23734 => to_signed(24963, LUT_AMPL_WIDTH),
		23735 => to_signed(24961, LUT_AMPL_WIDTH),
		23736 => to_signed(24959, LUT_AMPL_WIDTH),
		23737 => to_signed(24957, LUT_AMPL_WIDTH),
		23738 => to_signed(24955, LUT_AMPL_WIDTH),
		23739 => to_signed(24953, LUT_AMPL_WIDTH),
		23740 => to_signed(24950, LUT_AMPL_WIDTH),
		23741 => to_signed(24948, LUT_AMPL_WIDTH),
		23742 => to_signed(24946, LUT_AMPL_WIDTH),
		23743 => to_signed(24944, LUT_AMPL_WIDTH),
		23744 => to_signed(24942, LUT_AMPL_WIDTH),
		23745 => to_signed(24940, LUT_AMPL_WIDTH),
		23746 => to_signed(24938, LUT_AMPL_WIDTH),
		23747 => to_signed(24936, LUT_AMPL_WIDTH),
		23748 => to_signed(24934, LUT_AMPL_WIDTH),
		23749 => to_signed(24932, LUT_AMPL_WIDTH),
		23750 => to_signed(24930, LUT_AMPL_WIDTH),
		23751 => to_signed(24928, LUT_AMPL_WIDTH),
		23752 => to_signed(24926, LUT_AMPL_WIDTH),
		23753 => to_signed(24924, LUT_AMPL_WIDTH),
		23754 => to_signed(24922, LUT_AMPL_WIDTH),
		23755 => to_signed(24920, LUT_AMPL_WIDTH),
		23756 => to_signed(24918, LUT_AMPL_WIDTH),
		23757 => to_signed(24916, LUT_AMPL_WIDTH),
		23758 => to_signed(24914, LUT_AMPL_WIDTH),
		23759 => to_signed(24912, LUT_AMPL_WIDTH),
		23760 => to_signed(24910, LUT_AMPL_WIDTH),
		23761 => to_signed(24908, LUT_AMPL_WIDTH),
		23762 => to_signed(24906, LUT_AMPL_WIDTH),
		23763 => to_signed(24904, LUT_AMPL_WIDTH),
		23764 => to_signed(24902, LUT_AMPL_WIDTH),
		23765 => to_signed(24899, LUT_AMPL_WIDTH),
		23766 => to_signed(24897, LUT_AMPL_WIDTH),
		23767 => to_signed(24895, LUT_AMPL_WIDTH),
		23768 => to_signed(24893, LUT_AMPL_WIDTH),
		23769 => to_signed(24891, LUT_AMPL_WIDTH),
		23770 => to_signed(24889, LUT_AMPL_WIDTH),
		23771 => to_signed(24887, LUT_AMPL_WIDTH),
		23772 => to_signed(24885, LUT_AMPL_WIDTH),
		23773 => to_signed(24883, LUT_AMPL_WIDTH),
		23774 => to_signed(24881, LUT_AMPL_WIDTH),
		23775 => to_signed(24879, LUT_AMPL_WIDTH),
		23776 => to_signed(24877, LUT_AMPL_WIDTH),
		23777 => to_signed(24875, LUT_AMPL_WIDTH),
		23778 => to_signed(24873, LUT_AMPL_WIDTH),
		23779 => to_signed(24871, LUT_AMPL_WIDTH),
		23780 => to_signed(24869, LUT_AMPL_WIDTH),
		23781 => to_signed(24867, LUT_AMPL_WIDTH),
		23782 => to_signed(24865, LUT_AMPL_WIDTH),
		23783 => to_signed(24863, LUT_AMPL_WIDTH),
		23784 => to_signed(24861, LUT_AMPL_WIDTH),
		23785 => to_signed(24859, LUT_AMPL_WIDTH),
		23786 => to_signed(24857, LUT_AMPL_WIDTH),
		23787 => to_signed(24855, LUT_AMPL_WIDTH),
		23788 => to_signed(24852, LUT_AMPL_WIDTH),
		23789 => to_signed(24850, LUT_AMPL_WIDTH),
		23790 => to_signed(24848, LUT_AMPL_WIDTH),
		23791 => to_signed(24846, LUT_AMPL_WIDTH),
		23792 => to_signed(24844, LUT_AMPL_WIDTH),
		23793 => to_signed(24842, LUT_AMPL_WIDTH),
		23794 => to_signed(24840, LUT_AMPL_WIDTH),
		23795 => to_signed(24838, LUT_AMPL_WIDTH),
		23796 => to_signed(24836, LUT_AMPL_WIDTH),
		23797 => to_signed(24834, LUT_AMPL_WIDTH),
		23798 => to_signed(24832, LUT_AMPL_WIDTH),
		23799 => to_signed(24830, LUT_AMPL_WIDTH),
		23800 => to_signed(24828, LUT_AMPL_WIDTH),
		23801 => to_signed(24826, LUT_AMPL_WIDTH),
		23802 => to_signed(24824, LUT_AMPL_WIDTH),
		23803 => to_signed(24822, LUT_AMPL_WIDTH),
		23804 => to_signed(24820, LUT_AMPL_WIDTH),
		23805 => to_signed(24818, LUT_AMPL_WIDTH),
		23806 => to_signed(24816, LUT_AMPL_WIDTH),
		23807 => to_signed(24814, LUT_AMPL_WIDTH),
		23808 => to_signed(24811, LUT_AMPL_WIDTH),
		23809 => to_signed(24809, LUT_AMPL_WIDTH),
		23810 => to_signed(24807, LUT_AMPL_WIDTH),
		23811 => to_signed(24805, LUT_AMPL_WIDTH),
		23812 => to_signed(24803, LUT_AMPL_WIDTH),
		23813 => to_signed(24801, LUT_AMPL_WIDTH),
		23814 => to_signed(24799, LUT_AMPL_WIDTH),
		23815 => to_signed(24797, LUT_AMPL_WIDTH),
		23816 => to_signed(24795, LUT_AMPL_WIDTH),
		23817 => to_signed(24793, LUT_AMPL_WIDTH),
		23818 => to_signed(24791, LUT_AMPL_WIDTH),
		23819 => to_signed(24789, LUT_AMPL_WIDTH),
		23820 => to_signed(24787, LUT_AMPL_WIDTH),
		23821 => to_signed(24785, LUT_AMPL_WIDTH),
		23822 => to_signed(24783, LUT_AMPL_WIDTH),
		23823 => to_signed(24781, LUT_AMPL_WIDTH),
		23824 => to_signed(24779, LUT_AMPL_WIDTH),
		23825 => to_signed(24777, LUT_AMPL_WIDTH),
		23826 => to_signed(24774, LUT_AMPL_WIDTH),
		23827 => to_signed(24772, LUT_AMPL_WIDTH),
		23828 => to_signed(24770, LUT_AMPL_WIDTH),
		23829 => to_signed(24768, LUT_AMPL_WIDTH),
		23830 => to_signed(24766, LUT_AMPL_WIDTH),
		23831 => to_signed(24764, LUT_AMPL_WIDTH),
		23832 => to_signed(24762, LUT_AMPL_WIDTH),
		23833 => to_signed(24760, LUT_AMPL_WIDTH),
		23834 => to_signed(24758, LUT_AMPL_WIDTH),
		23835 => to_signed(24756, LUT_AMPL_WIDTH),
		23836 => to_signed(24754, LUT_AMPL_WIDTH),
		23837 => to_signed(24752, LUT_AMPL_WIDTH),
		23838 => to_signed(24750, LUT_AMPL_WIDTH),
		23839 => to_signed(24748, LUT_AMPL_WIDTH),
		23840 => to_signed(24746, LUT_AMPL_WIDTH),
		23841 => to_signed(24744, LUT_AMPL_WIDTH),
		23842 => to_signed(24742, LUT_AMPL_WIDTH),
		23843 => to_signed(24740, LUT_AMPL_WIDTH),
		23844 => to_signed(24737, LUT_AMPL_WIDTH),
		23845 => to_signed(24735, LUT_AMPL_WIDTH),
		23846 => to_signed(24733, LUT_AMPL_WIDTH),
		23847 => to_signed(24731, LUT_AMPL_WIDTH),
		23848 => to_signed(24729, LUT_AMPL_WIDTH),
		23849 => to_signed(24727, LUT_AMPL_WIDTH),
		23850 => to_signed(24725, LUT_AMPL_WIDTH),
		23851 => to_signed(24723, LUT_AMPL_WIDTH),
		23852 => to_signed(24721, LUT_AMPL_WIDTH),
		23853 => to_signed(24719, LUT_AMPL_WIDTH),
		23854 => to_signed(24717, LUT_AMPL_WIDTH),
		23855 => to_signed(24715, LUT_AMPL_WIDTH),
		23856 => to_signed(24713, LUT_AMPL_WIDTH),
		23857 => to_signed(24711, LUT_AMPL_WIDTH),
		23858 => to_signed(24709, LUT_AMPL_WIDTH),
		23859 => to_signed(24707, LUT_AMPL_WIDTH),
		23860 => to_signed(24704, LUT_AMPL_WIDTH),
		23861 => to_signed(24702, LUT_AMPL_WIDTH),
		23862 => to_signed(24700, LUT_AMPL_WIDTH),
		23863 => to_signed(24698, LUT_AMPL_WIDTH),
		23864 => to_signed(24696, LUT_AMPL_WIDTH),
		23865 => to_signed(24694, LUT_AMPL_WIDTH),
		23866 => to_signed(24692, LUT_AMPL_WIDTH),
		23867 => to_signed(24690, LUT_AMPL_WIDTH),
		23868 => to_signed(24688, LUT_AMPL_WIDTH),
		23869 => to_signed(24686, LUT_AMPL_WIDTH),
		23870 => to_signed(24684, LUT_AMPL_WIDTH),
		23871 => to_signed(24682, LUT_AMPL_WIDTH),
		23872 => to_signed(24680, LUT_AMPL_WIDTH),
		23873 => to_signed(24678, LUT_AMPL_WIDTH),
		23874 => to_signed(24676, LUT_AMPL_WIDTH),
		23875 => to_signed(24673, LUT_AMPL_WIDTH),
		23876 => to_signed(24671, LUT_AMPL_WIDTH),
		23877 => to_signed(24669, LUT_AMPL_WIDTH),
		23878 => to_signed(24667, LUT_AMPL_WIDTH),
		23879 => to_signed(24665, LUT_AMPL_WIDTH),
		23880 => to_signed(24663, LUT_AMPL_WIDTH),
		23881 => to_signed(24661, LUT_AMPL_WIDTH),
		23882 => to_signed(24659, LUT_AMPL_WIDTH),
		23883 => to_signed(24657, LUT_AMPL_WIDTH),
		23884 => to_signed(24655, LUT_AMPL_WIDTH),
		23885 => to_signed(24653, LUT_AMPL_WIDTH),
		23886 => to_signed(24651, LUT_AMPL_WIDTH),
		23887 => to_signed(24649, LUT_AMPL_WIDTH),
		23888 => to_signed(24647, LUT_AMPL_WIDTH),
		23889 => to_signed(24645, LUT_AMPL_WIDTH),
		23890 => to_signed(24642, LUT_AMPL_WIDTH),
		23891 => to_signed(24640, LUT_AMPL_WIDTH),
		23892 => to_signed(24638, LUT_AMPL_WIDTH),
		23893 => to_signed(24636, LUT_AMPL_WIDTH),
		23894 => to_signed(24634, LUT_AMPL_WIDTH),
		23895 => to_signed(24632, LUT_AMPL_WIDTH),
		23896 => to_signed(24630, LUT_AMPL_WIDTH),
		23897 => to_signed(24628, LUT_AMPL_WIDTH),
		23898 => to_signed(24626, LUT_AMPL_WIDTH),
		23899 => to_signed(24624, LUT_AMPL_WIDTH),
		23900 => to_signed(24622, LUT_AMPL_WIDTH),
		23901 => to_signed(24620, LUT_AMPL_WIDTH),
		23902 => to_signed(24618, LUT_AMPL_WIDTH),
		23903 => to_signed(24616, LUT_AMPL_WIDTH),
		23904 => to_signed(24613, LUT_AMPL_WIDTH),
		23905 => to_signed(24611, LUT_AMPL_WIDTH),
		23906 => to_signed(24609, LUT_AMPL_WIDTH),
		23907 => to_signed(24607, LUT_AMPL_WIDTH),
		23908 => to_signed(24605, LUT_AMPL_WIDTH),
		23909 => to_signed(24603, LUT_AMPL_WIDTH),
		23910 => to_signed(24601, LUT_AMPL_WIDTH),
		23911 => to_signed(24599, LUT_AMPL_WIDTH),
		23912 => to_signed(24597, LUT_AMPL_WIDTH),
		23913 => to_signed(24595, LUT_AMPL_WIDTH),
		23914 => to_signed(24593, LUT_AMPL_WIDTH),
		23915 => to_signed(24591, LUT_AMPL_WIDTH),
		23916 => to_signed(24589, LUT_AMPL_WIDTH),
		23917 => to_signed(24586, LUT_AMPL_WIDTH),
		23918 => to_signed(24584, LUT_AMPL_WIDTH),
		23919 => to_signed(24582, LUT_AMPL_WIDTH),
		23920 => to_signed(24580, LUT_AMPL_WIDTH),
		23921 => to_signed(24578, LUT_AMPL_WIDTH),
		23922 => to_signed(24576, LUT_AMPL_WIDTH),
		23923 => to_signed(24574, LUT_AMPL_WIDTH),
		23924 => to_signed(24572, LUT_AMPL_WIDTH),
		23925 => to_signed(24570, LUT_AMPL_WIDTH),
		23926 => to_signed(24568, LUT_AMPL_WIDTH),
		23927 => to_signed(24566, LUT_AMPL_WIDTH),
		23928 => to_signed(24564, LUT_AMPL_WIDTH),
		23929 => to_signed(24562, LUT_AMPL_WIDTH),
		23930 => to_signed(24559, LUT_AMPL_WIDTH),
		23931 => to_signed(24557, LUT_AMPL_WIDTH),
		23932 => to_signed(24555, LUT_AMPL_WIDTH),
		23933 => to_signed(24553, LUT_AMPL_WIDTH),
		23934 => to_signed(24551, LUT_AMPL_WIDTH),
		23935 => to_signed(24549, LUT_AMPL_WIDTH),
		23936 => to_signed(24547, LUT_AMPL_WIDTH),
		23937 => to_signed(24545, LUT_AMPL_WIDTH),
		23938 => to_signed(24543, LUT_AMPL_WIDTH),
		23939 => to_signed(24541, LUT_AMPL_WIDTH),
		23940 => to_signed(24539, LUT_AMPL_WIDTH),
		23941 => to_signed(24537, LUT_AMPL_WIDTH),
		23942 => to_signed(24534, LUT_AMPL_WIDTH),
		23943 => to_signed(24532, LUT_AMPL_WIDTH),
		23944 => to_signed(24530, LUT_AMPL_WIDTH),
		23945 => to_signed(24528, LUT_AMPL_WIDTH),
		23946 => to_signed(24526, LUT_AMPL_WIDTH),
		23947 => to_signed(24524, LUT_AMPL_WIDTH),
		23948 => to_signed(24522, LUT_AMPL_WIDTH),
		23949 => to_signed(24520, LUT_AMPL_WIDTH),
		23950 => to_signed(24518, LUT_AMPL_WIDTH),
		23951 => to_signed(24516, LUT_AMPL_WIDTH),
		23952 => to_signed(24514, LUT_AMPL_WIDTH),
		23953 => to_signed(24512, LUT_AMPL_WIDTH),
		23954 => to_signed(24509, LUT_AMPL_WIDTH),
		23955 => to_signed(24507, LUT_AMPL_WIDTH),
		23956 => to_signed(24505, LUT_AMPL_WIDTH),
		23957 => to_signed(24503, LUT_AMPL_WIDTH),
		23958 => to_signed(24501, LUT_AMPL_WIDTH),
		23959 => to_signed(24499, LUT_AMPL_WIDTH),
		23960 => to_signed(24497, LUT_AMPL_WIDTH),
		23961 => to_signed(24495, LUT_AMPL_WIDTH),
		23962 => to_signed(24493, LUT_AMPL_WIDTH),
		23963 => to_signed(24491, LUT_AMPL_WIDTH),
		23964 => to_signed(24489, LUT_AMPL_WIDTH),
		23965 => to_signed(24487, LUT_AMPL_WIDTH),
		23966 => to_signed(24484, LUT_AMPL_WIDTH),
		23967 => to_signed(24482, LUT_AMPL_WIDTH),
		23968 => to_signed(24480, LUT_AMPL_WIDTH),
		23969 => to_signed(24478, LUT_AMPL_WIDTH),
		23970 => to_signed(24476, LUT_AMPL_WIDTH),
		23971 => to_signed(24474, LUT_AMPL_WIDTH),
		23972 => to_signed(24472, LUT_AMPL_WIDTH),
		23973 => to_signed(24470, LUT_AMPL_WIDTH),
		23974 => to_signed(24468, LUT_AMPL_WIDTH),
		23975 => to_signed(24466, LUT_AMPL_WIDTH),
		23976 => to_signed(24464, LUT_AMPL_WIDTH),
		23977 => to_signed(24461, LUT_AMPL_WIDTH),
		23978 => to_signed(24459, LUT_AMPL_WIDTH),
		23979 => to_signed(24457, LUT_AMPL_WIDTH),
		23980 => to_signed(24455, LUT_AMPL_WIDTH),
		23981 => to_signed(24453, LUT_AMPL_WIDTH),
		23982 => to_signed(24451, LUT_AMPL_WIDTH),
		23983 => to_signed(24449, LUT_AMPL_WIDTH),
		23984 => to_signed(24447, LUT_AMPL_WIDTH),
		23985 => to_signed(24445, LUT_AMPL_WIDTH),
		23986 => to_signed(24443, LUT_AMPL_WIDTH),
		23987 => to_signed(24441, LUT_AMPL_WIDTH),
		23988 => to_signed(24438, LUT_AMPL_WIDTH),
		23989 => to_signed(24436, LUT_AMPL_WIDTH),
		23990 => to_signed(24434, LUT_AMPL_WIDTH),
		23991 => to_signed(24432, LUT_AMPL_WIDTH),
		23992 => to_signed(24430, LUT_AMPL_WIDTH),
		23993 => to_signed(24428, LUT_AMPL_WIDTH),
		23994 => to_signed(24426, LUT_AMPL_WIDTH),
		23995 => to_signed(24424, LUT_AMPL_WIDTH),
		23996 => to_signed(24422, LUT_AMPL_WIDTH),
		23997 => to_signed(24420, LUT_AMPL_WIDTH),
		23998 => to_signed(24417, LUT_AMPL_WIDTH),
		23999 => to_signed(24415, LUT_AMPL_WIDTH),
		24000 => to_signed(24413, LUT_AMPL_WIDTH),
		24001 => to_signed(24411, LUT_AMPL_WIDTH),
		24002 => to_signed(24409, LUT_AMPL_WIDTH),
		24003 => to_signed(24407, LUT_AMPL_WIDTH),
		24004 => to_signed(24405, LUT_AMPL_WIDTH),
		24005 => to_signed(24403, LUT_AMPL_WIDTH),
		24006 => to_signed(24401, LUT_AMPL_WIDTH),
		24007 => to_signed(24399, LUT_AMPL_WIDTH),
		24008 => to_signed(24397, LUT_AMPL_WIDTH),
		24009 => to_signed(24394, LUT_AMPL_WIDTH),
		24010 => to_signed(24392, LUT_AMPL_WIDTH),
		24011 => to_signed(24390, LUT_AMPL_WIDTH),
		24012 => to_signed(24388, LUT_AMPL_WIDTH),
		24013 => to_signed(24386, LUT_AMPL_WIDTH),
		24014 => to_signed(24384, LUT_AMPL_WIDTH),
		24015 => to_signed(24382, LUT_AMPL_WIDTH),
		24016 => to_signed(24380, LUT_AMPL_WIDTH),
		24017 => to_signed(24378, LUT_AMPL_WIDTH),
		24018 => to_signed(24376, LUT_AMPL_WIDTH),
		24019 => to_signed(24373, LUT_AMPL_WIDTH),
		24020 => to_signed(24371, LUT_AMPL_WIDTH),
		24021 => to_signed(24369, LUT_AMPL_WIDTH),
		24022 => to_signed(24367, LUT_AMPL_WIDTH),
		24023 => to_signed(24365, LUT_AMPL_WIDTH),
		24024 => to_signed(24363, LUT_AMPL_WIDTH),
		24025 => to_signed(24361, LUT_AMPL_WIDTH),
		24026 => to_signed(24359, LUT_AMPL_WIDTH),
		24027 => to_signed(24357, LUT_AMPL_WIDTH),
		24028 => to_signed(24355, LUT_AMPL_WIDTH),
		24029 => to_signed(24352, LUT_AMPL_WIDTH),
		24030 => to_signed(24350, LUT_AMPL_WIDTH),
		24031 => to_signed(24348, LUT_AMPL_WIDTH),
		24032 => to_signed(24346, LUT_AMPL_WIDTH),
		24033 => to_signed(24344, LUT_AMPL_WIDTH),
		24034 => to_signed(24342, LUT_AMPL_WIDTH),
		24035 => to_signed(24340, LUT_AMPL_WIDTH),
		24036 => to_signed(24338, LUT_AMPL_WIDTH),
		24037 => to_signed(24336, LUT_AMPL_WIDTH),
		24038 => to_signed(24334, LUT_AMPL_WIDTH),
		24039 => to_signed(24331, LUT_AMPL_WIDTH),
		24040 => to_signed(24329, LUT_AMPL_WIDTH),
		24041 => to_signed(24327, LUT_AMPL_WIDTH),
		24042 => to_signed(24325, LUT_AMPL_WIDTH),
		24043 => to_signed(24323, LUT_AMPL_WIDTH),
		24044 => to_signed(24321, LUT_AMPL_WIDTH),
		24045 => to_signed(24319, LUT_AMPL_WIDTH),
		24046 => to_signed(24317, LUT_AMPL_WIDTH),
		24047 => to_signed(24315, LUT_AMPL_WIDTH),
		24048 => to_signed(24312, LUT_AMPL_WIDTH),
		24049 => to_signed(24310, LUT_AMPL_WIDTH),
		24050 => to_signed(24308, LUT_AMPL_WIDTH),
		24051 => to_signed(24306, LUT_AMPL_WIDTH),
		24052 => to_signed(24304, LUT_AMPL_WIDTH),
		24053 => to_signed(24302, LUT_AMPL_WIDTH),
		24054 => to_signed(24300, LUT_AMPL_WIDTH),
		24055 => to_signed(24298, LUT_AMPL_WIDTH),
		24056 => to_signed(24296, LUT_AMPL_WIDTH),
		24057 => to_signed(24294, LUT_AMPL_WIDTH),
		24058 => to_signed(24291, LUT_AMPL_WIDTH),
		24059 => to_signed(24289, LUT_AMPL_WIDTH),
		24060 => to_signed(24287, LUT_AMPL_WIDTH),
		24061 => to_signed(24285, LUT_AMPL_WIDTH),
		24062 => to_signed(24283, LUT_AMPL_WIDTH),
		24063 => to_signed(24281, LUT_AMPL_WIDTH),
		24064 => to_signed(24279, LUT_AMPL_WIDTH),
		24065 => to_signed(24277, LUT_AMPL_WIDTH),
		24066 => to_signed(24275, LUT_AMPL_WIDTH),
		24067 => to_signed(24272, LUT_AMPL_WIDTH),
		24068 => to_signed(24270, LUT_AMPL_WIDTH),
		24069 => to_signed(24268, LUT_AMPL_WIDTH),
		24070 => to_signed(24266, LUT_AMPL_WIDTH),
		24071 => to_signed(24264, LUT_AMPL_WIDTH),
		24072 => to_signed(24262, LUT_AMPL_WIDTH),
		24073 => to_signed(24260, LUT_AMPL_WIDTH),
		24074 => to_signed(24258, LUT_AMPL_WIDTH),
		24075 => to_signed(24256, LUT_AMPL_WIDTH),
		24076 => to_signed(24253, LUT_AMPL_WIDTH),
		24077 => to_signed(24251, LUT_AMPL_WIDTH),
		24078 => to_signed(24249, LUT_AMPL_WIDTH),
		24079 => to_signed(24247, LUT_AMPL_WIDTH),
		24080 => to_signed(24245, LUT_AMPL_WIDTH),
		24081 => to_signed(24243, LUT_AMPL_WIDTH),
		24082 => to_signed(24241, LUT_AMPL_WIDTH),
		24083 => to_signed(24239, LUT_AMPL_WIDTH),
		24084 => to_signed(24237, LUT_AMPL_WIDTH),
		24085 => to_signed(24234, LUT_AMPL_WIDTH),
		24086 => to_signed(24232, LUT_AMPL_WIDTH),
		24087 => to_signed(24230, LUT_AMPL_WIDTH),
		24088 => to_signed(24228, LUT_AMPL_WIDTH),
		24089 => to_signed(24226, LUT_AMPL_WIDTH),
		24090 => to_signed(24224, LUT_AMPL_WIDTH),
		24091 => to_signed(24222, LUT_AMPL_WIDTH),
		24092 => to_signed(24220, LUT_AMPL_WIDTH),
		24093 => to_signed(24217, LUT_AMPL_WIDTH),
		24094 => to_signed(24215, LUT_AMPL_WIDTH),
		24095 => to_signed(24213, LUT_AMPL_WIDTH),
		24096 => to_signed(24211, LUT_AMPL_WIDTH),
		24097 => to_signed(24209, LUT_AMPL_WIDTH),
		24098 => to_signed(24207, LUT_AMPL_WIDTH),
		24099 => to_signed(24205, LUT_AMPL_WIDTH),
		24100 => to_signed(24203, LUT_AMPL_WIDTH),
		24101 => to_signed(24201, LUT_AMPL_WIDTH),
		24102 => to_signed(24198, LUT_AMPL_WIDTH),
		24103 => to_signed(24196, LUT_AMPL_WIDTH),
		24104 => to_signed(24194, LUT_AMPL_WIDTH),
		24105 => to_signed(24192, LUT_AMPL_WIDTH),
		24106 => to_signed(24190, LUT_AMPL_WIDTH),
		24107 => to_signed(24188, LUT_AMPL_WIDTH),
		24108 => to_signed(24186, LUT_AMPL_WIDTH),
		24109 => to_signed(24184, LUT_AMPL_WIDTH),
		24110 => to_signed(24181, LUT_AMPL_WIDTH),
		24111 => to_signed(24179, LUT_AMPL_WIDTH),
		24112 => to_signed(24177, LUT_AMPL_WIDTH),
		24113 => to_signed(24175, LUT_AMPL_WIDTH),
		24114 => to_signed(24173, LUT_AMPL_WIDTH),
		24115 => to_signed(24171, LUT_AMPL_WIDTH),
		24116 => to_signed(24169, LUT_AMPL_WIDTH),
		24117 => to_signed(24167, LUT_AMPL_WIDTH),
		24118 => to_signed(24164, LUT_AMPL_WIDTH),
		24119 => to_signed(24162, LUT_AMPL_WIDTH),
		24120 => to_signed(24160, LUT_AMPL_WIDTH),
		24121 => to_signed(24158, LUT_AMPL_WIDTH),
		24122 => to_signed(24156, LUT_AMPL_WIDTH),
		24123 => to_signed(24154, LUT_AMPL_WIDTH),
		24124 => to_signed(24152, LUT_AMPL_WIDTH),
		24125 => to_signed(24150, LUT_AMPL_WIDTH),
		24126 => to_signed(24148, LUT_AMPL_WIDTH),
		24127 => to_signed(24145, LUT_AMPL_WIDTH),
		24128 => to_signed(24143, LUT_AMPL_WIDTH),
		24129 => to_signed(24141, LUT_AMPL_WIDTH),
		24130 => to_signed(24139, LUT_AMPL_WIDTH),
		24131 => to_signed(24137, LUT_AMPL_WIDTH),
		24132 => to_signed(24135, LUT_AMPL_WIDTH),
		24133 => to_signed(24133, LUT_AMPL_WIDTH),
		24134 => to_signed(24131, LUT_AMPL_WIDTH),
		24135 => to_signed(24128, LUT_AMPL_WIDTH),
		24136 => to_signed(24126, LUT_AMPL_WIDTH),
		24137 => to_signed(24124, LUT_AMPL_WIDTH),
		24138 => to_signed(24122, LUT_AMPL_WIDTH),
		24139 => to_signed(24120, LUT_AMPL_WIDTH),
		24140 => to_signed(24118, LUT_AMPL_WIDTH),
		24141 => to_signed(24116, LUT_AMPL_WIDTH),
		24142 => to_signed(24114, LUT_AMPL_WIDTH),
		24143 => to_signed(24111, LUT_AMPL_WIDTH),
		24144 => to_signed(24109, LUT_AMPL_WIDTH),
		24145 => to_signed(24107, LUT_AMPL_WIDTH),
		24146 => to_signed(24105, LUT_AMPL_WIDTH),
		24147 => to_signed(24103, LUT_AMPL_WIDTH),
		24148 => to_signed(24101, LUT_AMPL_WIDTH),
		24149 => to_signed(24099, LUT_AMPL_WIDTH),
		24150 => to_signed(24096, LUT_AMPL_WIDTH),
		24151 => to_signed(24094, LUT_AMPL_WIDTH),
		24152 => to_signed(24092, LUT_AMPL_WIDTH),
		24153 => to_signed(24090, LUT_AMPL_WIDTH),
		24154 => to_signed(24088, LUT_AMPL_WIDTH),
		24155 => to_signed(24086, LUT_AMPL_WIDTH),
		24156 => to_signed(24084, LUT_AMPL_WIDTH),
		24157 => to_signed(24082, LUT_AMPL_WIDTH),
		24158 => to_signed(24079, LUT_AMPL_WIDTH),
		24159 => to_signed(24077, LUT_AMPL_WIDTH),
		24160 => to_signed(24075, LUT_AMPL_WIDTH),
		24161 => to_signed(24073, LUT_AMPL_WIDTH),
		24162 => to_signed(24071, LUT_AMPL_WIDTH),
		24163 => to_signed(24069, LUT_AMPL_WIDTH),
		24164 => to_signed(24067, LUT_AMPL_WIDTH),
		24165 => to_signed(24065, LUT_AMPL_WIDTH),
		24166 => to_signed(24062, LUT_AMPL_WIDTH),
		24167 => to_signed(24060, LUT_AMPL_WIDTH),
		24168 => to_signed(24058, LUT_AMPL_WIDTH),
		24169 => to_signed(24056, LUT_AMPL_WIDTH),
		24170 => to_signed(24054, LUT_AMPL_WIDTH),
		24171 => to_signed(24052, LUT_AMPL_WIDTH),
		24172 => to_signed(24050, LUT_AMPL_WIDTH),
		24173 => to_signed(24047, LUT_AMPL_WIDTH),
		24174 => to_signed(24045, LUT_AMPL_WIDTH),
		24175 => to_signed(24043, LUT_AMPL_WIDTH),
		24176 => to_signed(24041, LUT_AMPL_WIDTH),
		24177 => to_signed(24039, LUT_AMPL_WIDTH),
		24178 => to_signed(24037, LUT_AMPL_WIDTH),
		24179 => to_signed(24035, LUT_AMPL_WIDTH),
		24180 => to_signed(24033, LUT_AMPL_WIDTH),
		24181 => to_signed(24030, LUT_AMPL_WIDTH),
		24182 => to_signed(24028, LUT_AMPL_WIDTH),
		24183 => to_signed(24026, LUT_AMPL_WIDTH),
		24184 => to_signed(24024, LUT_AMPL_WIDTH),
		24185 => to_signed(24022, LUT_AMPL_WIDTH),
		24186 => to_signed(24020, LUT_AMPL_WIDTH),
		24187 => to_signed(24018, LUT_AMPL_WIDTH),
		24188 => to_signed(24015, LUT_AMPL_WIDTH),
		24189 => to_signed(24013, LUT_AMPL_WIDTH),
		24190 => to_signed(24011, LUT_AMPL_WIDTH),
		24191 => to_signed(24009, LUT_AMPL_WIDTH),
		24192 => to_signed(24007, LUT_AMPL_WIDTH),
		24193 => to_signed(24005, LUT_AMPL_WIDTH),
		24194 => to_signed(24003, LUT_AMPL_WIDTH),
		24195 => to_signed(24000, LUT_AMPL_WIDTH),
		24196 => to_signed(23998, LUT_AMPL_WIDTH),
		24197 => to_signed(23996, LUT_AMPL_WIDTH),
		24198 => to_signed(23994, LUT_AMPL_WIDTH),
		24199 => to_signed(23992, LUT_AMPL_WIDTH),
		24200 => to_signed(23990, LUT_AMPL_WIDTH),
		24201 => to_signed(23988, LUT_AMPL_WIDTH),
		24202 => to_signed(23985, LUT_AMPL_WIDTH),
		24203 => to_signed(23983, LUT_AMPL_WIDTH),
		24204 => to_signed(23981, LUT_AMPL_WIDTH),
		24205 => to_signed(23979, LUT_AMPL_WIDTH),
		24206 => to_signed(23977, LUT_AMPL_WIDTH),
		24207 => to_signed(23975, LUT_AMPL_WIDTH),
		24208 => to_signed(23973, LUT_AMPL_WIDTH),
		24209 => to_signed(23971, LUT_AMPL_WIDTH),
		24210 => to_signed(23968, LUT_AMPL_WIDTH),
		24211 => to_signed(23966, LUT_AMPL_WIDTH),
		24212 => to_signed(23964, LUT_AMPL_WIDTH),
		24213 => to_signed(23962, LUT_AMPL_WIDTH),
		24214 => to_signed(23960, LUT_AMPL_WIDTH),
		24215 => to_signed(23958, LUT_AMPL_WIDTH),
		24216 => to_signed(23956, LUT_AMPL_WIDTH),
		24217 => to_signed(23953, LUT_AMPL_WIDTH),
		24218 => to_signed(23951, LUT_AMPL_WIDTH),
		24219 => to_signed(23949, LUT_AMPL_WIDTH),
		24220 => to_signed(23947, LUT_AMPL_WIDTH),
		24221 => to_signed(23945, LUT_AMPL_WIDTH),
		24222 => to_signed(23943, LUT_AMPL_WIDTH),
		24223 => to_signed(23940, LUT_AMPL_WIDTH),
		24224 => to_signed(23938, LUT_AMPL_WIDTH),
		24225 => to_signed(23936, LUT_AMPL_WIDTH),
		24226 => to_signed(23934, LUT_AMPL_WIDTH),
		24227 => to_signed(23932, LUT_AMPL_WIDTH),
		24228 => to_signed(23930, LUT_AMPL_WIDTH),
		24229 => to_signed(23928, LUT_AMPL_WIDTH),
		24230 => to_signed(23925, LUT_AMPL_WIDTH),
		24231 => to_signed(23923, LUT_AMPL_WIDTH),
		24232 => to_signed(23921, LUT_AMPL_WIDTH),
		24233 => to_signed(23919, LUT_AMPL_WIDTH),
		24234 => to_signed(23917, LUT_AMPL_WIDTH),
		24235 => to_signed(23915, LUT_AMPL_WIDTH),
		24236 => to_signed(23913, LUT_AMPL_WIDTH),
		24237 => to_signed(23910, LUT_AMPL_WIDTH),
		24238 => to_signed(23908, LUT_AMPL_WIDTH),
		24239 => to_signed(23906, LUT_AMPL_WIDTH),
		24240 => to_signed(23904, LUT_AMPL_WIDTH),
		24241 => to_signed(23902, LUT_AMPL_WIDTH),
		24242 => to_signed(23900, LUT_AMPL_WIDTH),
		24243 => to_signed(23898, LUT_AMPL_WIDTH),
		24244 => to_signed(23895, LUT_AMPL_WIDTH),
		24245 => to_signed(23893, LUT_AMPL_WIDTH),
		24246 => to_signed(23891, LUT_AMPL_WIDTH),
		24247 => to_signed(23889, LUT_AMPL_WIDTH),
		24248 => to_signed(23887, LUT_AMPL_WIDTH),
		24249 => to_signed(23885, LUT_AMPL_WIDTH),
		24250 => to_signed(23883, LUT_AMPL_WIDTH),
		24251 => to_signed(23880, LUT_AMPL_WIDTH),
		24252 => to_signed(23878, LUT_AMPL_WIDTH),
		24253 => to_signed(23876, LUT_AMPL_WIDTH),
		24254 => to_signed(23874, LUT_AMPL_WIDTH),
		24255 => to_signed(23872, LUT_AMPL_WIDTH),
		24256 => to_signed(23870, LUT_AMPL_WIDTH),
		24257 => to_signed(23867, LUT_AMPL_WIDTH),
		24258 => to_signed(23865, LUT_AMPL_WIDTH),
		24259 => to_signed(23863, LUT_AMPL_WIDTH),
		24260 => to_signed(23861, LUT_AMPL_WIDTH),
		24261 => to_signed(23859, LUT_AMPL_WIDTH),
		24262 => to_signed(23857, LUT_AMPL_WIDTH),
		24263 => to_signed(23855, LUT_AMPL_WIDTH),
		24264 => to_signed(23852, LUT_AMPL_WIDTH),
		24265 => to_signed(23850, LUT_AMPL_WIDTH),
		24266 => to_signed(23848, LUT_AMPL_WIDTH),
		24267 => to_signed(23846, LUT_AMPL_WIDTH),
		24268 => to_signed(23844, LUT_AMPL_WIDTH),
		24269 => to_signed(23842, LUT_AMPL_WIDTH),
		24270 => to_signed(23839, LUT_AMPL_WIDTH),
		24271 => to_signed(23837, LUT_AMPL_WIDTH),
		24272 => to_signed(23835, LUT_AMPL_WIDTH),
		24273 => to_signed(23833, LUT_AMPL_WIDTH),
		24274 => to_signed(23831, LUT_AMPL_WIDTH),
		24275 => to_signed(23829, LUT_AMPL_WIDTH),
		24276 => to_signed(23827, LUT_AMPL_WIDTH),
		24277 => to_signed(23824, LUT_AMPL_WIDTH),
		24278 => to_signed(23822, LUT_AMPL_WIDTH),
		24279 => to_signed(23820, LUT_AMPL_WIDTH),
		24280 => to_signed(23818, LUT_AMPL_WIDTH),
		24281 => to_signed(23816, LUT_AMPL_WIDTH),
		24282 => to_signed(23814, LUT_AMPL_WIDTH),
		24283 => to_signed(23811, LUT_AMPL_WIDTH),
		24284 => to_signed(23809, LUT_AMPL_WIDTH),
		24285 => to_signed(23807, LUT_AMPL_WIDTH),
		24286 => to_signed(23805, LUT_AMPL_WIDTH),
		24287 => to_signed(23803, LUT_AMPL_WIDTH),
		24288 => to_signed(23801, LUT_AMPL_WIDTH),
		24289 => to_signed(23798, LUT_AMPL_WIDTH),
		24290 => to_signed(23796, LUT_AMPL_WIDTH),
		24291 => to_signed(23794, LUT_AMPL_WIDTH),
		24292 => to_signed(23792, LUT_AMPL_WIDTH),
		24293 => to_signed(23790, LUT_AMPL_WIDTH),
		24294 => to_signed(23788, LUT_AMPL_WIDTH),
		24295 => to_signed(23785, LUT_AMPL_WIDTH),
		24296 => to_signed(23783, LUT_AMPL_WIDTH),
		24297 => to_signed(23781, LUT_AMPL_WIDTH),
		24298 => to_signed(23779, LUT_AMPL_WIDTH),
		24299 => to_signed(23777, LUT_AMPL_WIDTH),
		24300 => to_signed(23775, LUT_AMPL_WIDTH),
		24301 => to_signed(23773, LUT_AMPL_WIDTH),
		24302 => to_signed(23770, LUT_AMPL_WIDTH),
		24303 => to_signed(23768, LUT_AMPL_WIDTH),
		24304 => to_signed(23766, LUT_AMPL_WIDTH),
		24305 => to_signed(23764, LUT_AMPL_WIDTH),
		24306 => to_signed(23762, LUT_AMPL_WIDTH),
		24307 => to_signed(23760, LUT_AMPL_WIDTH),
		24308 => to_signed(23757, LUT_AMPL_WIDTH),
		24309 => to_signed(23755, LUT_AMPL_WIDTH),
		24310 => to_signed(23753, LUT_AMPL_WIDTH),
		24311 => to_signed(23751, LUT_AMPL_WIDTH),
		24312 => to_signed(23749, LUT_AMPL_WIDTH),
		24313 => to_signed(23747, LUT_AMPL_WIDTH),
		24314 => to_signed(23744, LUT_AMPL_WIDTH),
		24315 => to_signed(23742, LUT_AMPL_WIDTH),
		24316 => to_signed(23740, LUT_AMPL_WIDTH),
		24317 => to_signed(23738, LUT_AMPL_WIDTH),
		24318 => to_signed(23736, LUT_AMPL_WIDTH),
		24319 => to_signed(23734, LUT_AMPL_WIDTH),
		24320 => to_signed(23731, LUT_AMPL_WIDTH),
		24321 => to_signed(23729, LUT_AMPL_WIDTH),
		24322 => to_signed(23727, LUT_AMPL_WIDTH),
		24323 => to_signed(23725, LUT_AMPL_WIDTH),
		24324 => to_signed(23723, LUT_AMPL_WIDTH),
		24325 => to_signed(23721, LUT_AMPL_WIDTH),
		24326 => to_signed(23718, LUT_AMPL_WIDTH),
		24327 => to_signed(23716, LUT_AMPL_WIDTH),
		24328 => to_signed(23714, LUT_AMPL_WIDTH),
		24329 => to_signed(23712, LUT_AMPL_WIDTH),
		24330 => to_signed(23710, LUT_AMPL_WIDTH),
		24331 => to_signed(23708, LUT_AMPL_WIDTH),
		24332 => to_signed(23705, LUT_AMPL_WIDTH),
		24333 => to_signed(23703, LUT_AMPL_WIDTH),
		24334 => to_signed(23701, LUT_AMPL_WIDTH),
		24335 => to_signed(23699, LUT_AMPL_WIDTH),
		24336 => to_signed(23697, LUT_AMPL_WIDTH),
		24337 => to_signed(23695, LUT_AMPL_WIDTH),
		24338 => to_signed(23692, LUT_AMPL_WIDTH),
		24339 => to_signed(23690, LUT_AMPL_WIDTH),
		24340 => to_signed(23688, LUT_AMPL_WIDTH),
		24341 => to_signed(23686, LUT_AMPL_WIDTH),
		24342 => to_signed(23684, LUT_AMPL_WIDTH),
		24343 => to_signed(23682, LUT_AMPL_WIDTH),
		24344 => to_signed(23679, LUT_AMPL_WIDTH),
		24345 => to_signed(23677, LUT_AMPL_WIDTH),
		24346 => to_signed(23675, LUT_AMPL_WIDTH),
		24347 => to_signed(23673, LUT_AMPL_WIDTH),
		24348 => to_signed(23671, LUT_AMPL_WIDTH),
		24349 => to_signed(23668, LUT_AMPL_WIDTH),
		24350 => to_signed(23666, LUT_AMPL_WIDTH),
		24351 => to_signed(23664, LUT_AMPL_WIDTH),
		24352 => to_signed(23662, LUT_AMPL_WIDTH),
		24353 => to_signed(23660, LUT_AMPL_WIDTH),
		24354 => to_signed(23658, LUT_AMPL_WIDTH),
		24355 => to_signed(23655, LUT_AMPL_WIDTH),
		24356 => to_signed(23653, LUT_AMPL_WIDTH),
		24357 => to_signed(23651, LUT_AMPL_WIDTH),
		24358 => to_signed(23649, LUT_AMPL_WIDTH),
		24359 => to_signed(23647, LUT_AMPL_WIDTH),
		24360 => to_signed(23645, LUT_AMPL_WIDTH),
		24361 => to_signed(23642, LUT_AMPL_WIDTH),
		24362 => to_signed(23640, LUT_AMPL_WIDTH),
		24363 => to_signed(23638, LUT_AMPL_WIDTH),
		24364 => to_signed(23636, LUT_AMPL_WIDTH),
		24365 => to_signed(23634, LUT_AMPL_WIDTH),
		24366 => to_signed(23632, LUT_AMPL_WIDTH),
		24367 => to_signed(23629, LUT_AMPL_WIDTH),
		24368 => to_signed(23627, LUT_AMPL_WIDTH),
		24369 => to_signed(23625, LUT_AMPL_WIDTH),
		24370 => to_signed(23623, LUT_AMPL_WIDTH),
		24371 => to_signed(23621, LUT_AMPL_WIDTH),
		24372 => to_signed(23618, LUT_AMPL_WIDTH),
		24373 => to_signed(23616, LUT_AMPL_WIDTH),
		24374 => to_signed(23614, LUT_AMPL_WIDTH),
		24375 => to_signed(23612, LUT_AMPL_WIDTH),
		24376 => to_signed(23610, LUT_AMPL_WIDTH),
		24377 => to_signed(23608, LUT_AMPL_WIDTH),
		24378 => to_signed(23605, LUT_AMPL_WIDTH),
		24379 => to_signed(23603, LUT_AMPL_WIDTH),
		24380 => to_signed(23601, LUT_AMPL_WIDTH),
		24381 => to_signed(23599, LUT_AMPL_WIDTH),
		24382 => to_signed(23597, LUT_AMPL_WIDTH),
		24383 => to_signed(23595, LUT_AMPL_WIDTH),
		24384 => to_signed(23592, LUT_AMPL_WIDTH),
		24385 => to_signed(23590, LUT_AMPL_WIDTH),
		24386 => to_signed(23588, LUT_AMPL_WIDTH),
		24387 => to_signed(23586, LUT_AMPL_WIDTH),
		24388 => to_signed(23584, LUT_AMPL_WIDTH),
		24389 => to_signed(23581, LUT_AMPL_WIDTH),
		24390 => to_signed(23579, LUT_AMPL_WIDTH),
		24391 => to_signed(23577, LUT_AMPL_WIDTH),
		24392 => to_signed(23575, LUT_AMPL_WIDTH),
		24393 => to_signed(23573, LUT_AMPL_WIDTH),
		24394 => to_signed(23571, LUT_AMPL_WIDTH),
		24395 => to_signed(23568, LUT_AMPL_WIDTH),
		24396 => to_signed(23566, LUT_AMPL_WIDTH),
		24397 => to_signed(23564, LUT_AMPL_WIDTH),
		24398 => to_signed(23562, LUT_AMPL_WIDTH),
		24399 => to_signed(23560, LUT_AMPL_WIDTH),
		24400 => to_signed(23557, LUT_AMPL_WIDTH),
		24401 => to_signed(23555, LUT_AMPL_WIDTH),
		24402 => to_signed(23553, LUT_AMPL_WIDTH),
		24403 => to_signed(23551, LUT_AMPL_WIDTH),
		24404 => to_signed(23549, LUT_AMPL_WIDTH),
		24405 => to_signed(23546, LUT_AMPL_WIDTH),
		24406 => to_signed(23544, LUT_AMPL_WIDTH),
		24407 => to_signed(23542, LUT_AMPL_WIDTH),
		24408 => to_signed(23540, LUT_AMPL_WIDTH),
		24409 => to_signed(23538, LUT_AMPL_WIDTH),
		24410 => to_signed(23536, LUT_AMPL_WIDTH),
		24411 => to_signed(23533, LUT_AMPL_WIDTH),
		24412 => to_signed(23531, LUT_AMPL_WIDTH),
		24413 => to_signed(23529, LUT_AMPL_WIDTH),
		24414 => to_signed(23527, LUT_AMPL_WIDTH),
		24415 => to_signed(23525, LUT_AMPL_WIDTH),
		24416 => to_signed(23522, LUT_AMPL_WIDTH),
		24417 => to_signed(23520, LUT_AMPL_WIDTH),
		24418 => to_signed(23518, LUT_AMPL_WIDTH),
		24419 => to_signed(23516, LUT_AMPL_WIDTH),
		24420 => to_signed(23514, LUT_AMPL_WIDTH),
		24421 => to_signed(23512, LUT_AMPL_WIDTH),
		24422 => to_signed(23509, LUT_AMPL_WIDTH),
		24423 => to_signed(23507, LUT_AMPL_WIDTH),
		24424 => to_signed(23505, LUT_AMPL_WIDTH),
		24425 => to_signed(23503, LUT_AMPL_WIDTH),
		24426 => to_signed(23501, LUT_AMPL_WIDTH),
		24427 => to_signed(23498, LUT_AMPL_WIDTH),
		24428 => to_signed(23496, LUT_AMPL_WIDTH),
		24429 => to_signed(23494, LUT_AMPL_WIDTH),
		24430 => to_signed(23492, LUT_AMPL_WIDTH),
		24431 => to_signed(23490, LUT_AMPL_WIDTH),
		24432 => to_signed(23487, LUT_AMPL_WIDTH),
		24433 => to_signed(23485, LUT_AMPL_WIDTH),
		24434 => to_signed(23483, LUT_AMPL_WIDTH),
		24435 => to_signed(23481, LUT_AMPL_WIDTH),
		24436 => to_signed(23479, LUT_AMPL_WIDTH),
		24437 => to_signed(23476, LUT_AMPL_WIDTH),
		24438 => to_signed(23474, LUT_AMPL_WIDTH),
		24439 => to_signed(23472, LUT_AMPL_WIDTH),
		24440 => to_signed(23470, LUT_AMPL_WIDTH),
		24441 => to_signed(23468, LUT_AMPL_WIDTH),
		24442 => to_signed(23466, LUT_AMPL_WIDTH),
		24443 => to_signed(23463, LUT_AMPL_WIDTH),
		24444 => to_signed(23461, LUT_AMPL_WIDTH),
		24445 => to_signed(23459, LUT_AMPL_WIDTH),
		24446 => to_signed(23457, LUT_AMPL_WIDTH),
		24447 => to_signed(23455, LUT_AMPL_WIDTH),
		24448 => to_signed(23452, LUT_AMPL_WIDTH),
		24449 => to_signed(23450, LUT_AMPL_WIDTH),
		24450 => to_signed(23448, LUT_AMPL_WIDTH),
		24451 => to_signed(23446, LUT_AMPL_WIDTH),
		24452 => to_signed(23444, LUT_AMPL_WIDTH),
		24453 => to_signed(23441, LUT_AMPL_WIDTH),
		24454 => to_signed(23439, LUT_AMPL_WIDTH),
		24455 => to_signed(23437, LUT_AMPL_WIDTH),
		24456 => to_signed(23435, LUT_AMPL_WIDTH),
		24457 => to_signed(23433, LUT_AMPL_WIDTH),
		24458 => to_signed(23430, LUT_AMPL_WIDTH),
		24459 => to_signed(23428, LUT_AMPL_WIDTH),
		24460 => to_signed(23426, LUT_AMPL_WIDTH),
		24461 => to_signed(23424, LUT_AMPL_WIDTH),
		24462 => to_signed(23422, LUT_AMPL_WIDTH),
		24463 => to_signed(23419, LUT_AMPL_WIDTH),
		24464 => to_signed(23417, LUT_AMPL_WIDTH),
		24465 => to_signed(23415, LUT_AMPL_WIDTH),
		24466 => to_signed(23413, LUT_AMPL_WIDTH),
		24467 => to_signed(23411, LUT_AMPL_WIDTH),
		24468 => to_signed(23408, LUT_AMPL_WIDTH),
		24469 => to_signed(23406, LUT_AMPL_WIDTH),
		24470 => to_signed(23404, LUT_AMPL_WIDTH),
		24471 => to_signed(23402, LUT_AMPL_WIDTH),
		24472 => to_signed(23400, LUT_AMPL_WIDTH),
		24473 => to_signed(23397, LUT_AMPL_WIDTH),
		24474 => to_signed(23395, LUT_AMPL_WIDTH),
		24475 => to_signed(23393, LUT_AMPL_WIDTH),
		24476 => to_signed(23391, LUT_AMPL_WIDTH),
		24477 => to_signed(23389, LUT_AMPL_WIDTH),
		24478 => to_signed(23386, LUT_AMPL_WIDTH),
		24479 => to_signed(23384, LUT_AMPL_WIDTH),
		24480 => to_signed(23382, LUT_AMPL_WIDTH),
		24481 => to_signed(23380, LUT_AMPL_WIDTH),
		24482 => to_signed(23378, LUT_AMPL_WIDTH),
		24483 => to_signed(23375, LUT_AMPL_WIDTH),
		24484 => to_signed(23373, LUT_AMPL_WIDTH),
		24485 => to_signed(23371, LUT_AMPL_WIDTH),
		24486 => to_signed(23369, LUT_AMPL_WIDTH),
		24487 => to_signed(23367, LUT_AMPL_WIDTH),
		24488 => to_signed(23364, LUT_AMPL_WIDTH),
		24489 => to_signed(23362, LUT_AMPL_WIDTH),
		24490 => to_signed(23360, LUT_AMPL_WIDTH),
		24491 => to_signed(23358, LUT_AMPL_WIDTH),
		24492 => to_signed(23356, LUT_AMPL_WIDTH),
		24493 => to_signed(23353, LUT_AMPL_WIDTH),
		24494 => to_signed(23351, LUT_AMPL_WIDTH),
		24495 => to_signed(23349, LUT_AMPL_WIDTH),
		24496 => to_signed(23347, LUT_AMPL_WIDTH),
		24497 => to_signed(23345, LUT_AMPL_WIDTH),
		24498 => to_signed(23342, LUT_AMPL_WIDTH),
		24499 => to_signed(23340, LUT_AMPL_WIDTH),
		24500 => to_signed(23338, LUT_AMPL_WIDTH),
		24501 => to_signed(23336, LUT_AMPL_WIDTH),
		24502 => to_signed(23334, LUT_AMPL_WIDTH),
		24503 => to_signed(23331, LUT_AMPL_WIDTH),
		24504 => to_signed(23329, LUT_AMPL_WIDTH),
		24505 => to_signed(23327, LUT_AMPL_WIDTH),
		24506 => to_signed(23325, LUT_AMPL_WIDTH),
		24507 => to_signed(23323, LUT_AMPL_WIDTH),
		24508 => to_signed(23320, LUT_AMPL_WIDTH),
		24509 => to_signed(23318, LUT_AMPL_WIDTH),
		24510 => to_signed(23316, LUT_AMPL_WIDTH),
		24511 => to_signed(23314, LUT_AMPL_WIDTH),
		24512 => to_signed(23311, LUT_AMPL_WIDTH),
		24513 => to_signed(23309, LUT_AMPL_WIDTH),
		24514 => to_signed(23307, LUT_AMPL_WIDTH),
		24515 => to_signed(23305, LUT_AMPL_WIDTH),
		24516 => to_signed(23303, LUT_AMPL_WIDTH),
		24517 => to_signed(23300, LUT_AMPL_WIDTH),
		24518 => to_signed(23298, LUT_AMPL_WIDTH),
		24519 => to_signed(23296, LUT_AMPL_WIDTH),
		24520 => to_signed(23294, LUT_AMPL_WIDTH),
		24521 => to_signed(23292, LUT_AMPL_WIDTH),
		24522 => to_signed(23289, LUT_AMPL_WIDTH),
		24523 => to_signed(23287, LUT_AMPL_WIDTH),
		24524 => to_signed(23285, LUT_AMPL_WIDTH),
		24525 => to_signed(23283, LUT_AMPL_WIDTH),
		24526 => to_signed(23281, LUT_AMPL_WIDTH),
		24527 => to_signed(23278, LUT_AMPL_WIDTH),
		24528 => to_signed(23276, LUT_AMPL_WIDTH),
		24529 => to_signed(23274, LUT_AMPL_WIDTH),
		24530 => to_signed(23272, LUT_AMPL_WIDTH),
		24531 => to_signed(23270, LUT_AMPL_WIDTH),
		24532 => to_signed(23267, LUT_AMPL_WIDTH),
		24533 => to_signed(23265, LUT_AMPL_WIDTH),
		24534 => to_signed(23263, LUT_AMPL_WIDTH),
		24535 => to_signed(23261, LUT_AMPL_WIDTH),
		24536 => to_signed(23258, LUT_AMPL_WIDTH),
		24537 => to_signed(23256, LUT_AMPL_WIDTH),
		24538 => to_signed(23254, LUT_AMPL_WIDTH),
		24539 => to_signed(23252, LUT_AMPL_WIDTH),
		24540 => to_signed(23250, LUT_AMPL_WIDTH),
		24541 => to_signed(23247, LUT_AMPL_WIDTH),
		24542 => to_signed(23245, LUT_AMPL_WIDTH),
		24543 => to_signed(23243, LUT_AMPL_WIDTH),
		24544 => to_signed(23241, LUT_AMPL_WIDTH),
		24545 => to_signed(23239, LUT_AMPL_WIDTH),
		24546 => to_signed(23236, LUT_AMPL_WIDTH),
		24547 => to_signed(23234, LUT_AMPL_WIDTH),
		24548 => to_signed(23232, LUT_AMPL_WIDTH),
		24549 => to_signed(23230, LUT_AMPL_WIDTH),
		24550 => to_signed(23227, LUT_AMPL_WIDTH),
		24551 => to_signed(23225, LUT_AMPL_WIDTH),
		24552 => to_signed(23223, LUT_AMPL_WIDTH),
		24553 => to_signed(23221, LUT_AMPL_WIDTH),
		24554 => to_signed(23219, LUT_AMPL_WIDTH),
		24555 => to_signed(23216, LUT_AMPL_WIDTH),
		24556 => to_signed(23214, LUT_AMPL_WIDTH),
		24557 => to_signed(23212, LUT_AMPL_WIDTH),
		24558 => to_signed(23210, LUT_AMPL_WIDTH),
		24559 => to_signed(23208, LUT_AMPL_WIDTH),
		24560 => to_signed(23205, LUT_AMPL_WIDTH),
		24561 => to_signed(23203, LUT_AMPL_WIDTH),
		24562 => to_signed(23201, LUT_AMPL_WIDTH),
		24563 => to_signed(23199, LUT_AMPL_WIDTH),
		24564 => to_signed(23196, LUT_AMPL_WIDTH),
		24565 => to_signed(23194, LUT_AMPL_WIDTH),
		24566 => to_signed(23192, LUT_AMPL_WIDTH),
		24567 => to_signed(23190, LUT_AMPL_WIDTH),
		24568 => to_signed(23188, LUT_AMPL_WIDTH),
		24569 => to_signed(23185, LUT_AMPL_WIDTH),
		24570 => to_signed(23183, LUT_AMPL_WIDTH),
		24571 => to_signed(23181, LUT_AMPL_WIDTH),
		24572 => to_signed(23179, LUT_AMPL_WIDTH),
		24573 => to_signed(23176, LUT_AMPL_WIDTH),
		24574 => to_signed(23174, LUT_AMPL_WIDTH),
		24575 => to_signed(23172, LUT_AMPL_WIDTH),
		24576 => to_signed(23170, LUT_AMPL_WIDTH),
		24577 => to_signed(23168, LUT_AMPL_WIDTH),
		24578 => to_signed(23165, LUT_AMPL_WIDTH),
		24579 => to_signed(23163, LUT_AMPL_WIDTH),
		24580 => to_signed(23161, LUT_AMPL_WIDTH),
		24581 => to_signed(23159, LUT_AMPL_WIDTH),
		24582 => to_signed(23156, LUT_AMPL_WIDTH),
		24583 => to_signed(23154, LUT_AMPL_WIDTH),
		24584 => to_signed(23152, LUT_AMPL_WIDTH),
		24585 => to_signed(23150, LUT_AMPL_WIDTH),
		24586 => to_signed(23148, LUT_AMPL_WIDTH),
		24587 => to_signed(23145, LUT_AMPL_WIDTH),
		24588 => to_signed(23143, LUT_AMPL_WIDTH),
		24589 => to_signed(23141, LUT_AMPL_WIDTH),
		24590 => to_signed(23139, LUT_AMPL_WIDTH),
		24591 => to_signed(23136, LUT_AMPL_WIDTH),
		24592 => to_signed(23134, LUT_AMPL_WIDTH),
		24593 => to_signed(23132, LUT_AMPL_WIDTH),
		24594 => to_signed(23130, LUT_AMPL_WIDTH),
		24595 => to_signed(23128, LUT_AMPL_WIDTH),
		24596 => to_signed(23125, LUT_AMPL_WIDTH),
		24597 => to_signed(23123, LUT_AMPL_WIDTH),
		24598 => to_signed(23121, LUT_AMPL_WIDTH),
		24599 => to_signed(23119, LUT_AMPL_WIDTH),
		24600 => to_signed(23116, LUT_AMPL_WIDTH),
		24601 => to_signed(23114, LUT_AMPL_WIDTH),
		24602 => to_signed(23112, LUT_AMPL_WIDTH),
		24603 => to_signed(23110, LUT_AMPL_WIDTH),
		24604 => to_signed(23107, LUT_AMPL_WIDTH),
		24605 => to_signed(23105, LUT_AMPL_WIDTH),
		24606 => to_signed(23103, LUT_AMPL_WIDTH),
		24607 => to_signed(23101, LUT_AMPL_WIDTH),
		24608 => to_signed(23099, LUT_AMPL_WIDTH),
		24609 => to_signed(23096, LUT_AMPL_WIDTH),
		24610 => to_signed(23094, LUT_AMPL_WIDTH),
		24611 => to_signed(23092, LUT_AMPL_WIDTH),
		24612 => to_signed(23090, LUT_AMPL_WIDTH),
		24613 => to_signed(23087, LUT_AMPL_WIDTH),
		24614 => to_signed(23085, LUT_AMPL_WIDTH),
		24615 => to_signed(23083, LUT_AMPL_WIDTH),
		24616 => to_signed(23081, LUT_AMPL_WIDTH),
		24617 => to_signed(23079, LUT_AMPL_WIDTH),
		24618 => to_signed(23076, LUT_AMPL_WIDTH),
		24619 => to_signed(23074, LUT_AMPL_WIDTH),
		24620 => to_signed(23072, LUT_AMPL_WIDTH),
		24621 => to_signed(23070, LUT_AMPL_WIDTH),
		24622 => to_signed(23067, LUT_AMPL_WIDTH),
		24623 => to_signed(23065, LUT_AMPL_WIDTH),
		24624 => to_signed(23063, LUT_AMPL_WIDTH),
		24625 => to_signed(23061, LUT_AMPL_WIDTH),
		24626 => to_signed(23058, LUT_AMPL_WIDTH),
		24627 => to_signed(23056, LUT_AMPL_WIDTH),
		24628 => to_signed(23054, LUT_AMPL_WIDTH),
		24629 => to_signed(23052, LUT_AMPL_WIDTH),
		24630 => to_signed(23050, LUT_AMPL_WIDTH),
		24631 => to_signed(23047, LUT_AMPL_WIDTH),
		24632 => to_signed(23045, LUT_AMPL_WIDTH),
		24633 => to_signed(23043, LUT_AMPL_WIDTH),
		24634 => to_signed(23041, LUT_AMPL_WIDTH),
		24635 => to_signed(23038, LUT_AMPL_WIDTH),
		24636 => to_signed(23036, LUT_AMPL_WIDTH),
		24637 => to_signed(23034, LUT_AMPL_WIDTH),
		24638 => to_signed(23032, LUT_AMPL_WIDTH),
		24639 => to_signed(23029, LUT_AMPL_WIDTH),
		24640 => to_signed(23027, LUT_AMPL_WIDTH),
		24641 => to_signed(23025, LUT_AMPL_WIDTH),
		24642 => to_signed(23023, LUT_AMPL_WIDTH),
		24643 => to_signed(23020, LUT_AMPL_WIDTH),
		24644 => to_signed(23018, LUT_AMPL_WIDTH),
		24645 => to_signed(23016, LUT_AMPL_WIDTH),
		24646 => to_signed(23014, LUT_AMPL_WIDTH),
		24647 => to_signed(23012, LUT_AMPL_WIDTH),
		24648 => to_signed(23009, LUT_AMPL_WIDTH),
		24649 => to_signed(23007, LUT_AMPL_WIDTH),
		24650 => to_signed(23005, LUT_AMPL_WIDTH),
		24651 => to_signed(23003, LUT_AMPL_WIDTH),
		24652 => to_signed(23000, LUT_AMPL_WIDTH),
		24653 => to_signed(22998, LUT_AMPL_WIDTH),
		24654 => to_signed(22996, LUT_AMPL_WIDTH),
		24655 => to_signed(22994, LUT_AMPL_WIDTH),
		24656 => to_signed(22991, LUT_AMPL_WIDTH),
		24657 => to_signed(22989, LUT_AMPL_WIDTH),
		24658 => to_signed(22987, LUT_AMPL_WIDTH),
		24659 => to_signed(22985, LUT_AMPL_WIDTH),
		24660 => to_signed(22982, LUT_AMPL_WIDTH),
		24661 => to_signed(22980, LUT_AMPL_WIDTH),
		24662 => to_signed(22978, LUT_AMPL_WIDTH),
		24663 => to_signed(22976, LUT_AMPL_WIDTH),
		24664 => to_signed(22973, LUT_AMPL_WIDTH),
		24665 => to_signed(22971, LUT_AMPL_WIDTH),
		24666 => to_signed(22969, LUT_AMPL_WIDTH),
		24667 => to_signed(22967, LUT_AMPL_WIDTH),
		24668 => to_signed(22965, LUT_AMPL_WIDTH),
		24669 => to_signed(22962, LUT_AMPL_WIDTH),
		24670 => to_signed(22960, LUT_AMPL_WIDTH),
		24671 => to_signed(22958, LUT_AMPL_WIDTH),
		24672 => to_signed(22956, LUT_AMPL_WIDTH),
		24673 => to_signed(22953, LUT_AMPL_WIDTH),
		24674 => to_signed(22951, LUT_AMPL_WIDTH),
		24675 => to_signed(22949, LUT_AMPL_WIDTH),
		24676 => to_signed(22947, LUT_AMPL_WIDTH),
		24677 => to_signed(22944, LUT_AMPL_WIDTH),
		24678 => to_signed(22942, LUT_AMPL_WIDTH),
		24679 => to_signed(22940, LUT_AMPL_WIDTH),
		24680 => to_signed(22938, LUT_AMPL_WIDTH),
		24681 => to_signed(22935, LUT_AMPL_WIDTH),
		24682 => to_signed(22933, LUT_AMPL_WIDTH),
		24683 => to_signed(22931, LUT_AMPL_WIDTH),
		24684 => to_signed(22929, LUT_AMPL_WIDTH),
		24685 => to_signed(22926, LUT_AMPL_WIDTH),
		24686 => to_signed(22924, LUT_AMPL_WIDTH),
		24687 => to_signed(22922, LUT_AMPL_WIDTH),
		24688 => to_signed(22920, LUT_AMPL_WIDTH),
		24689 => to_signed(22917, LUT_AMPL_WIDTH),
		24690 => to_signed(22915, LUT_AMPL_WIDTH),
		24691 => to_signed(22913, LUT_AMPL_WIDTH),
		24692 => to_signed(22911, LUT_AMPL_WIDTH),
		24693 => to_signed(22908, LUT_AMPL_WIDTH),
		24694 => to_signed(22906, LUT_AMPL_WIDTH),
		24695 => to_signed(22904, LUT_AMPL_WIDTH),
		24696 => to_signed(22902, LUT_AMPL_WIDTH),
		24697 => to_signed(22899, LUT_AMPL_WIDTH),
		24698 => to_signed(22897, LUT_AMPL_WIDTH),
		24699 => to_signed(22895, LUT_AMPL_WIDTH),
		24700 => to_signed(22893, LUT_AMPL_WIDTH),
		24701 => to_signed(22890, LUT_AMPL_WIDTH),
		24702 => to_signed(22888, LUT_AMPL_WIDTH),
		24703 => to_signed(22886, LUT_AMPL_WIDTH),
		24704 => to_signed(22884, LUT_AMPL_WIDTH),
		24705 => to_signed(22881, LUT_AMPL_WIDTH),
		24706 => to_signed(22879, LUT_AMPL_WIDTH),
		24707 => to_signed(22877, LUT_AMPL_WIDTH),
		24708 => to_signed(22875, LUT_AMPL_WIDTH),
		24709 => to_signed(22872, LUT_AMPL_WIDTH),
		24710 => to_signed(22870, LUT_AMPL_WIDTH),
		24711 => to_signed(22868, LUT_AMPL_WIDTH),
		24712 => to_signed(22866, LUT_AMPL_WIDTH),
		24713 => to_signed(22863, LUT_AMPL_WIDTH),
		24714 => to_signed(22861, LUT_AMPL_WIDTH),
		24715 => to_signed(22859, LUT_AMPL_WIDTH),
		24716 => to_signed(22857, LUT_AMPL_WIDTH),
		24717 => to_signed(22854, LUT_AMPL_WIDTH),
		24718 => to_signed(22852, LUT_AMPL_WIDTH),
		24719 => to_signed(22850, LUT_AMPL_WIDTH),
		24720 => to_signed(22848, LUT_AMPL_WIDTH),
		24721 => to_signed(22845, LUT_AMPL_WIDTH),
		24722 => to_signed(22843, LUT_AMPL_WIDTH),
		24723 => to_signed(22841, LUT_AMPL_WIDTH),
		24724 => to_signed(22839, LUT_AMPL_WIDTH),
		24725 => to_signed(22836, LUT_AMPL_WIDTH),
		24726 => to_signed(22834, LUT_AMPL_WIDTH),
		24727 => to_signed(22832, LUT_AMPL_WIDTH),
		24728 => to_signed(22830, LUT_AMPL_WIDTH),
		24729 => to_signed(22827, LUT_AMPL_WIDTH),
		24730 => to_signed(22825, LUT_AMPL_WIDTH),
		24731 => to_signed(22823, LUT_AMPL_WIDTH),
		24732 => to_signed(22821, LUT_AMPL_WIDTH),
		24733 => to_signed(22818, LUT_AMPL_WIDTH),
		24734 => to_signed(22816, LUT_AMPL_WIDTH),
		24735 => to_signed(22814, LUT_AMPL_WIDTH),
		24736 => to_signed(22812, LUT_AMPL_WIDTH),
		24737 => to_signed(22809, LUT_AMPL_WIDTH),
		24738 => to_signed(22807, LUT_AMPL_WIDTH),
		24739 => to_signed(22805, LUT_AMPL_WIDTH),
		24740 => to_signed(22803, LUT_AMPL_WIDTH),
		24741 => to_signed(22800, LUT_AMPL_WIDTH),
		24742 => to_signed(22798, LUT_AMPL_WIDTH),
		24743 => to_signed(22796, LUT_AMPL_WIDTH),
		24744 => to_signed(22794, LUT_AMPL_WIDTH),
		24745 => to_signed(22791, LUT_AMPL_WIDTH),
		24746 => to_signed(22789, LUT_AMPL_WIDTH),
		24747 => to_signed(22787, LUT_AMPL_WIDTH),
		24748 => to_signed(22785, LUT_AMPL_WIDTH),
		24749 => to_signed(22782, LUT_AMPL_WIDTH),
		24750 => to_signed(22780, LUT_AMPL_WIDTH),
		24751 => to_signed(22778, LUT_AMPL_WIDTH),
		24752 => to_signed(22776, LUT_AMPL_WIDTH),
		24753 => to_signed(22773, LUT_AMPL_WIDTH),
		24754 => to_signed(22771, LUT_AMPL_WIDTH),
		24755 => to_signed(22769, LUT_AMPL_WIDTH),
		24756 => to_signed(22766, LUT_AMPL_WIDTH),
		24757 => to_signed(22764, LUT_AMPL_WIDTH),
		24758 => to_signed(22762, LUT_AMPL_WIDTH),
		24759 => to_signed(22760, LUT_AMPL_WIDTH),
		24760 => to_signed(22757, LUT_AMPL_WIDTH),
		24761 => to_signed(22755, LUT_AMPL_WIDTH),
		24762 => to_signed(22753, LUT_AMPL_WIDTH),
		24763 => to_signed(22751, LUT_AMPL_WIDTH),
		24764 => to_signed(22748, LUT_AMPL_WIDTH),
		24765 => to_signed(22746, LUT_AMPL_WIDTH),
		24766 => to_signed(22744, LUT_AMPL_WIDTH),
		24767 => to_signed(22742, LUT_AMPL_WIDTH),
		24768 => to_signed(22739, LUT_AMPL_WIDTH),
		24769 => to_signed(22737, LUT_AMPL_WIDTH),
		24770 => to_signed(22735, LUT_AMPL_WIDTH),
		24771 => to_signed(22733, LUT_AMPL_WIDTH),
		24772 => to_signed(22730, LUT_AMPL_WIDTH),
		24773 => to_signed(22728, LUT_AMPL_WIDTH),
		24774 => to_signed(22726, LUT_AMPL_WIDTH),
		24775 => to_signed(22724, LUT_AMPL_WIDTH),
		24776 => to_signed(22721, LUT_AMPL_WIDTH),
		24777 => to_signed(22719, LUT_AMPL_WIDTH),
		24778 => to_signed(22717, LUT_AMPL_WIDTH),
		24779 => to_signed(22714, LUT_AMPL_WIDTH),
		24780 => to_signed(22712, LUT_AMPL_WIDTH),
		24781 => to_signed(22710, LUT_AMPL_WIDTH),
		24782 => to_signed(22708, LUT_AMPL_WIDTH),
		24783 => to_signed(22705, LUT_AMPL_WIDTH),
		24784 => to_signed(22703, LUT_AMPL_WIDTH),
		24785 => to_signed(22701, LUT_AMPL_WIDTH),
		24786 => to_signed(22699, LUT_AMPL_WIDTH),
		24787 => to_signed(22696, LUT_AMPL_WIDTH),
		24788 => to_signed(22694, LUT_AMPL_WIDTH),
		24789 => to_signed(22692, LUT_AMPL_WIDTH),
		24790 => to_signed(22690, LUT_AMPL_WIDTH),
		24791 => to_signed(22687, LUT_AMPL_WIDTH),
		24792 => to_signed(22685, LUT_AMPL_WIDTH),
		24793 => to_signed(22683, LUT_AMPL_WIDTH),
		24794 => to_signed(22680, LUT_AMPL_WIDTH),
		24795 => to_signed(22678, LUT_AMPL_WIDTH),
		24796 => to_signed(22676, LUT_AMPL_WIDTH),
		24797 => to_signed(22674, LUT_AMPL_WIDTH),
		24798 => to_signed(22671, LUT_AMPL_WIDTH),
		24799 => to_signed(22669, LUT_AMPL_WIDTH),
		24800 => to_signed(22667, LUT_AMPL_WIDTH),
		24801 => to_signed(22665, LUT_AMPL_WIDTH),
		24802 => to_signed(22662, LUT_AMPL_WIDTH),
		24803 => to_signed(22660, LUT_AMPL_WIDTH),
		24804 => to_signed(22658, LUT_AMPL_WIDTH),
		24805 => to_signed(22656, LUT_AMPL_WIDTH),
		24806 => to_signed(22653, LUT_AMPL_WIDTH),
		24807 => to_signed(22651, LUT_AMPL_WIDTH),
		24808 => to_signed(22649, LUT_AMPL_WIDTH),
		24809 => to_signed(22646, LUT_AMPL_WIDTH),
		24810 => to_signed(22644, LUT_AMPL_WIDTH),
		24811 => to_signed(22642, LUT_AMPL_WIDTH),
		24812 => to_signed(22640, LUT_AMPL_WIDTH),
		24813 => to_signed(22637, LUT_AMPL_WIDTH),
		24814 => to_signed(22635, LUT_AMPL_WIDTH),
		24815 => to_signed(22633, LUT_AMPL_WIDTH),
		24816 => to_signed(22631, LUT_AMPL_WIDTH),
		24817 => to_signed(22628, LUT_AMPL_WIDTH),
		24818 => to_signed(22626, LUT_AMPL_WIDTH),
		24819 => to_signed(22624, LUT_AMPL_WIDTH),
		24820 => to_signed(22621, LUT_AMPL_WIDTH),
		24821 => to_signed(22619, LUT_AMPL_WIDTH),
		24822 => to_signed(22617, LUT_AMPL_WIDTH),
		24823 => to_signed(22615, LUT_AMPL_WIDTH),
		24824 => to_signed(22612, LUT_AMPL_WIDTH),
		24825 => to_signed(22610, LUT_AMPL_WIDTH),
		24826 => to_signed(22608, LUT_AMPL_WIDTH),
		24827 => to_signed(22606, LUT_AMPL_WIDTH),
		24828 => to_signed(22603, LUT_AMPL_WIDTH),
		24829 => to_signed(22601, LUT_AMPL_WIDTH),
		24830 => to_signed(22599, LUT_AMPL_WIDTH),
		24831 => to_signed(22596, LUT_AMPL_WIDTH),
		24832 => to_signed(22594, LUT_AMPL_WIDTH),
		24833 => to_signed(22592, LUT_AMPL_WIDTH),
		24834 => to_signed(22590, LUT_AMPL_WIDTH),
		24835 => to_signed(22587, LUT_AMPL_WIDTH),
		24836 => to_signed(22585, LUT_AMPL_WIDTH),
		24837 => to_signed(22583, LUT_AMPL_WIDTH),
		24838 => to_signed(22581, LUT_AMPL_WIDTH),
		24839 => to_signed(22578, LUT_AMPL_WIDTH),
		24840 => to_signed(22576, LUT_AMPL_WIDTH),
		24841 => to_signed(22574, LUT_AMPL_WIDTH),
		24842 => to_signed(22571, LUT_AMPL_WIDTH),
		24843 => to_signed(22569, LUT_AMPL_WIDTH),
		24844 => to_signed(22567, LUT_AMPL_WIDTH),
		24845 => to_signed(22565, LUT_AMPL_WIDTH),
		24846 => to_signed(22562, LUT_AMPL_WIDTH),
		24847 => to_signed(22560, LUT_AMPL_WIDTH),
		24848 => to_signed(22558, LUT_AMPL_WIDTH),
		24849 => to_signed(22555, LUT_AMPL_WIDTH),
		24850 => to_signed(22553, LUT_AMPL_WIDTH),
		24851 => to_signed(22551, LUT_AMPL_WIDTH),
		24852 => to_signed(22549, LUT_AMPL_WIDTH),
		24853 => to_signed(22546, LUT_AMPL_WIDTH),
		24854 => to_signed(22544, LUT_AMPL_WIDTH),
		24855 => to_signed(22542, LUT_AMPL_WIDTH),
		24856 => to_signed(22540, LUT_AMPL_WIDTH),
		24857 => to_signed(22537, LUT_AMPL_WIDTH),
		24858 => to_signed(22535, LUT_AMPL_WIDTH),
		24859 => to_signed(22533, LUT_AMPL_WIDTH),
		24860 => to_signed(22530, LUT_AMPL_WIDTH),
		24861 => to_signed(22528, LUT_AMPL_WIDTH),
		24862 => to_signed(22526, LUT_AMPL_WIDTH),
		24863 => to_signed(22524, LUT_AMPL_WIDTH),
		24864 => to_signed(22521, LUT_AMPL_WIDTH),
		24865 => to_signed(22519, LUT_AMPL_WIDTH),
		24866 => to_signed(22517, LUT_AMPL_WIDTH),
		24867 => to_signed(22514, LUT_AMPL_WIDTH),
		24868 => to_signed(22512, LUT_AMPL_WIDTH),
		24869 => to_signed(22510, LUT_AMPL_WIDTH),
		24870 => to_signed(22508, LUT_AMPL_WIDTH),
		24871 => to_signed(22505, LUT_AMPL_WIDTH),
		24872 => to_signed(22503, LUT_AMPL_WIDTH),
		24873 => to_signed(22501, LUT_AMPL_WIDTH),
		24874 => to_signed(22498, LUT_AMPL_WIDTH),
		24875 => to_signed(22496, LUT_AMPL_WIDTH),
		24876 => to_signed(22494, LUT_AMPL_WIDTH),
		24877 => to_signed(22492, LUT_AMPL_WIDTH),
		24878 => to_signed(22489, LUT_AMPL_WIDTH),
		24879 => to_signed(22487, LUT_AMPL_WIDTH),
		24880 => to_signed(22485, LUT_AMPL_WIDTH),
		24881 => to_signed(22482, LUT_AMPL_WIDTH),
		24882 => to_signed(22480, LUT_AMPL_WIDTH),
		24883 => to_signed(22478, LUT_AMPL_WIDTH),
		24884 => to_signed(22476, LUT_AMPL_WIDTH),
		24885 => to_signed(22473, LUT_AMPL_WIDTH),
		24886 => to_signed(22471, LUT_AMPL_WIDTH),
		24887 => to_signed(22469, LUT_AMPL_WIDTH),
		24888 => to_signed(22466, LUT_AMPL_WIDTH),
		24889 => to_signed(22464, LUT_AMPL_WIDTH),
		24890 => to_signed(22462, LUT_AMPL_WIDTH),
		24891 => to_signed(22460, LUT_AMPL_WIDTH),
		24892 => to_signed(22457, LUT_AMPL_WIDTH),
		24893 => to_signed(22455, LUT_AMPL_WIDTH),
		24894 => to_signed(22453, LUT_AMPL_WIDTH),
		24895 => to_signed(22450, LUT_AMPL_WIDTH),
		24896 => to_signed(22448, LUT_AMPL_WIDTH),
		24897 => to_signed(22446, LUT_AMPL_WIDTH),
		24898 => to_signed(22444, LUT_AMPL_WIDTH),
		24899 => to_signed(22441, LUT_AMPL_WIDTH),
		24900 => to_signed(22439, LUT_AMPL_WIDTH),
		24901 => to_signed(22437, LUT_AMPL_WIDTH),
		24902 => to_signed(22434, LUT_AMPL_WIDTH),
		24903 => to_signed(22432, LUT_AMPL_WIDTH),
		24904 => to_signed(22430, LUT_AMPL_WIDTH),
		24905 => to_signed(22428, LUT_AMPL_WIDTH),
		24906 => to_signed(22425, LUT_AMPL_WIDTH),
		24907 => to_signed(22423, LUT_AMPL_WIDTH),
		24908 => to_signed(22421, LUT_AMPL_WIDTH),
		24909 => to_signed(22418, LUT_AMPL_WIDTH),
		24910 => to_signed(22416, LUT_AMPL_WIDTH),
		24911 => to_signed(22414, LUT_AMPL_WIDTH),
		24912 => to_signed(22411, LUT_AMPL_WIDTH),
		24913 => to_signed(22409, LUT_AMPL_WIDTH),
		24914 => to_signed(22407, LUT_AMPL_WIDTH),
		24915 => to_signed(22405, LUT_AMPL_WIDTH),
		24916 => to_signed(22402, LUT_AMPL_WIDTH),
		24917 => to_signed(22400, LUT_AMPL_WIDTH),
		24918 => to_signed(22398, LUT_AMPL_WIDTH),
		24919 => to_signed(22395, LUT_AMPL_WIDTH),
		24920 => to_signed(22393, LUT_AMPL_WIDTH),
		24921 => to_signed(22391, LUT_AMPL_WIDTH),
		24922 => to_signed(22389, LUT_AMPL_WIDTH),
		24923 => to_signed(22386, LUT_AMPL_WIDTH),
		24924 => to_signed(22384, LUT_AMPL_WIDTH),
		24925 => to_signed(22382, LUT_AMPL_WIDTH),
		24926 => to_signed(22379, LUT_AMPL_WIDTH),
		24927 => to_signed(22377, LUT_AMPL_WIDTH),
		24928 => to_signed(22375, LUT_AMPL_WIDTH),
		24929 => to_signed(22373, LUT_AMPL_WIDTH),
		24930 => to_signed(22370, LUT_AMPL_WIDTH),
		24931 => to_signed(22368, LUT_AMPL_WIDTH),
		24932 => to_signed(22366, LUT_AMPL_WIDTH),
		24933 => to_signed(22363, LUT_AMPL_WIDTH),
		24934 => to_signed(22361, LUT_AMPL_WIDTH),
		24935 => to_signed(22359, LUT_AMPL_WIDTH),
		24936 => to_signed(22356, LUT_AMPL_WIDTH),
		24937 => to_signed(22354, LUT_AMPL_WIDTH),
		24938 => to_signed(22352, LUT_AMPL_WIDTH),
		24939 => to_signed(22350, LUT_AMPL_WIDTH),
		24940 => to_signed(22347, LUT_AMPL_WIDTH),
		24941 => to_signed(22345, LUT_AMPL_WIDTH),
		24942 => to_signed(22343, LUT_AMPL_WIDTH),
		24943 => to_signed(22340, LUT_AMPL_WIDTH),
		24944 => to_signed(22338, LUT_AMPL_WIDTH),
		24945 => to_signed(22336, LUT_AMPL_WIDTH),
		24946 => to_signed(22333, LUT_AMPL_WIDTH),
		24947 => to_signed(22331, LUT_AMPL_WIDTH),
		24948 => to_signed(22329, LUT_AMPL_WIDTH),
		24949 => to_signed(22327, LUT_AMPL_WIDTH),
		24950 => to_signed(22324, LUT_AMPL_WIDTH),
		24951 => to_signed(22322, LUT_AMPL_WIDTH),
		24952 => to_signed(22320, LUT_AMPL_WIDTH),
		24953 => to_signed(22317, LUT_AMPL_WIDTH),
		24954 => to_signed(22315, LUT_AMPL_WIDTH),
		24955 => to_signed(22313, LUT_AMPL_WIDTH),
		24956 => to_signed(22310, LUT_AMPL_WIDTH),
		24957 => to_signed(22308, LUT_AMPL_WIDTH),
		24958 => to_signed(22306, LUT_AMPL_WIDTH),
		24959 => to_signed(22304, LUT_AMPL_WIDTH),
		24960 => to_signed(22301, LUT_AMPL_WIDTH),
		24961 => to_signed(22299, LUT_AMPL_WIDTH),
		24962 => to_signed(22297, LUT_AMPL_WIDTH),
		24963 => to_signed(22294, LUT_AMPL_WIDTH),
		24964 => to_signed(22292, LUT_AMPL_WIDTH),
		24965 => to_signed(22290, LUT_AMPL_WIDTH),
		24966 => to_signed(22287, LUT_AMPL_WIDTH),
		24967 => to_signed(22285, LUT_AMPL_WIDTH),
		24968 => to_signed(22283, LUT_AMPL_WIDTH),
		24969 => to_signed(22281, LUT_AMPL_WIDTH),
		24970 => to_signed(22278, LUT_AMPL_WIDTH),
		24971 => to_signed(22276, LUT_AMPL_WIDTH),
		24972 => to_signed(22274, LUT_AMPL_WIDTH),
		24973 => to_signed(22271, LUT_AMPL_WIDTH),
		24974 => to_signed(22269, LUT_AMPL_WIDTH),
		24975 => to_signed(22267, LUT_AMPL_WIDTH),
		24976 => to_signed(22264, LUT_AMPL_WIDTH),
		24977 => to_signed(22262, LUT_AMPL_WIDTH),
		24978 => to_signed(22260, LUT_AMPL_WIDTH),
		24979 => to_signed(22257, LUT_AMPL_WIDTH),
		24980 => to_signed(22255, LUT_AMPL_WIDTH),
		24981 => to_signed(22253, LUT_AMPL_WIDTH),
		24982 => to_signed(22251, LUT_AMPL_WIDTH),
		24983 => to_signed(22248, LUT_AMPL_WIDTH),
		24984 => to_signed(22246, LUT_AMPL_WIDTH),
		24985 => to_signed(22244, LUT_AMPL_WIDTH),
		24986 => to_signed(22241, LUT_AMPL_WIDTH),
		24987 => to_signed(22239, LUT_AMPL_WIDTH),
		24988 => to_signed(22237, LUT_AMPL_WIDTH),
		24989 => to_signed(22234, LUT_AMPL_WIDTH),
		24990 => to_signed(22232, LUT_AMPL_WIDTH),
		24991 => to_signed(22230, LUT_AMPL_WIDTH),
		24992 => to_signed(22227, LUT_AMPL_WIDTH),
		24993 => to_signed(22225, LUT_AMPL_WIDTH),
		24994 => to_signed(22223, LUT_AMPL_WIDTH),
		24995 => to_signed(22221, LUT_AMPL_WIDTH),
		24996 => to_signed(22218, LUT_AMPL_WIDTH),
		24997 => to_signed(22216, LUT_AMPL_WIDTH),
		24998 => to_signed(22214, LUT_AMPL_WIDTH),
		24999 => to_signed(22211, LUT_AMPL_WIDTH),
		25000 => to_signed(22209, LUT_AMPL_WIDTH),
		25001 => to_signed(22207, LUT_AMPL_WIDTH),
		25002 => to_signed(22204, LUT_AMPL_WIDTH),
		25003 => to_signed(22202, LUT_AMPL_WIDTH),
		25004 => to_signed(22200, LUT_AMPL_WIDTH),
		25005 => to_signed(22197, LUT_AMPL_WIDTH),
		25006 => to_signed(22195, LUT_AMPL_WIDTH),
		25007 => to_signed(22193, LUT_AMPL_WIDTH),
		25008 => to_signed(22191, LUT_AMPL_WIDTH),
		25009 => to_signed(22188, LUT_AMPL_WIDTH),
		25010 => to_signed(22186, LUT_AMPL_WIDTH),
		25011 => to_signed(22184, LUT_AMPL_WIDTH),
		25012 => to_signed(22181, LUT_AMPL_WIDTH),
		25013 => to_signed(22179, LUT_AMPL_WIDTH),
		25014 => to_signed(22177, LUT_AMPL_WIDTH),
		25015 => to_signed(22174, LUT_AMPL_WIDTH),
		25016 => to_signed(22172, LUT_AMPL_WIDTH),
		25017 => to_signed(22170, LUT_AMPL_WIDTH),
		25018 => to_signed(22167, LUT_AMPL_WIDTH),
		25019 => to_signed(22165, LUT_AMPL_WIDTH),
		25020 => to_signed(22163, LUT_AMPL_WIDTH),
		25021 => to_signed(22160, LUT_AMPL_WIDTH),
		25022 => to_signed(22158, LUT_AMPL_WIDTH),
		25023 => to_signed(22156, LUT_AMPL_WIDTH),
		25024 => to_signed(22154, LUT_AMPL_WIDTH),
		25025 => to_signed(22151, LUT_AMPL_WIDTH),
		25026 => to_signed(22149, LUT_AMPL_WIDTH),
		25027 => to_signed(22147, LUT_AMPL_WIDTH),
		25028 => to_signed(22144, LUT_AMPL_WIDTH),
		25029 => to_signed(22142, LUT_AMPL_WIDTH),
		25030 => to_signed(22140, LUT_AMPL_WIDTH),
		25031 => to_signed(22137, LUT_AMPL_WIDTH),
		25032 => to_signed(22135, LUT_AMPL_WIDTH),
		25033 => to_signed(22133, LUT_AMPL_WIDTH),
		25034 => to_signed(22130, LUT_AMPL_WIDTH),
		25035 => to_signed(22128, LUT_AMPL_WIDTH),
		25036 => to_signed(22126, LUT_AMPL_WIDTH),
		25037 => to_signed(22123, LUT_AMPL_WIDTH),
		25038 => to_signed(22121, LUT_AMPL_WIDTH),
		25039 => to_signed(22119, LUT_AMPL_WIDTH),
		25040 => to_signed(22116, LUT_AMPL_WIDTH),
		25041 => to_signed(22114, LUT_AMPL_WIDTH),
		25042 => to_signed(22112, LUT_AMPL_WIDTH),
		25043 => to_signed(22110, LUT_AMPL_WIDTH),
		25044 => to_signed(22107, LUT_AMPL_WIDTH),
		25045 => to_signed(22105, LUT_AMPL_WIDTH),
		25046 => to_signed(22103, LUT_AMPL_WIDTH),
		25047 => to_signed(22100, LUT_AMPL_WIDTH),
		25048 => to_signed(22098, LUT_AMPL_WIDTH),
		25049 => to_signed(22096, LUT_AMPL_WIDTH),
		25050 => to_signed(22093, LUT_AMPL_WIDTH),
		25051 => to_signed(22091, LUT_AMPL_WIDTH),
		25052 => to_signed(22089, LUT_AMPL_WIDTH),
		25053 => to_signed(22086, LUT_AMPL_WIDTH),
		25054 => to_signed(22084, LUT_AMPL_WIDTH),
		25055 => to_signed(22082, LUT_AMPL_WIDTH),
		25056 => to_signed(22079, LUT_AMPL_WIDTH),
		25057 => to_signed(22077, LUT_AMPL_WIDTH),
		25058 => to_signed(22075, LUT_AMPL_WIDTH),
		25059 => to_signed(22072, LUT_AMPL_WIDTH),
		25060 => to_signed(22070, LUT_AMPL_WIDTH),
		25061 => to_signed(22068, LUT_AMPL_WIDTH),
		25062 => to_signed(22065, LUT_AMPL_WIDTH),
		25063 => to_signed(22063, LUT_AMPL_WIDTH),
		25064 => to_signed(22061, LUT_AMPL_WIDTH),
		25065 => to_signed(22058, LUT_AMPL_WIDTH),
		25066 => to_signed(22056, LUT_AMPL_WIDTH),
		25067 => to_signed(22054, LUT_AMPL_WIDTH),
		25068 => to_signed(22051, LUT_AMPL_WIDTH),
		25069 => to_signed(22049, LUT_AMPL_WIDTH),
		25070 => to_signed(22047, LUT_AMPL_WIDTH),
		25071 => to_signed(22045, LUT_AMPL_WIDTH),
		25072 => to_signed(22042, LUT_AMPL_WIDTH),
		25073 => to_signed(22040, LUT_AMPL_WIDTH),
		25074 => to_signed(22038, LUT_AMPL_WIDTH),
		25075 => to_signed(22035, LUT_AMPL_WIDTH),
		25076 => to_signed(22033, LUT_AMPL_WIDTH),
		25077 => to_signed(22031, LUT_AMPL_WIDTH),
		25078 => to_signed(22028, LUT_AMPL_WIDTH),
		25079 => to_signed(22026, LUT_AMPL_WIDTH),
		25080 => to_signed(22024, LUT_AMPL_WIDTH),
		25081 => to_signed(22021, LUT_AMPL_WIDTH),
		25082 => to_signed(22019, LUT_AMPL_WIDTH),
		25083 => to_signed(22017, LUT_AMPL_WIDTH),
		25084 => to_signed(22014, LUT_AMPL_WIDTH),
		25085 => to_signed(22012, LUT_AMPL_WIDTH),
		25086 => to_signed(22010, LUT_AMPL_WIDTH),
		25087 => to_signed(22007, LUT_AMPL_WIDTH),
		25088 => to_signed(22005, LUT_AMPL_WIDTH),
		25089 => to_signed(22003, LUT_AMPL_WIDTH),
		25090 => to_signed(22000, LUT_AMPL_WIDTH),
		25091 => to_signed(21998, LUT_AMPL_WIDTH),
		25092 => to_signed(21996, LUT_AMPL_WIDTH),
		25093 => to_signed(21993, LUT_AMPL_WIDTH),
		25094 => to_signed(21991, LUT_AMPL_WIDTH),
		25095 => to_signed(21989, LUT_AMPL_WIDTH),
		25096 => to_signed(21986, LUT_AMPL_WIDTH),
		25097 => to_signed(21984, LUT_AMPL_WIDTH),
		25098 => to_signed(21982, LUT_AMPL_WIDTH),
		25099 => to_signed(21979, LUT_AMPL_WIDTH),
		25100 => to_signed(21977, LUT_AMPL_WIDTH),
		25101 => to_signed(21975, LUT_AMPL_WIDTH),
		25102 => to_signed(21972, LUT_AMPL_WIDTH),
		25103 => to_signed(21970, LUT_AMPL_WIDTH),
		25104 => to_signed(21968, LUT_AMPL_WIDTH),
		25105 => to_signed(21965, LUT_AMPL_WIDTH),
		25106 => to_signed(21963, LUT_AMPL_WIDTH),
		25107 => to_signed(21961, LUT_AMPL_WIDTH),
		25108 => to_signed(21958, LUT_AMPL_WIDTH),
		25109 => to_signed(21956, LUT_AMPL_WIDTH),
		25110 => to_signed(21954, LUT_AMPL_WIDTH),
		25111 => to_signed(21951, LUT_AMPL_WIDTH),
		25112 => to_signed(21949, LUT_AMPL_WIDTH),
		25113 => to_signed(21947, LUT_AMPL_WIDTH),
		25114 => to_signed(21944, LUT_AMPL_WIDTH),
		25115 => to_signed(21942, LUT_AMPL_WIDTH),
		25116 => to_signed(21940, LUT_AMPL_WIDTH),
		25117 => to_signed(21937, LUT_AMPL_WIDTH),
		25118 => to_signed(21935, LUT_AMPL_WIDTH),
		25119 => to_signed(21933, LUT_AMPL_WIDTH),
		25120 => to_signed(21930, LUT_AMPL_WIDTH),
		25121 => to_signed(21928, LUT_AMPL_WIDTH),
		25122 => to_signed(21926, LUT_AMPL_WIDTH),
		25123 => to_signed(21923, LUT_AMPL_WIDTH),
		25124 => to_signed(21921, LUT_AMPL_WIDTH),
		25125 => to_signed(21919, LUT_AMPL_WIDTH),
		25126 => to_signed(21916, LUT_AMPL_WIDTH),
		25127 => to_signed(21914, LUT_AMPL_WIDTH),
		25128 => to_signed(21912, LUT_AMPL_WIDTH),
		25129 => to_signed(21909, LUT_AMPL_WIDTH),
		25130 => to_signed(21907, LUT_AMPL_WIDTH),
		25131 => to_signed(21905, LUT_AMPL_WIDTH),
		25132 => to_signed(21902, LUT_AMPL_WIDTH),
		25133 => to_signed(21900, LUT_AMPL_WIDTH),
		25134 => to_signed(21898, LUT_AMPL_WIDTH),
		25135 => to_signed(21895, LUT_AMPL_WIDTH),
		25136 => to_signed(21893, LUT_AMPL_WIDTH),
		25137 => to_signed(21891, LUT_AMPL_WIDTH),
		25138 => to_signed(21888, LUT_AMPL_WIDTH),
		25139 => to_signed(21886, LUT_AMPL_WIDTH),
		25140 => to_signed(21884, LUT_AMPL_WIDTH),
		25141 => to_signed(21881, LUT_AMPL_WIDTH),
		25142 => to_signed(21879, LUT_AMPL_WIDTH),
		25143 => to_signed(21877, LUT_AMPL_WIDTH),
		25144 => to_signed(21874, LUT_AMPL_WIDTH),
		25145 => to_signed(21872, LUT_AMPL_WIDTH),
		25146 => to_signed(21870, LUT_AMPL_WIDTH),
		25147 => to_signed(21867, LUT_AMPL_WIDTH),
		25148 => to_signed(21865, LUT_AMPL_WIDTH),
		25149 => to_signed(21863, LUT_AMPL_WIDTH),
		25150 => to_signed(21860, LUT_AMPL_WIDTH),
		25151 => to_signed(21858, LUT_AMPL_WIDTH),
		25152 => to_signed(21856, LUT_AMPL_WIDTH),
		25153 => to_signed(21853, LUT_AMPL_WIDTH),
		25154 => to_signed(21851, LUT_AMPL_WIDTH),
		25155 => to_signed(21849, LUT_AMPL_WIDTH),
		25156 => to_signed(21846, LUT_AMPL_WIDTH),
		25157 => to_signed(21844, LUT_AMPL_WIDTH),
		25158 => to_signed(21842, LUT_AMPL_WIDTH),
		25159 => to_signed(21839, LUT_AMPL_WIDTH),
		25160 => to_signed(21837, LUT_AMPL_WIDTH),
		25161 => to_signed(21835, LUT_AMPL_WIDTH),
		25162 => to_signed(21832, LUT_AMPL_WIDTH),
		25163 => to_signed(21830, LUT_AMPL_WIDTH),
		25164 => to_signed(21827, LUT_AMPL_WIDTH),
		25165 => to_signed(21825, LUT_AMPL_WIDTH),
		25166 => to_signed(21823, LUT_AMPL_WIDTH),
		25167 => to_signed(21820, LUT_AMPL_WIDTH),
		25168 => to_signed(21818, LUT_AMPL_WIDTH),
		25169 => to_signed(21816, LUT_AMPL_WIDTH),
		25170 => to_signed(21813, LUT_AMPL_WIDTH),
		25171 => to_signed(21811, LUT_AMPL_WIDTH),
		25172 => to_signed(21809, LUT_AMPL_WIDTH),
		25173 => to_signed(21806, LUT_AMPL_WIDTH),
		25174 => to_signed(21804, LUT_AMPL_WIDTH),
		25175 => to_signed(21802, LUT_AMPL_WIDTH),
		25176 => to_signed(21799, LUT_AMPL_WIDTH),
		25177 => to_signed(21797, LUT_AMPL_WIDTH),
		25178 => to_signed(21795, LUT_AMPL_WIDTH),
		25179 => to_signed(21792, LUT_AMPL_WIDTH),
		25180 => to_signed(21790, LUT_AMPL_WIDTH),
		25181 => to_signed(21788, LUT_AMPL_WIDTH),
		25182 => to_signed(21785, LUT_AMPL_WIDTH),
		25183 => to_signed(21783, LUT_AMPL_WIDTH),
		25184 => to_signed(21781, LUT_AMPL_WIDTH),
		25185 => to_signed(21778, LUT_AMPL_WIDTH),
		25186 => to_signed(21776, LUT_AMPL_WIDTH),
		25187 => to_signed(21774, LUT_AMPL_WIDTH),
		25188 => to_signed(21771, LUT_AMPL_WIDTH),
		25189 => to_signed(21769, LUT_AMPL_WIDTH),
		25190 => to_signed(21766, LUT_AMPL_WIDTH),
		25191 => to_signed(21764, LUT_AMPL_WIDTH),
		25192 => to_signed(21762, LUT_AMPL_WIDTH),
		25193 => to_signed(21759, LUT_AMPL_WIDTH),
		25194 => to_signed(21757, LUT_AMPL_WIDTH),
		25195 => to_signed(21755, LUT_AMPL_WIDTH),
		25196 => to_signed(21752, LUT_AMPL_WIDTH),
		25197 => to_signed(21750, LUT_AMPL_WIDTH),
		25198 => to_signed(21748, LUT_AMPL_WIDTH),
		25199 => to_signed(21745, LUT_AMPL_WIDTH),
		25200 => to_signed(21743, LUT_AMPL_WIDTH),
		25201 => to_signed(21741, LUT_AMPL_WIDTH),
		25202 => to_signed(21738, LUT_AMPL_WIDTH),
		25203 => to_signed(21736, LUT_AMPL_WIDTH),
		25204 => to_signed(21734, LUT_AMPL_WIDTH),
		25205 => to_signed(21731, LUT_AMPL_WIDTH),
		25206 => to_signed(21729, LUT_AMPL_WIDTH),
		25207 => to_signed(21727, LUT_AMPL_WIDTH),
		25208 => to_signed(21724, LUT_AMPL_WIDTH),
		25209 => to_signed(21722, LUT_AMPL_WIDTH),
		25210 => to_signed(21719, LUT_AMPL_WIDTH),
		25211 => to_signed(21717, LUT_AMPL_WIDTH),
		25212 => to_signed(21715, LUT_AMPL_WIDTH),
		25213 => to_signed(21712, LUT_AMPL_WIDTH),
		25214 => to_signed(21710, LUT_AMPL_WIDTH),
		25215 => to_signed(21708, LUT_AMPL_WIDTH),
		25216 => to_signed(21705, LUT_AMPL_WIDTH),
		25217 => to_signed(21703, LUT_AMPL_WIDTH),
		25218 => to_signed(21701, LUT_AMPL_WIDTH),
		25219 => to_signed(21698, LUT_AMPL_WIDTH),
		25220 => to_signed(21696, LUT_AMPL_WIDTH),
		25221 => to_signed(21694, LUT_AMPL_WIDTH),
		25222 => to_signed(21691, LUT_AMPL_WIDTH),
		25223 => to_signed(21689, LUT_AMPL_WIDTH),
		25224 => to_signed(21687, LUT_AMPL_WIDTH),
		25225 => to_signed(21684, LUT_AMPL_WIDTH),
		25226 => to_signed(21682, LUT_AMPL_WIDTH),
		25227 => to_signed(21679, LUT_AMPL_WIDTH),
		25228 => to_signed(21677, LUT_AMPL_WIDTH),
		25229 => to_signed(21675, LUT_AMPL_WIDTH),
		25230 => to_signed(21672, LUT_AMPL_WIDTH),
		25231 => to_signed(21670, LUT_AMPL_WIDTH),
		25232 => to_signed(21668, LUT_AMPL_WIDTH),
		25233 => to_signed(21665, LUT_AMPL_WIDTH),
		25234 => to_signed(21663, LUT_AMPL_WIDTH),
		25235 => to_signed(21661, LUT_AMPL_WIDTH),
		25236 => to_signed(21658, LUT_AMPL_WIDTH),
		25237 => to_signed(21656, LUT_AMPL_WIDTH),
		25238 => to_signed(21654, LUT_AMPL_WIDTH),
		25239 => to_signed(21651, LUT_AMPL_WIDTH),
		25240 => to_signed(21649, LUT_AMPL_WIDTH),
		25241 => to_signed(21646, LUT_AMPL_WIDTH),
		25242 => to_signed(21644, LUT_AMPL_WIDTH),
		25243 => to_signed(21642, LUT_AMPL_WIDTH),
		25244 => to_signed(21639, LUT_AMPL_WIDTH),
		25245 => to_signed(21637, LUT_AMPL_WIDTH),
		25246 => to_signed(21635, LUT_AMPL_WIDTH),
		25247 => to_signed(21632, LUT_AMPL_WIDTH),
		25248 => to_signed(21630, LUT_AMPL_WIDTH),
		25249 => to_signed(21628, LUT_AMPL_WIDTH),
		25250 => to_signed(21625, LUT_AMPL_WIDTH),
		25251 => to_signed(21623, LUT_AMPL_WIDTH),
		25252 => to_signed(21621, LUT_AMPL_WIDTH),
		25253 => to_signed(21618, LUT_AMPL_WIDTH),
		25254 => to_signed(21616, LUT_AMPL_WIDTH),
		25255 => to_signed(21613, LUT_AMPL_WIDTH),
		25256 => to_signed(21611, LUT_AMPL_WIDTH),
		25257 => to_signed(21609, LUT_AMPL_WIDTH),
		25258 => to_signed(21606, LUT_AMPL_WIDTH),
		25259 => to_signed(21604, LUT_AMPL_WIDTH),
		25260 => to_signed(21602, LUT_AMPL_WIDTH),
		25261 => to_signed(21599, LUT_AMPL_WIDTH),
		25262 => to_signed(21597, LUT_AMPL_WIDTH),
		25263 => to_signed(21595, LUT_AMPL_WIDTH),
		25264 => to_signed(21592, LUT_AMPL_WIDTH),
		25265 => to_signed(21590, LUT_AMPL_WIDTH),
		25266 => to_signed(21587, LUT_AMPL_WIDTH),
		25267 => to_signed(21585, LUT_AMPL_WIDTH),
		25268 => to_signed(21583, LUT_AMPL_WIDTH),
		25269 => to_signed(21580, LUT_AMPL_WIDTH),
		25270 => to_signed(21578, LUT_AMPL_WIDTH),
		25271 => to_signed(21576, LUT_AMPL_WIDTH),
		25272 => to_signed(21573, LUT_AMPL_WIDTH),
		25273 => to_signed(21571, LUT_AMPL_WIDTH),
		25274 => to_signed(21569, LUT_AMPL_WIDTH),
		25275 => to_signed(21566, LUT_AMPL_WIDTH),
		25276 => to_signed(21564, LUT_AMPL_WIDTH),
		25277 => to_signed(21561, LUT_AMPL_WIDTH),
		25278 => to_signed(21559, LUT_AMPL_WIDTH),
		25279 => to_signed(21557, LUT_AMPL_WIDTH),
		25280 => to_signed(21554, LUT_AMPL_WIDTH),
		25281 => to_signed(21552, LUT_AMPL_WIDTH),
		25282 => to_signed(21550, LUT_AMPL_WIDTH),
		25283 => to_signed(21547, LUT_AMPL_WIDTH),
		25284 => to_signed(21545, LUT_AMPL_WIDTH),
		25285 => to_signed(21543, LUT_AMPL_WIDTH),
		25286 => to_signed(21540, LUT_AMPL_WIDTH),
		25287 => to_signed(21538, LUT_AMPL_WIDTH),
		25288 => to_signed(21535, LUT_AMPL_WIDTH),
		25289 => to_signed(21533, LUT_AMPL_WIDTH),
		25290 => to_signed(21531, LUT_AMPL_WIDTH),
		25291 => to_signed(21528, LUT_AMPL_WIDTH),
		25292 => to_signed(21526, LUT_AMPL_WIDTH),
		25293 => to_signed(21524, LUT_AMPL_WIDTH),
		25294 => to_signed(21521, LUT_AMPL_WIDTH),
		25295 => to_signed(21519, LUT_AMPL_WIDTH),
		25296 => to_signed(21516, LUT_AMPL_WIDTH),
		25297 => to_signed(21514, LUT_AMPL_WIDTH),
		25298 => to_signed(21512, LUT_AMPL_WIDTH),
		25299 => to_signed(21509, LUT_AMPL_WIDTH),
		25300 => to_signed(21507, LUT_AMPL_WIDTH),
		25301 => to_signed(21505, LUT_AMPL_WIDTH),
		25302 => to_signed(21502, LUT_AMPL_WIDTH),
		25303 => to_signed(21500, LUT_AMPL_WIDTH),
		25304 => to_signed(21498, LUT_AMPL_WIDTH),
		25305 => to_signed(21495, LUT_AMPL_WIDTH),
		25306 => to_signed(21493, LUT_AMPL_WIDTH),
		25307 => to_signed(21490, LUT_AMPL_WIDTH),
		25308 => to_signed(21488, LUT_AMPL_WIDTH),
		25309 => to_signed(21486, LUT_AMPL_WIDTH),
		25310 => to_signed(21483, LUT_AMPL_WIDTH),
		25311 => to_signed(21481, LUT_AMPL_WIDTH),
		25312 => to_signed(21479, LUT_AMPL_WIDTH),
		25313 => to_signed(21476, LUT_AMPL_WIDTH),
		25314 => to_signed(21474, LUT_AMPL_WIDTH),
		25315 => to_signed(21471, LUT_AMPL_WIDTH),
		25316 => to_signed(21469, LUT_AMPL_WIDTH),
		25317 => to_signed(21467, LUT_AMPL_WIDTH),
		25318 => to_signed(21464, LUT_AMPL_WIDTH),
		25319 => to_signed(21462, LUT_AMPL_WIDTH),
		25320 => to_signed(21460, LUT_AMPL_WIDTH),
		25321 => to_signed(21457, LUT_AMPL_WIDTH),
		25322 => to_signed(21455, LUT_AMPL_WIDTH),
		25323 => to_signed(21452, LUT_AMPL_WIDTH),
		25324 => to_signed(21450, LUT_AMPL_WIDTH),
		25325 => to_signed(21448, LUT_AMPL_WIDTH),
		25326 => to_signed(21445, LUT_AMPL_WIDTH),
		25327 => to_signed(21443, LUT_AMPL_WIDTH),
		25328 => to_signed(21441, LUT_AMPL_WIDTH),
		25329 => to_signed(21438, LUT_AMPL_WIDTH),
		25330 => to_signed(21436, LUT_AMPL_WIDTH),
		25331 => to_signed(21433, LUT_AMPL_WIDTH),
		25332 => to_signed(21431, LUT_AMPL_WIDTH),
		25333 => to_signed(21429, LUT_AMPL_WIDTH),
		25334 => to_signed(21426, LUT_AMPL_WIDTH),
		25335 => to_signed(21424, LUT_AMPL_WIDTH),
		25336 => to_signed(21422, LUT_AMPL_WIDTH),
		25337 => to_signed(21419, LUT_AMPL_WIDTH),
		25338 => to_signed(21417, LUT_AMPL_WIDTH),
		25339 => to_signed(21414, LUT_AMPL_WIDTH),
		25340 => to_signed(21412, LUT_AMPL_WIDTH),
		25341 => to_signed(21410, LUT_AMPL_WIDTH),
		25342 => to_signed(21407, LUT_AMPL_WIDTH),
		25343 => to_signed(21405, LUT_AMPL_WIDTH),
		25344 => to_signed(21403, LUT_AMPL_WIDTH),
		25345 => to_signed(21400, LUT_AMPL_WIDTH),
		25346 => to_signed(21398, LUT_AMPL_WIDTH),
		25347 => to_signed(21395, LUT_AMPL_WIDTH),
		25348 => to_signed(21393, LUT_AMPL_WIDTH),
		25349 => to_signed(21391, LUT_AMPL_WIDTH),
		25350 => to_signed(21388, LUT_AMPL_WIDTH),
		25351 => to_signed(21386, LUT_AMPL_WIDTH),
		25352 => to_signed(21383, LUT_AMPL_WIDTH),
		25353 => to_signed(21381, LUT_AMPL_WIDTH),
		25354 => to_signed(21379, LUT_AMPL_WIDTH),
		25355 => to_signed(21376, LUT_AMPL_WIDTH),
		25356 => to_signed(21374, LUT_AMPL_WIDTH),
		25357 => to_signed(21372, LUT_AMPL_WIDTH),
		25358 => to_signed(21369, LUT_AMPL_WIDTH),
		25359 => to_signed(21367, LUT_AMPL_WIDTH),
		25360 => to_signed(21364, LUT_AMPL_WIDTH),
		25361 => to_signed(21362, LUT_AMPL_WIDTH),
		25362 => to_signed(21360, LUT_AMPL_WIDTH),
		25363 => to_signed(21357, LUT_AMPL_WIDTH),
		25364 => to_signed(21355, LUT_AMPL_WIDTH),
		25365 => to_signed(21353, LUT_AMPL_WIDTH),
		25366 => to_signed(21350, LUT_AMPL_WIDTH),
		25367 => to_signed(21348, LUT_AMPL_WIDTH),
		25368 => to_signed(21345, LUT_AMPL_WIDTH),
		25369 => to_signed(21343, LUT_AMPL_WIDTH),
		25370 => to_signed(21341, LUT_AMPL_WIDTH),
		25371 => to_signed(21338, LUT_AMPL_WIDTH),
		25372 => to_signed(21336, LUT_AMPL_WIDTH),
		25373 => to_signed(21333, LUT_AMPL_WIDTH),
		25374 => to_signed(21331, LUT_AMPL_WIDTH),
		25375 => to_signed(21329, LUT_AMPL_WIDTH),
		25376 => to_signed(21326, LUT_AMPL_WIDTH),
		25377 => to_signed(21324, LUT_AMPL_WIDTH),
		25378 => to_signed(21322, LUT_AMPL_WIDTH),
		25379 => to_signed(21319, LUT_AMPL_WIDTH),
		25380 => to_signed(21317, LUT_AMPL_WIDTH),
		25381 => to_signed(21314, LUT_AMPL_WIDTH),
		25382 => to_signed(21312, LUT_AMPL_WIDTH),
		25383 => to_signed(21310, LUT_AMPL_WIDTH),
		25384 => to_signed(21307, LUT_AMPL_WIDTH),
		25385 => to_signed(21305, LUT_AMPL_WIDTH),
		25386 => to_signed(21302, LUT_AMPL_WIDTH),
		25387 => to_signed(21300, LUT_AMPL_WIDTH),
		25388 => to_signed(21298, LUT_AMPL_WIDTH),
		25389 => to_signed(21295, LUT_AMPL_WIDTH),
		25390 => to_signed(21293, LUT_AMPL_WIDTH),
		25391 => to_signed(21290, LUT_AMPL_WIDTH),
		25392 => to_signed(21288, LUT_AMPL_WIDTH),
		25393 => to_signed(21286, LUT_AMPL_WIDTH),
		25394 => to_signed(21283, LUT_AMPL_WIDTH),
		25395 => to_signed(21281, LUT_AMPL_WIDTH),
		25396 => to_signed(21279, LUT_AMPL_WIDTH),
		25397 => to_signed(21276, LUT_AMPL_WIDTH),
		25398 => to_signed(21274, LUT_AMPL_WIDTH),
		25399 => to_signed(21271, LUT_AMPL_WIDTH),
		25400 => to_signed(21269, LUT_AMPL_WIDTH),
		25401 => to_signed(21267, LUT_AMPL_WIDTH),
		25402 => to_signed(21264, LUT_AMPL_WIDTH),
		25403 => to_signed(21262, LUT_AMPL_WIDTH),
		25404 => to_signed(21259, LUT_AMPL_WIDTH),
		25405 => to_signed(21257, LUT_AMPL_WIDTH),
		25406 => to_signed(21255, LUT_AMPL_WIDTH),
		25407 => to_signed(21252, LUT_AMPL_WIDTH),
		25408 => to_signed(21250, LUT_AMPL_WIDTH),
		25409 => to_signed(21247, LUT_AMPL_WIDTH),
		25410 => to_signed(21245, LUT_AMPL_WIDTH),
		25411 => to_signed(21243, LUT_AMPL_WIDTH),
		25412 => to_signed(21240, LUT_AMPL_WIDTH),
		25413 => to_signed(21238, LUT_AMPL_WIDTH),
		25414 => to_signed(21236, LUT_AMPL_WIDTH),
		25415 => to_signed(21233, LUT_AMPL_WIDTH),
		25416 => to_signed(21231, LUT_AMPL_WIDTH),
		25417 => to_signed(21228, LUT_AMPL_WIDTH),
		25418 => to_signed(21226, LUT_AMPL_WIDTH),
		25419 => to_signed(21224, LUT_AMPL_WIDTH),
		25420 => to_signed(21221, LUT_AMPL_WIDTH),
		25421 => to_signed(21219, LUT_AMPL_WIDTH),
		25422 => to_signed(21216, LUT_AMPL_WIDTH),
		25423 => to_signed(21214, LUT_AMPL_WIDTH),
		25424 => to_signed(21212, LUT_AMPL_WIDTH),
		25425 => to_signed(21209, LUT_AMPL_WIDTH),
		25426 => to_signed(21207, LUT_AMPL_WIDTH),
		25427 => to_signed(21204, LUT_AMPL_WIDTH),
		25428 => to_signed(21202, LUT_AMPL_WIDTH),
		25429 => to_signed(21200, LUT_AMPL_WIDTH),
		25430 => to_signed(21197, LUT_AMPL_WIDTH),
		25431 => to_signed(21195, LUT_AMPL_WIDTH),
		25432 => to_signed(21192, LUT_AMPL_WIDTH),
		25433 => to_signed(21190, LUT_AMPL_WIDTH),
		25434 => to_signed(21188, LUT_AMPL_WIDTH),
		25435 => to_signed(21185, LUT_AMPL_WIDTH),
		25436 => to_signed(21183, LUT_AMPL_WIDTH),
		25437 => to_signed(21180, LUT_AMPL_WIDTH),
		25438 => to_signed(21178, LUT_AMPL_WIDTH),
		25439 => to_signed(21176, LUT_AMPL_WIDTH),
		25440 => to_signed(21173, LUT_AMPL_WIDTH),
		25441 => to_signed(21171, LUT_AMPL_WIDTH),
		25442 => to_signed(21168, LUT_AMPL_WIDTH),
		25443 => to_signed(21166, LUT_AMPL_WIDTH),
		25444 => to_signed(21164, LUT_AMPL_WIDTH),
		25445 => to_signed(21161, LUT_AMPL_WIDTH),
		25446 => to_signed(21159, LUT_AMPL_WIDTH),
		25447 => to_signed(21156, LUT_AMPL_WIDTH),
		25448 => to_signed(21154, LUT_AMPL_WIDTH),
		25449 => to_signed(21152, LUT_AMPL_WIDTH),
		25450 => to_signed(21149, LUT_AMPL_WIDTH),
		25451 => to_signed(21147, LUT_AMPL_WIDTH),
		25452 => to_signed(21144, LUT_AMPL_WIDTH),
		25453 => to_signed(21142, LUT_AMPL_WIDTH),
		25454 => to_signed(21140, LUT_AMPL_WIDTH),
		25455 => to_signed(21137, LUT_AMPL_WIDTH),
		25456 => to_signed(21135, LUT_AMPL_WIDTH),
		25457 => to_signed(21132, LUT_AMPL_WIDTH),
		25458 => to_signed(21130, LUT_AMPL_WIDTH),
		25459 => to_signed(21128, LUT_AMPL_WIDTH),
		25460 => to_signed(21125, LUT_AMPL_WIDTH),
		25461 => to_signed(21123, LUT_AMPL_WIDTH),
		25462 => to_signed(21120, LUT_AMPL_WIDTH),
		25463 => to_signed(21118, LUT_AMPL_WIDTH),
		25464 => to_signed(21116, LUT_AMPL_WIDTH),
		25465 => to_signed(21113, LUT_AMPL_WIDTH),
		25466 => to_signed(21111, LUT_AMPL_WIDTH),
		25467 => to_signed(21108, LUT_AMPL_WIDTH),
		25468 => to_signed(21106, LUT_AMPL_WIDTH),
		25469 => to_signed(21104, LUT_AMPL_WIDTH),
		25470 => to_signed(21101, LUT_AMPL_WIDTH),
		25471 => to_signed(21099, LUT_AMPL_WIDTH),
		25472 => to_signed(21096, LUT_AMPL_WIDTH),
		25473 => to_signed(21094, LUT_AMPL_WIDTH),
		25474 => to_signed(21092, LUT_AMPL_WIDTH),
		25475 => to_signed(21089, LUT_AMPL_WIDTH),
		25476 => to_signed(21087, LUT_AMPL_WIDTH),
		25477 => to_signed(21084, LUT_AMPL_WIDTH),
		25478 => to_signed(21082, LUT_AMPL_WIDTH),
		25479 => to_signed(21080, LUT_AMPL_WIDTH),
		25480 => to_signed(21077, LUT_AMPL_WIDTH),
		25481 => to_signed(21075, LUT_AMPL_WIDTH),
		25482 => to_signed(21072, LUT_AMPL_WIDTH),
		25483 => to_signed(21070, LUT_AMPL_WIDTH),
		25484 => to_signed(21068, LUT_AMPL_WIDTH),
		25485 => to_signed(21065, LUT_AMPL_WIDTH),
		25486 => to_signed(21063, LUT_AMPL_WIDTH),
		25487 => to_signed(21060, LUT_AMPL_WIDTH),
		25488 => to_signed(21058, LUT_AMPL_WIDTH),
		25489 => to_signed(21056, LUT_AMPL_WIDTH),
		25490 => to_signed(21053, LUT_AMPL_WIDTH),
		25491 => to_signed(21051, LUT_AMPL_WIDTH),
		25492 => to_signed(21048, LUT_AMPL_WIDTH),
		25493 => to_signed(21046, LUT_AMPL_WIDTH),
		25494 => to_signed(21043, LUT_AMPL_WIDTH),
		25495 => to_signed(21041, LUT_AMPL_WIDTH),
		25496 => to_signed(21039, LUT_AMPL_WIDTH),
		25497 => to_signed(21036, LUT_AMPL_WIDTH),
		25498 => to_signed(21034, LUT_AMPL_WIDTH),
		25499 => to_signed(21031, LUT_AMPL_WIDTH),
		25500 => to_signed(21029, LUT_AMPL_WIDTH),
		25501 => to_signed(21027, LUT_AMPL_WIDTH),
		25502 => to_signed(21024, LUT_AMPL_WIDTH),
		25503 => to_signed(21022, LUT_AMPL_WIDTH),
		25504 => to_signed(21019, LUT_AMPL_WIDTH),
		25505 => to_signed(21017, LUT_AMPL_WIDTH),
		25506 => to_signed(21015, LUT_AMPL_WIDTH),
		25507 => to_signed(21012, LUT_AMPL_WIDTH),
		25508 => to_signed(21010, LUT_AMPL_WIDTH),
		25509 => to_signed(21007, LUT_AMPL_WIDTH),
		25510 => to_signed(21005, LUT_AMPL_WIDTH),
		25511 => to_signed(21003, LUT_AMPL_WIDTH),
		25512 => to_signed(21000, LUT_AMPL_WIDTH),
		25513 => to_signed(20998, LUT_AMPL_WIDTH),
		25514 => to_signed(20995, LUT_AMPL_WIDTH),
		25515 => to_signed(20993, LUT_AMPL_WIDTH),
		25516 => to_signed(20990, LUT_AMPL_WIDTH),
		25517 => to_signed(20988, LUT_AMPL_WIDTH),
		25518 => to_signed(20986, LUT_AMPL_WIDTH),
		25519 => to_signed(20983, LUT_AMPL_WIDTH),
		25520 => to_signed(20981, LUT_AMPL_WIDTH),
		25521 => to_signed(20978, LUT_AMPL_WIDTH),
		25522 => to_signed(20976, LUT_AMPL_WIDTH),
		25523 => to_signed(20974, LUT_AMPL_WIDTH),
		25524 => to_signed(20971, LUT_AMPL_WIDTH),
		25525 => to_signed(20969, LUT_AMPL_WIDTH),
		25526 => to_signed(20966, LUT_AMPL_WIDTH),
		25527 => to_signed(20964, LUT_AMPL_WIDTH),
		25528 => to_signed(20962, LUT_AMPL_WIDTH),
		25529 => to_signed(20959, LUT_AMPL_WIDTH),
		25530 => to_signed(20957, LUT_AMPL_WIDTH),
		25531 => to_signed(20954, LUT_AMPL_WIDTH),
		25532 => to_signed(20952, LUT_AMPL_WIDTH),
		25533 => to_signed(20949, LUT_AMPL_WIDTH),
		25534 => to_signed(20947, LUT_AMPL_WIDTH),
		25535 => to_signed(20945, LUT_AMPL_WIDTH),
		25536 => to_signed(20942, LUT_AMPL_WIDTH),
		25537 => to_signed(20940, LUT_AMPL_WIDTH),
		25538 => to_signed(20937, LUT_AMPL_WIDTH),
		25539 => to_signed(20935, LUT_AMPL_WIDTH),
		25540 => to_signed(20933, LUT_AMPL_WIDTH),
		25541 => to_signed(20930, LUT_AMPL_WIDTH),
		25542 => to_signed(20928, LUT_AMPL_WIDTH),
		25543 => to_signed(20925, LUT_AMPL_WIDTH),
		25544 => to_signed(20923, LUT_AMPL_WIDTH),
		25545 => to_signed(20920, LUT_AMPL_WIDTH),
		25546 => to_signed(20918, LUT_AMPL_WIDTH),
		25547 => to_signed(20916, LUT_AMPL_WIDTH),
		25548 => to_signed(20913, LUT_AMPL_WIDTH),
		25549 => to_signed(20911, LUT_AMPL_WIDTH),
		25550 => to_signed(20908, LUT_AMPL_WIDTH),
		25551 => to_signed(20906, LUT_AMPL_WIDTH),
		25552 => to_signed(20904, LUT_AMPL_WIDTH),
		25553 => to_signed(20901, LUT_AMPL_WIDTH),
		25554 => to_signed(20899, LUT_AMPL_WIDTH),
		25555 => to_signed(20896, LUT_AMPL_WIDTH),
		25556 => to_signed(20894, LUT_AMPL_WIDTH),
		25557 => to_signed(20891, LUT_AMPL_WIDTH),
		25558 => to_signed(20889, LUT_AMPL_WIDTH),
		25559 => to_signed(20887, LUT_AMPL_WIDTH),
		25560 => to_signed(20884, LUT_AMPL_WIDTH),
		25561 => to_signed(20882, LUT_AMPL_WIDTH),
		25562 => to_signed(20879, LUT_AMPL_WIDTH),
		25563 => to_signed(20877, LUT_AMPL_WIDTH),
		25564 => to_signed(20874, LUT_AMPL_WIDTH),
		25565 => to_signed(20872, LUT_AMPL_WIDTH),
		25566 => to_signed(20870, LUT_AMPL_WIDTH),
		25567 => to_signed(20867, LUT_AMPL_WIDTH),
		25568 => to_signed(20865, LUT_AMPL_WIDTH),
		25569 => to_signed(20862, LUT_AMPL_WIDTH),
		25570 => to_signed(20860, LUT_AMPL_WIDTH),
		25571 => to_signed(20858, LUT_AMPL_WIDTH),
		25572 => to_signed(20855, LUT_AMPL_WIDTH),
		25573 => to_signed(20853, LUT_AMPL_WIDTH),
		25574 => to_signed(20850, LUT_AMPL_WIDTH),
		25575 => to_signed(20848, LUT_AMPL_WIDTH),
		25576 => to_signed(20845, LUT_AMPL_WIDTH),
		25577 => to_signed(20843, LUT_AMPL_WIDTH),
		25578 => to_signed(20841, LUT_AMPL_WIDTH),
		25579 => to_signed(20838, LUT_AMPL_WIDTH),
		25580 => to_signed(20836, LUT_AMPL_WIDTH),
		25581 => to_signed(20833, LUT_AMPL_WIDTH),
		25582 => to_signed(20831, LUT_AMPL_WIDTH),
		25583 => to_signed(20828, LUT_AMPL_WIDTH),
		25584 => to_signed(20826, LUT_AMPL_WIDTH),
		25585 => to_signed(20824, LUT_AMPL_WIDTH),
		25586 => to_signed(20821, LUT_AMPL_WIDTH),
		25587 => to_signed(20819, LUT_AMPL_WIDTH),
		25588 => to_signed(20816, LUT_AMPL_WIDTH),
		25589 => to_signed(20814, LUT_AMPL_WIDTH),
		25590 => to_signed(20811, LUT_AMPL_WIDTH),
		25591 => to_signed(20809, LUT_AMPL_WIDTH),
		25592 => to_signed(20807, LUT_AMPL_WIDTH),
		25593 => to_signed(20804, LUT_AMPL_WIDTH),
		25594 => to_signed(20802, LUT_AMPL_WIDTH),
		25595 => to_signed(20799, LUT_AMPL_WIDTH),
		25596 => to_signed(20797, LUT_AMPL_WIDTH),
		25597 => to_signed(20794, LUT_AMPL_WIDTH),
		25598 => to_signed(20792, LUT_AMPL_WIDTH),
		25599 => to_signed(20790, LUT_AMPL_WIDTH),
		25600 => to_signed(20787, LUT_AMPL_WIDTH),
		25601 => to_signed(20785, LUT_AMPL_WIDTH),
		25602 => to_signed(20782, LUT_AMPL_WIDTH),
		25603 => to_signed(20780, LUT_AMPL_WIDTH),
		25604 => to_signed(20777, LUT_AMPL_WIDTH),
		25605 => to_signed(20775, LUT_AMPL_WIDTH),
		25606 => to_signed(20773, LUT_AMPL_WIDTH),
		25607 => to_signed(20770, LUT_AMPL_WIDTH),
		25608 => to_signed(20768, LUT_AMPL_WIDTH),
		25609 => to_signed(20765, LUT_AMPL_WIDTH),
		25610 => to_signed(20763, LUT_AMPL_WIDTH),
		25611 => to_signed(20760, LUT_AMPL_WIDTH),
		25612 => to_signed(20758, LUT_AMPL_WIDTH),
		25613 => to_signed(20756, LUT_AMPL_WIDTH),
		25614 => to_signed(20753, LUT_AMPL_WIDTH),
		25615 => to_signed(20751, LUT_AMPL_WIDTH),
		25616 => to_signed(20748, LUT_AMPL_WIDTH),
		25617 => to_signed(20746, LUT_AMPL_WIDTH),
		25618 => to_signed(20743, LUT_AMPL_WIDTH),
		25619 => to_signed(20741, LUT_AMPL_WIDTH),
		25620 => to_signed(20739, LUT_AMPL_WIDTH),
		25621 => to_signed(20736, LUT_AMPL_WIDTH),
		25622 => to_signed(20734, LUT_AMPL_WIDTH),
		25623 => to_signed(20731, LUT_AMPL_WIDTH),
		25624 => to_signed(20729, LUT_AMPL_WIDTH),
		25625 => to_signed(20726, LUT_AMPL_WIDTH),
		25626 => to_signed(20724, LUT_AMPL_WIDTH),
		25627 => to_signed(20722, LUT_AMPL_WIDTH),
		25628 => to_signed(20719, LUT_AMPL_WIDTH),
		25629 => to_signed(20717, LUT_AMPL_WIDTH),
		25630 => to_signed(20714, LUT_AMPL_WIDTH),
		25631 => to_signed(20712, LUT_AMPL_WIDTH),
		25632 => to_signed(20709, LUT_AMPL_WIDTH),
		25633 => to_signed(20707, LUT_AMPL_WIDTH),
		25634 => to_signed(20704, LUT_AMPL_WIDTH),
		25635 => to_signed(20702, LUT_AMPL_WIDTH),
		25636 => to_signed(20700, LUT_AMPL_WIDTH),
		25637 => to_signed(20697, LUT_AMPL_WIDTH),
		25638 => to_signed(20695, LUT_AMPL_WIDTH),
		25639 => to_signed(20692, LUT_AMPL_WIDTH),
		25640 => to_signed(20690, LUT_AMPL_WIDTH),
		25641 => to_signed(20687, LUT_AMPL_WIDTH),
		25642 => to_signed(20685, LUT_AMPL_WIDTH),
		25643 => to_signed(20683, LUT_AMPL_WIDTH),
		25644 => to_signed(20680, LUT_AMPL_WIDTH),
		25645 => to_signed(20678, LUT_AMPL_WIDTH),
		25646 => to_signed(20675, LUT_AMPL_WIDTH),
		25647 => to_signed(20673, LUT_AMPL_WIDTH),
		25648 => to_signed(20670, LUT_AMPL_WIDTH),
		25649 => to_signed(20668, LUT_AMPL_WIDTH),
		25650 => to_signed(20666, LUT_AMPL_WIDTH),
		25651 => to_signed(20663, LUT_AMPL_WIDTH),
		25652 => to_signed(20661, LUT_AMPL_WIDTH),
		25653 => to_signed(20658, LUT_AMPL_WIDTH),
		25654 => to_signed(20656, LUT_AMPL_WIDTH),
		25655 => to_signed(20653, LUT_AMPL_WIDTH),
		25656 => to_signed(20651, LUT_AMPL_WIDTH),
		25657 => to_signed(20648, LUT_AMPL_WIDTH),
		25658 => to_signed(20646, LUT_AMPL_WIDTH),
		25659 => to_signed(20644, LUT_AMPL_WIDTH),
		25660 => to_signed(20641, LUT_AMPL_WIDTH),
		25661 => to_signed(20639, LUT_AMPL_WIDTH),
		25662 => to_signed(20636, LUT_AMPL_WIDTH),
		25663 => to_signed(20634, LUT_AMPL_WIDTH),
		25664 => to_signed(20631, LUT_AMPL_WIDTH),
		25665 => to_signed(20629, LUT_AMPL_WIDTH),
		25666 => to_signed(20626, LUT_AMPL_WIDTH),
		25667 => to_signed(20624, LUT_AMPL_WIDTH),
		25668 => to_signed(20622, LUT_AMPL_WIDTH),
		25669 => to_signed(20619, LUT_AMPL_WIDTH),
		25670 => to_signed(20617, LUT_AMPL_WIDTH),
		25671 => to_signed(20614, LUT_AMPL_WIDTH),
		25672 => to_signed(20612, LUT_AMPL_WIDTH),
		25673 => to_signed(20609, LUT_AMPL_WIDTH),
		25674 => to_signed(20607, LUT_AMPL_WIDTH),
		25675 => to_signed(20604, LUT_AMPL_WIDTH),
		25676 => to_signed(20602, LUT_AMPL_WIDTH),
		25677 => to_signed(20600, LUT_AMPL_WIDTH),
		25678 => to_signed(20597, LUT_AMPL_WIDTH),
		25679 => to_signed(20595, LUT_AMPL_WIDTH),
		25680 => to_signed(20592, LUT_AMPL_WIDTH),
		25681 => to_signed(20590, LUT_AMPL_WIDTH),
		25682 => to_signed(20587, LUT_AMPL_WIDTH),
		25683 => to_signed(20585, LUT_AMPL_WIDTH),
		25684 => to_signed(20583, LUT_AMPL_WIDTH),
		25685 => to_signed(20580, LUT_AMPL_WIDTH),
		25686 => to_signed(20578, LUT_AMPL_WIDTH),
		25687 => to_signed(20575, LUT_AMPL_WIDTH),
		25688 => to_signed(20573, LUT_AMPL_WIDTH),
		25689 => to_signed(20570, LUT_AMPL_WIDTH),
		25690 => to_signed(20568, LUT_AMPL_WIDTH),
		25691 => to_signed(20565, LUT_AMPL_WIDTH),
		25692 => to_signed(20563, LUT_AMPL_WIDTH),
		25693 => to_signed(20560, LUT_AMPL_WIDTH),
		25694 => to_signed(20558, LUT_AMPL_WIDTH),
		25695 => to_signed(20556, LUT_AMPL_WIDTH),
		25696 => to_signed(20553, LUT_AMPL_WIDTH),
		25697 => to_signed(20551, LUT_AMPL_WIDTH),
		25698 => to_signed(20548, LUT_AMPL_WIDTH),
		25699 => to_signed(20546, LUT_AMPL_WIDTH),
		25700 => to_signed(20543, LUT_AMPL_WIDTH),
		25701 => to_signed(20541, LUT_AMPL_WIDTH),
		25702 => to_signed(20538, LUT_AMPL_WIDTH),
		25703 => to_signed(20536, LUT_AMPL_WIDTH),
		25704 => to_signed(20534, LUT_AMPL_WIDTH),
		25705 => to_signed(20531, LUT_AMPL_WIDTH),
		25706 => to_signed(20529, LUT_AMPL_WIDTH),
		25707 => to_signed(20526, LUT_AMPL_WIDTH),
		25708 => to_signed(20524, LUT_AMPL_WIDTH),
		25709 => to_signed(20521, LUT_AMPL_WIDTH),
		25710 => to_signed(20519, LUT_AMPL_WIDTH),
		25711 => to_signed(20516, LUT_AMPL_WIDTH),
		25712 => to_signed(20514, LUT_AMPL_WIDTH),
		25713 => to_signed(20512, LUT_AMPL_WIDTH),
		25714 => to_signed(20509, LUT_AMPL_WIDTH),
		25715 => to_signed(20507, LUT_AMPL_WIDTH),
		25716 => to_signed(20504, LUT_AMPL_WIDTH),
		25717 => to_signed(20502, LUT_AMPL_WIDTH),
		25718 => to_signed(20499, LUT_AMPL_WIDTH),
		25719 => to_signed(20497, LUT_AMPL_WIDTH),
		25720 => to_signed(20494, LUT_AMPL_WIDTH),
		25721 => to_signed(20492, LUT_AMPL_WIDTH),
		25722 => to_signed(20489, LUT_AMPL_WIDTH),
		25723 => to_signed(20487, LUT_AMPL_WIDTH),
		25724 => to_signed(20485, LUT_AMPL_WIDTH),
		25725 => to_signed(20482, LUT_AMPL_WIDTH),
		25726 => to_signed(20480, LUT_AMPL_WIDTH),
		25727 => to_signed(20477, LUT_AMPL_WIDTH),
		25728 => to_signed(20475, LUT_AMPL_WIDTH),
		25729 => to_signed(20472, LUT_AMPL_WIDTH),
		25730 => to_signed(20470, LUT_AMPL_WIDTH),
		25731 => to_signed(20467, LUT_AMPL_WIDTH),
		25732 => to_signed(20465, LUT_AMPL_WIDTH),
		25733 => to_signed(20463, LUT_AMPL_WIDTH),
		25734 => to_signed(20460, LUT_AMPL_WIDTH),
		25735 => to_signed(20458, LUT_AMPL_WIDTH),
		25736 => to_signed(20455, LUT_AMPL_WIDTH),
		25737 => to_signed(20453, LUT_AMPL_WIDTH),
		25738 => to_signed(20450, LUT_AMPL_WIDTH),
		25739 => to_signed(20448, LUT_AMPL_WIDTH),
		25740 => to_signed(20445, LUT_AMPL_WIDTH),
		25741 => to_signed(20443, LUT_AMPL_WIDTH),
		25742 => to_signed(20440, LUT_AMPL_WIDTH),
		25743 => to_signed(20438, LUT_AMPL_WIDTH),
		25744 => to_signed(20436, LUT_AMPL_WIDTH),
		25745 => to_signed(20433, LUT_AMPL_WIDTH),
		25746 => to_signed(20431, LUT_AMPL_WIDTH),
		25747 => to_signed(20428, LUT_AMPL_WIDTH),
		25748 => to_signed(20426, LUT_AMPL_WIDTH),
		25749 => to_signed(20423, LUT_AMPL_WIDTH),
		25750 => to_signed(20421, LUT_AMPL_WIDTH),
		25751 => to_signed(20418, LUT_AMPL_WIDTH),
		25752 => to_signed(20416, LUT_AMPL_WIDTH),
		25753 => to_signed(20413, LUT_AMPL_WIDTH),
		25754 => to_signed(20411, LUT_AMPL_WIDTH),
		25755 => to_signed(20408, LUT_AMPL_WIDTH),
		25756 => to_signed(20406, LUT_AMPL_WIDTH),
		25757 => to_signed(20404, LUT_AMPL_WIDTH),
		25758 => to_signed(20401, LUT_AMPL_WIDTH),
		25759 => to_signed(20399, LUT_AMPL_WIDTH),
		25760 => to_signed(20396, LUT_AMPL_WIDTH),
		25761 => to_signed(20394, LUT_AMPL_WIDTH),
		25762 => to_signed(20391, LUT_AMPL_WIDTH),
		25763 => to_signed(20389, LUT_AMPL_WIDTH),
		25764 => to_signed(20386, LUT_AMPL_WIDTH),
		25765 => to_signed(20384, LUT_AMPL_WIDTH),
		25766 => to_signed(20381, LUT_AMPL_WIDTH),
		25767 => to_signed(20379, LUT_AMPL_WIDTH),
		25768 => to_signed(20377, LUT_AMPL_WIDTH),
		25769 => to_signed(20374, LUT_AMPL_WIDTH),
		25770 => to_signed(20372, LUT_AMPL_WIDTH),
		25771 => to_signed(20369, LUT_AMPL_WIDTH),
		25772 => to_signed(20367, LUT_AMPL_WIDTH),
		25773 => to_signed(20364, LUT_AMPL_WIDTH),
		25774 => to_signed(20362, LUT_AMPL_WIDTH),
		25775 => to_signed(20359, LUT_AMPL_WIDTH),
		25776 => to_signed(20357, LUT_AMPL_WIDTH),
		25777 => to_signed(20354, LUT_AMPL_WIDTH),
		25778 => to_signed(20352, LUT_AMPL_WIDTH),
		25779 => to_signed(20349, LUT_AMPL_WIDTH),
		25780 => to_signed(20347, LUT_AMPL_WIDTH),
		25781 => to_signed(20345, LUT_AMPL_WIDTH),
		25782 => to_signed(20342, LUT_AMPL_WIDTH),
		25783 => to_signed(20340, LUT_AMPL_WIDTH),
		25784 => to_signed(20337, LUT_AMPL_WIDTH),
		25785 => to_signed(20335, LUT_AMPL_WIDTH),
		25786 => to_signed(20332, LUT_AMPL_WIDTH),
		25787 => to_signed(20330, LUT_AMPL_WIDTH),
		25788 => to_signed(20327, LUT_AMPL_WIDTH),
		25789 => to_signed(20325, LUT_AMPL_WIDTH),
		25790 => to_signed(20322, LUT_AMPL_WIDTH),
		25791 => to_signed(20320, LUT_AMPL_WIDTH),
		25792 => to_signed(20317, LUT_AMPL_WIDTH),
		25793 => to_signed(20315, LUT_AMPL_WIDTH),
		25794 => to_signed(20312, LUT_AMPL_WIDTH),
		25795 => to_signed(20310, LUT_AMPL_WIDTH),
		25796 => to_signed(20308, LUT_AMPL_WIDTH),
		25797 => to_signed(20305, LUT_AMPL_WIDTH),
		25798 => to_signed(20303, LUT_AMPL_WIDTH),
		25799 => to_signed(20300, LUT_AMPL_WIDTH),
		25800 => to_signed(20298, LUT_AMPL_WIDTH),
		25801 => to_signed(20295, LUT_AMPL_WIDTH),
		25802 => to_signed(20293, LUT_AMPL_WIDTH),
		25803 => to_signed(20290, LUT_AMPL_WIDTH),
		25804 => to_signed(20288, LUT_AMPL_WIDTH),
		25805 => to_signed(20285, LUT_AMPL_WIDTH),
		25806 => to_signed(20283, LUT_AMPL_WIDTH),
		25807 => to_signed(20280, LUT_AMPL_WIDTH),
		25808 => to_signed(20278, LUT_AMPL_WIDTH),
		25809 => to_signed(20275, LUT_AMPL_WIDTH),
		25810 => to_signed(20273, LUT_AMPL_WIDTH),
		25811 => to_signed(20271, LUT_AMPL_WIDTH),
		25812 => to_signed(20268, LUT_AMPL_WIDTH),
		25813 => to_signed(20266, LUT_AMPL_WIDTH),
		25814 => to_signed(20263, LUT_AMPL_WIDTH),
		25815 => to_signed(20261, LUT_AMPL_WIDTH),
		25816 => to_signed(20258, LUT_AMPL_WIDTH),
		25817 => to_signed(20256, LUT_AMPL_WIDTH),
		25818 => to_signed(20253, LUT_AMPL_WIDTH),
		25819 => to_signed(20251, LUT_AMPL_WIDTH),
		25820 => to_signed(20248, LUT_AMPL_WIDTH),
		25821 => to_signed(20246, LUT_AMPL_WIDTH),
		25822 => to_signed(20243, LUT_AMPL_WIDTH),
		25823 => to_signed(20241, LUT_AMPL_WIDTH),
		25824 => to_signed(20238, LUT_AMPL_WIDTH),
		25825 => to_signed(20236, LUT_AMPL_WIDTH),
		25826 => to_signed(20234, LUT_AMPL_WIDTH),
		25827 => to_signed(20231, LUT_AMPL_WIDTH),
		25828 => to_signed(20229, LUT_AMPL_WIDTH),
		25829 => to_signed(20226, LUT_AMPL_WIDTH),
		25830 => to_signed(20224, LUT_AMPL_WIDTH),
		25831 => to_signed(20221, LUT_AMPL_WIDTH),
		25832 => to_signed(20219, LUT_AMPL_WIDTH),
		25833 => to_signed(20216, LUT_AMPL_WIDTH),
		25834 => to_signed(20214, LUT_AMPL_WIDTH),
		25835 => to_signed(20211, LUT_AMPL_WIDTH),
		25836 => to_signed(20209, LUT_AMPL_WIDTH),
		25837 => to_signed(20206, LUT_AMPL_WIDTH),
		25838 => to_signed(20204, LUT_AMPL_WIDTH),
		25839 => to_signed(20201, LUT_AMPL_WIDTH),
		25840 => to_signed(20199, LUT_AMPL_WIDTH),
		25841 => to_signed(20196, LUT_AMPL_WIDTH),
		25842 => to_signed(20194, LUT_AMPL_WIDTH),
		25843 => to_signed(20191, LUT_AMPL_WIDTH),
		25844 => to_signed(20189, LUT_AMPL_WIDTH),
		25845 => to_signed(20187, LUT_AMPL_WIDTH),
		25846 => to_signed(20184, LUT_AMPL_WIDTH),
		25847 => to_signed(20182, LUT_AMPL_WIDTH),
		25848 => to_signed(20179, LUT_AMPL_WIDTH),
		25849 => to_signed(20177, LUT_AMPL_WIDTH),
		25850 => to_signed(20174, LUT_AMPL_WIDTH),
		25851 => to_signed(20172, LUT_AMPL_WIDTH),
		25852 => to_signed(20169, LUT_AMPL_WIDTH),
		25853 => to_signed(20167, LUT_AMPL_WIDTH),
		25854 => to_signed(20164, LUT_AMPL_WIDTH),
		25855 => to_signed(20162, LUT_AMPL_WIDTH),
		25856 => to_signed(20159, LUT_AMPL_WIDTH),
		25857 => to_signed(20157, LUT_AMPL_WIDTH),
		25858 => to_signed(20154, LUT_AMPL_WIDTH),
		25859 => to_signed(20152, LUT_AMPL_WIDTH),
		25860 => to_signed(20149, LUT_AMPL_WIDTH),
		25861 => to_signed(20147, LUT_AMPL_WIDTH),
		25862 => to_signed(20144, LUT_AMPL_WIDTH),
		25863 => to_signed(20142, LUT_AMPL_WIDTH),
		25864 => to_signed(20139, LUT_AMPL_WIDTH),
		25865 => to_signed(20137, LUT_AMPL_WIDTH),
		25866 => to_signed(20135, LUT_AMPL_WIDTH),
		25867 => to_signed(20132, LUT_AMPL_WIDTH),
		25868 => to_signed(20130, LUT_AMPL_WIDTH),
		25869 => to_signed(20127, LUT_AMPL_WIDTH),
		25870 => to_signed(20125, LUT_AMPL_WIDTH),
		25871 => to_signed(20122, LUT_AMPL_WIDTH),
		25872 => to_signed(20120, LUT_AMPL_WIDTH),
		25873 => to_signed(20117, LUT_AMPL_WIDTH),
		25874 => to_signed(20115, LUT_AMPL_WIDTH),
		25875 => to_signed(20112, LUT_AMPL_WIDTH),
		25876 => to_signed(20110, LUT_AMPL_WIDTH),
		25877 => to_signed(20107, LUT_AMPL_WIDTH),
		25878 => to_signed(20105, LUT_AMPL_WIDTH),
		25879 => to_signed(20102, LUT_AMPL_WIDTH),
		25880 => to_signed(20100, LUT_AMPL_WIDTH),
		25881 => to_signed(20097, LUT_AMPL_WIDTH),
		25882 => to_signed(20095, LUT_AMPL_WIDTH),
		25883 => to_signed(20092, LUT_AMPL_WIDTH),
		25884 => to_signed(20090, LUT_AMPL_WIDTH),
		25885 => to_signed(20087, LUT_AMPL_WIDTH),
		25886 => to_signed(20085, LUT_AMPL_WIDTH),
		25887 => to_signed(20082, LUT_AMPL_WIDTH),
		25888 => to_signed(20080, LUT_AMPL_WIDTH),
		25889 => to_signed(20077, LUT_AMPL_WIDTH),
		25890 => to_signed(20075, LUT_AMPL_WIDTH),
		25891 => to_signed(20072, LUT_AMPL_WIDTH),
		25892 => to_signed(20070, LUT_AMPL_WIDTH),
		25893 => to_signed(20068, LUT_AMPL_WIDTH),
		25894 => to_signed(20065, LUT_AMPL_WIDTH),
		25895 => to_signed(20063, LUT_AMPL_WIDTH),
		25896 => to_signed(20060, LUT_AMPL_WIDTH),
		25897 => to_signed(20058, LUT_AMPL_WIDTH),
		25898 => to_signed(20055, LUT_AMPL_WIDTH),
		25899 => to_signed(20053, LUT_AMPL_WIDTH),
		25900 => to_signed(20050, LUT_AMPL_WIDTH),
		25901 => to_signed(20048, LUT_AMPL_WIDTH),
		25902 => to_signed(20045, LUT_AMPL_WIDTH),
		25903 => to_signed(20043, LUT_AMPL_WIDTH),
		25904 => to_signed(20040, LUT_AMPL_WIDTH),
		25905 => to_signed(20038, LUT_AMPL_WIDTH),
		25906 => to_signed(20035, LUT_AMPL_WIDTH),
		25907 => to_signed(20033, LUT_AMPL_WIDTH),
		25908 => to_signed(20030, LUT_AMPL_WIDTH),
		25909 => to_signed(20028, LUT_AMPL_WIDTH),
		25910 => to_signed(20025, LUT_AMPL_WIDTH),
		25911 => to_signed(20023, LUT_AMPL_WIDTH),
		25912 => to_signed(20020, LUT_AMPL_WIDTH),
		25913 => to_signed(20018, LUT_AMPL_WIDTH),
		25914 => to_signed(20015, LUT_AMPL_WIDTH),
		25915 => to_signed(20013, LUT_AMPL_WIDTH),
		25916 => to_signed(20010, LUT_AMPL_WIDTH),
		25917 => to_signed(20008, LUT_AMPL_WIDTH),
		25918 => to_signed(20005, LUT_AMPL_WIDTH),
		25919 => to_signed(20003, LUT_AMPL_WIDTH),
		25920 => to_signed(20000, LUT_AMPL_WIDTH),
		25921 => to_signed(19998, LUT_AMPL_WIDTH),
		25922 => to_signed(19995, LUT_AMPL_WIDTH),
		25923 => to_signed(19993, LUT_AMPL_WIDTH),
		25924 => to_signed(19990, LUT_AMPL_WIDTH),
		25925 => to_signed(19988, LUT_AMPL_WIDTH),
		25926 => to_signed(19985, LUT_AMPL_WIDTH),
		25927 => to_signed(19983, LUT_AMPL_WIDTH),
		25928 => to_signed(19981, LUT_AMPL_WIDTH),
		25929 => to_signed(19978, LUT_AMPL_WIDTH),
		25930 => to_signed(19976, LUT_AMPL_WIDTH),
		25931 => to_signed(19973, LUT_AMPL_WIDTH),
		25932 => to_signed(19971, LUT_AMPL_WIDTH),
		25933 => to_signed(19968, LUT_AMPL_WIDTH),
		25934 => to_signed(19966, LUT_AMPL_WIDTH),
		25935 => to_signed(19963, LUT_AMPL_WIDTH),
		25936 => to_signed(19961, LUT_AMPL_WIDTH),
		25937 => to_signed(19958, LUT_AMPL_WIDTH),
		25938 => to_signed(19956, LUT_AMPL_WIDTH),
		25939 => to_signed(19953, LUT_AMPL_WIDTH),
		25940 => to_signed(19951, LUT_AMPL_WIDTH),
		25941 => to_signed(19948, LUT_AMPL_WIDTH),
		25942 => to_signed(19946, LUT_AMPL_WIDTH),
		25943 => to_signed(19943, LUT_AMPL_WIDTH),
		25944 => to_signed(19941, LUT_AMPL_WIDTH),
		25945 => to_signed(19938, LUT_AMPL_WIDTH),
		25946 => to_signed(19936, LUT_AMPL_WIDTH),
		25947 => to_signed(19933, LUT_AMPL_WIDTH),
		25948 => to_signed(19931, LUT_AMPL_WIDTH),
		25949 => to_signed(19928, LUT_AMPL_WIDTH),
		25950 => to_signed(19926, LUT_AMPL_WIDTH),
		25951 => to_signed(19923, LUT_AMPL_WIDTH),
		25952 => to_signed(19921, LUT_AMPL_WIDTH),
		25953 => to_signed(19918, LUT_AMPL_WIDTH),
		25954 => to_signed(19916, LUT_AMPL_WIDTH),
		25955 => to_signed(19913, LUT_AMPL_WIDTH),
		25956 => to_signed(19911, LUT_AMPL_WIDTH),
		25957 => to_signed(19908, LUT_AMPL_WIDTH),
		25958 => to_signed(19906, LUT_AMPL_WIDTH),
		25959 => to_signed(19903, LUT_AMPL_WIDTH),
		25960 => to_signed(19901, LUT_AMPL_WIDTH),
		25961 => to_signed(19898, LUT_AMPL_WIDTH),
		25962 => to_signed(19896, LUT_AMPL_WIDTH),
		25963 => to_signed(19893, LUT_AMPL_WIDTH),
		25964 => to_signed(19891, LUT_AMPL_WIDTH),
		25965 => to_signed(19888, LUT_AMPL_WIDTH),
		25966 => to_signed(19886, LUT_AMPL_WIDTH),
		25967 => to_signed(19883, LUT_AMPL_WIDTH),
		25968 => to_signed(19881, LUT_AMPL_WIDTH),
		25969 => to_signed(19878, LUT_AMPL_WIDTH),
		25970 => to_signed(19876, LUT_AMPL_WIDTH),
		25971 => to_signed(19873, LUT_AMPL_WIDTH),
		25972 => to_signed(19871, LUT_AMPL_WIDTH),
		25973 => to_signed(19868, LUT_AMPL_WIDTH),
		25974 => to_signed(19866, LUT_AMPL_WIDTH),
		25975 => to_signed(19863, LUT_AMPL_WIDTH),
		25976 => to_signed(19861, LUT_AMPL_WIDTH),
		25977 => to_signed(19858, LUT_AMPL_WIDTH),
		25978 => to_signed(19856, LUT_AMPL_WIDTH),
		25979 => to_signed(19853, LUT_AMPL_WIDTH),
		25980 => to_signed(19851, LUT_AMPL_WIDTH),
		25981 => to_signed(19848, LUT_AMPL_WIDTH),
		25982 => to_signed(19846, LUT_AMPL_WIDTH),
		25983 => to_signed(19843, LUT_AMPL_WIDTH),
		25984 => to_signed(19841, LUT_AMPL_WIDTH),
		25985 => to_signed(19838, LUT_AMPL_WIDTH),
		25986 => to_signed(19836, LUT_AMPL_WIDTH),
		25987 => to_signed(19833, LUT_AMPL_WIDTH),
		25988 => to_signed(19831, LUT_AMPL_WIDTH),
		25989 => to_signed(19828, LUT_AMPL_WIDTH),
		25990 => to_signed(19826, LUT_AMPL_WIDTH),
		25991 => to_signed(19823, LUT_AMPL_WIDTH),
		25992 => to_signed(19821, LUT_AMPL_WIDTH),
		25993 => to_signed(19818, LUT_AMPL_WIDTH),
		25994 => to_signed(19816, LUT_AMPL_WIDTH),
		25995 => to_signed(19813, LUT_AMPL_WIDTH),
		25996 => to_signed(19811, LUT_AMPL_WIDTH),
		25997 => to_signed(19808, LUT_AMPL_WIDTH),
		25998 => to_signed(19806, LUT_AMPL_WIDTH),
		25999 => to_signed(19803, LUT_AMPL_WIDTH),
		26000 => to_signed(19801, LUT_AMPL_WIDTH),
		26001 => to_signed(19798, LUT_AMPL_WIDTH),
		26002 => to_signed(19796, LUT_AMPL_WIDTH),
		26003 => to_signed(19793, LUT_AMPL_WIDTH),
		26004 => to_signed(19791, LUT_AMPL_WIDTH),
		26005 => to_signed(19788, LUT_AMPL_WIDTH),
		26006 => to_signed(19786, LUT_AMPL_WIDTH),
		26007 => to_signed(19783, LUT_AMPL_WIDTH),
		26008 => to_signed(19781, LUT_AMPL_WIDTH),
		26009 => to_signed(19778, LUT_AMPL_WIDTH),
		26010 => to_signed(19776, LUT_AMPL_WIDTH),
		26011 => to_signed(19773, LUT_AMPL_WIDTH),
		26012 => to_signed(19771, LUT_AMPL_WIDTH),
		26013 => to_signed(19768, LUT_AMPL_WIDTH),
		26014 => to_signed(19766, LUT_AMPL_WIDTH),
		26015 => to_signed(19763, LUT_AMPL_WIDTH),
		26016 => to_signed(19761, LUT_AMPL_WIDTH),
		26017 => to_signed(19758, LUT_AMPL_WIDTH),
		26018 => to_signed(19756, LUT_AMPL_WIDTH),
		26019 => to_signed(19753, LUT_AMPL_WIDTH),
		26020 => to_signed(19751, LUT_AMPL_WIDTH),
		26021 => to_signed(19748, LUT_AMPL_WIDTH),
		26022 => to_signed(19746, LUT_AMPL_WIDTH),
		26023 => to_signed(19743, LUT_AMPL_WIDTH),
		26024 => to_signed(19741, LUT_AMPL_WIDTH),
		26025 => to_signed(19738, LUT_AMPL_WIDTH),
		26026 => to_signed(19736, LUT_AMPL_WIDTH),
		26027 => to_signed(19733, LUT_AMPL_WIDTH),
		26028 => to_signed(19731, LUT_AMPL_WIDTH),
		26029 => to_signed(19728, LUT_AMPL_WIDTH),
		26030 => to_signed(19726, LUT_AMPL_WIDTH),
		26031 => to_signed(19723, LUT_AMPL_WIDTH),
		26032 => to_signed(19721, LUT_AMPL_WIDTH),
		26033 => to_signed(19718, LUT_AMPL_WIDTH),
		26034 => to_signed(19716, LUT_AMPL_WIDTH),
		26035 => to_signed(19713, LUT_AMPL_WIDTH),
		26036 => to_signed(19711, LUT_AMPL_WIDTH),
		26037 => to_signed(19708, LUT_AMPL_WIDTH),
		26038 => to_signed(19706, LUT_AMPL_WIDTH),
		26039 => to_signed(19703, LUT_AMPL_WIDTH),
		26040 => to_signed(19700, LUT_AMPL_WIDTH),
		26041 => to_signed(19698, LUT_AMPL_WIDTH),
		26042 => to_signed(19695, LUT_AMPL_WIDTH),
		26043 => to_signed(19693, LUT_AMPL_WIDTH),
		26044 => to_signed(19690, LUT_AMPL_WIDTH),
		26045 => to_signed(19688, LUT_AMPL_WIDTH),
		26046 => to_signed(19685, LUT_AMPL_WIDTH),
		26047 => to_signed(19683, LUT_AMPL_WIDTH),
		26048 => to_signed(19680, LUT_AMPL_WIDTH),
		26049 => to_signed(19678, LUT_AMPL_WIDTH),
		26050 => to_signed(19675, LUT_AMPL_WIDTH),
		26051 => to_signed(19673, LUT_AMPL_WIDTH),
		26052 => to_signed(19670, LUT_AMPL_WIDTH),
		26053 => to_signed(19668, LUT_AMPL_WIDTH),
		26054 => to_signed(19665, LUT_AMPL_WIDTH),
		26055 => to_signed(19663, LUT_AMPL_WIDTH),
		26056 => to_signed(19660, LUT_AMPL_WIDTH),
		26057 => to_signed(19658, LUT_AMPL_WIDTH),
		26058 => to_signed(19655, LUT_AMPL_WIDTH),
		26059 => to_signed(19653, LUT_AMPL_WIDTH),
		26060 => to_signed(19650, LUT_AMPL_WIDTH),
		26061 => to_signed(19648, LUT_AMPL_WIDTH),
		26062 => to_signed(19645, LUT_AMPL_WIDTH),
		26063 => to_signed(19643, LUT_AMPL_WIDTH),
		26064 => to_signed(19640, LUT_AMPL_WIDTH),
		26065 => to_signed(19638, LUT_AMPL_WIDTH),
		26066 => to_signed(19635, LUT_AMPL_WIDTH),
		26067 => to_signed(19633, LUT_AMPL_WIDTH),
		26068 => to_signed(19630, LUT_AMPL_WIDTH),
		26069 => to_signed(19628, LUT_AMPL_WIDTH),
		26070 => to_signed(19625, LUT_AMPL_WIDTH),
		26071 => to_signed(19623, LUT_AMPL_WIDTH),
		26072 => to_signed(19620, LUT_AMPL_WIDTH),
		26073 => to_signed(19618, LUT_AMPL_WIDTH),
		26074 => to_signed(19615, LUT_AMPL_WIDTH),
		26075 => to_signed(19613, LUT_AMPL_WIDTH),
		26076 => to_signed(19610, LUT_AMPL_WIDTH),
		26077 => to_signed(19607, LUT_AMPL_WIDTH),
		26078 => to_signed(19605, LUT_AMPL_WIDTH),
		26079 => to_signed(19602, LUT_AMPL_WIDTH),
		26080 => to_signed(19600, LUT_AMPL_WIDTH),
		26081 => to_signed(19597, LUT_AMPL_WIDTH),
		26082 => to_signed(19595, LUT_AMPL_WIDTH),
		26083 => to_signed(19592, LUT_AMPL_WIDTH),
		26084 => to_signed(19590, LUT_AMPL_WIDTH),
		26085 => to_signed(19587, LUT_AMPL_WIDTH),
		26086 => to_signed(19585, LUT_AMPL_WIDTH),
		26087 => to_signed(19582, LUT_AMPL_WIDTH),
		26088 => to_signed(19580, LUT_AMPL_WIDTH),
		26089 => to_signed(19577, LUT_AMPL_WIDTH),
		26090 => to_signed(19575, LUT_AMPL_WIDTH),
		26091 => to_signed(19572, LUT_AMPL_WIDTH),
		26092 => to_signed(19570, LUT_AMPL_WIDTH),
		26093 => to_signed(19567, LUT_AMPL_WIDTH),
		26094 => to_signed(19565, LUT_AMPL_WIDTH),
		26095 => to_signed(19562, LUT_AMPL_WIDTH),
		26096 => to_signed(19560, LUT_AMPL_WIDTH),
		26097 => to_signed(19557, LUT_AMPL_WIDTH),
		26098 => to_signed(19555, LUT_AMPL_WIDTH),
		26099 => to_signed(19552, LUT_AMPL_WIDTH),
		26100 => to_signed(19550, LUT_AMPL_WIDTH),
		26101 => to_signed(19547, LUT_AMPL_WIDTH),
		26102 => to_signed(19545, LUT_AMPL_WIDTH),
		26103 => to_signed(19542, LUT_AMPL_WIDTH),
		26104 => to_signed(19539, LUT_AMPL_WIDTH),
		26105 => to_signed(19537, LUT_AMPL_WIDTH),
		26106 => to_signed(19534, LUT_AMPL_WIDTH),
		26107 => to_signed(19532, LUT_AMPL_WIDTH),
		26108 => to_signed(19529, LUT_AMPL_WIDTH),
		26109 => to_signed(19527, LUT_AMPL_WIDTH),
		26110 => to_signed(19524, LUT_AMPL_WIDTH),
		26111 => to_signed(19522, LUT_AMPL_WIDTH),
		26112 => to_signed(19519, LUT_AMPL_WIDTH),
		26113 => to_signed(19517, LUT_AMPL_WIDTH),
		26114 => to_signed(19514, LUT_AMPL_WIDTH),
		26115 => to_signed(19512, LUT_AMPL_WIDTH),
		26116 => to_signed(19509, LUT_AMPL_WIDTH),
		26117 => to_signed(19507, LUT_AMPL_WIDTH),
		26118 => to_signed(19504, LUT_AMPL_WIDTH),
		26119 => to_signed(19502, LUT_AMPL_WIDTH),
		26120 => to_signed(19499, LUT_AMPL_WIDTH),
		26121 => to_signed(19497, LUT_AMPL_WIDTH),
		26122 => to_signed(19494, LUT_AMPL_WIDTH),
		26123 => to_signed(19492, LUT_AMPL_WIDTH),
		26124 => to_signed(19489, LUT_AMPL_WIDTH),
		26125 => to_signed(19486, LUT_AMPL_WIDTH),
		26126 => to_signed(19484, LUT_AMPL_WIDTH),
		26127 => to_signed(19481, LUT_AMPL_WIDTH),
		26128 => to_signed(19479, LUT_AMPL_WIDTH),
		26129 => to_signed(19476, LUT_AMPL_WIDTH),
		26130 => to_signed(19474, LUT_AMPL_WIDTH),
		26131 => to_signed(19471, LUT_AMPL_WIDTH),
		26132 => to_signed(19469, LUT_AMPL_WIDTH),
		26133 => to_signed(19466, LUT_AMPL_WIDTH),
		26134 => to_signed(19464, LUT_AMPL_WIDTH),
		26135 => to_signed(19461, LUT_AMPL_WIDTH),
		26136 => to_signed(19459, LUT_AMPL_WIDTH),
		26137 => to_signed(19456, LUT_AMPL_WIDTH),
		26138 => to_signed(19454, LUT_AMPL_WIDTH),
		26139 => to_signed(19451, LUT_AMPL_WIDTH),
		26140 => to_signed(19449, LUT_AMPL_WIDTH),
		26141 => to_signed(19446, LUT_AMPL_WIDTH),
		26142 => to_signed(19444, LUT_AMPL_WIDTH),
		26143 => to_signed(19441, LUT_AMPL_WIDTH),
		26144 => to_signed(19438, LUT_AMPL_WIDTH),
		26145 => to_signed(19436, LUT_AMPL_WIDTH),
		26146 => to_signed(19433, LUT_AMPL_WIDTH),
		26147 => to_signed(19431, LUT_AMPL_WIDTH),
		26148 => to_signed(19428, LUT_AMPL_WIDTH),
		26149 => to_signed(19426, LUT_AMPL_WIDTH),
		26150 => to_signed(19423, LUT_AMPL_WIDTH),
		26151 => to_signed(19421, LUT_AMPL_WIDTH),
		26152 => to_signed(19418, LUT_AMPL_WIDTH),
		26153 => to_signed(19416, LUT_AMPL_WIDTH),
		26154 => to_signed(19413, LUT_AMPL_WIDTH),
		26155 => to_signed(19411, LUT_AMPL_WIDTH),
		26156 => to_signed(19408, LUT_AMPL_WIDTH),
		26157 => to_signed(19406, LUT_AMPL_WIDTH),
		26158 => to_signed(19403, LUT_AMPL_WIDTH),
		26159 => to_signed(19400, LUT_AMPL_WIDTH),
		26160 => to_signed(19398, LUT_AMPL_WIDTH),
		26161 => to_signed(19395, LUT_AMPL_WIDTH),
		26162 => to_signed(19393, LUT_AMPL_WIDTH),
		26163 => to_signed(19390, LUT_AMPL_WIDTH),
		26164 => to_signed(19388, LUT_AMPL_WIDTH),
		26165 => to_signed(19385, LUT_AMPL_WIDTH),
		26166 => to_signed(19383, LUT_AMPL_WIDTH),
		26167 => to_signed(19380, LUT_AMPL_WIDTH),
		26168 => to_signed(19378, LUT_AMPL_WIDTH),
		26169 => to_signed(19375, LUT_AMPL_WIDTH),
		26170 => to_signed(19373, LUT_AMPL_WIDTH),
		26171 => to_signed(19370, LUT_AMPL_WIDTH),
		26172 => to_signed(19368, LUT_AMPL_WIDTH),
		26173 => to_signed(19365, LUT_AMPL_WIDTH),
		26174 => to_signed(19362, LUT_AMPL_WIDTH),
		26175 => to_signed(19360, LUT_AMPL_WIDTH),
		26176 => to_signed(19357, LUT_AMPL_WIDTH),
		26177 => to_signed(19355, LUT_AMPL_WIDTH),
		26178 => to_signed(19352, LUT_AMPL_WIDTH),
		26179 => to_signed(19350, LUT_AMPL_WIDTH),
		26180 => to_signed(19347, LUT_AMPL_WIDTH),
		26181 => to_signed(19345, LUT_AMPL_WIDTH),
		26182 => to_signed(19342, LUT_AMPL_WIDTH),
		26183 => to_signed(19340, LUT_AMPL_WIDTH),
		26184 => to_signed(19337, LUT_AMPL_WIDTH),
		26185 => to_signed(19335, LUT_AMPL_WIDTH),
		26186 => to_signed(19332, LUT_AMPL_WIDTH),
		26187 => to_signed(19330, LUT_AMPL_WIDTH),
		26188 => to_signed(19327, LUT_AMPL_WIDTH),
		26189 => to_signed(19324, LUT_AMPL_WIDTH),
		26190 => to_signed(19322, LUT_AMPL_WIDTH),
		26191 => to_signed(19319, LUT_AMPL_WIDTH),
		26192 => to_signed(19317, LUT_AMPL_WIDTH),
		26193 => to_signed(19314, LUT_AMPL_WIDTH),
		26194 => to_signed(19312, LUT_AMPL_WIDTH),
		26195 => to_signed(19309, LUT_AMPL_WIDTH),
		26196 => to_signed(19307, LUT_AMPL_WIDTH),
		26197 => to_signed(19304, LUT_AMPL_WIDTH),
		26198 => to_signed(19302, LUT_AMPL_WIDTH),
		26199 => to_signed(19299, LUT_AMPL_WIDTH),
		26200 => to_signed(19297, LUT_AMPL_WIDTH),
		26201 => to_signed(19294, LUT_AMPL_WIDTH),
		26202 => to_signed(19291, LUT_AMPL_WIDTH),
		26203 => to_signed(19289, LUT_AMPL_WIDTH),
		26204 => to_signed(19286, LUT_AMPL_WIDTH),
		26205 => to_signed(19284, LUT_AMPL_WIDTH),
		26206 => to_signed(19281, LUT_AMPL_WIDTH),
		26207 => to_signed(19279, LUT_AMPL_WIDTH),
		26208 => to_signed(19276, LUT_AMPL_WIDTH),
		26209 => to_signed(19274, LUT_AMPL_WIDTH),
		26210 => to_signed(19271, LUT_AMPL_WIDTH),
		26211 => to_signed(19269, LUT_AMPL_WIDTH),
		26212 => to_signed(19266, LUT_AMPL_WIDTH),
		26213 => to_signed(19264, LUT_AMPL_WIDTH),
		26214 => to_signed(19261, LUT_AMPL_WIDTH),
		26215 => to_signed(19258, LUT_AMPL_WIDTH),
		26216 => to_signed(19256, LUT_AMPL_WIDTH),
		26217 => to_signed(19253, LUT_AMPL_WIDTH),
		26218 => to_signed(19251, LUT_AMPL_WIDTH),
		26219 => to_signed(19248, LUT_AMPL_WIDTH),
		26220 => to_signed(19246, LUT_AMPL_WIDTH),
		26221 => to_signed(19243, LUT_AMPL_WIDTH),
		26222 => to_signed(19241, LUT_AMPL_WIDTH),
		26223 => to_signed(19238, LUT_AMPL_WIDTH),
		26224 => to_signed(19236, LUT_AMPL_WIDTH),
		26225 => to_signed(19233, LUT_AMPL_WIDTH),
		26226 => to_signed(19230, LUT_AMPL_WIDTH),
		26227 => to_signed(19228, LUT_AMPL_WIDTH),
		26228 => to_signed(19225, LUT_AMPL_WIDTH),
		26229 => to_signed(19223, LUT_AMPL_WIDTH),
		26230 => to_signed(19220, LUT_AMPL_WIDTH),
		26231 => to_signed(19218, LUT_AMPL_WIDTH),
		26232 => to_signed(19215, LUT_AMPL_WIDTH),
		26233 => to_signed(19213, LUT_AMPL_WIDTH),
		26234 => to_signed(19210, LUT_AMPL_WIDTH),
		26235 => to_signed(19208, LUT_AMPL_WIDTH),
		26236 => to_signed(19205, LUT_AMPL_WIDTH),
		26237 => to_signed(19202, LUT_AMPL_WIDTH),
		26238 => to_signed(19200, LUT_AMPL_WIDTH),
		26239 => to_signed(19197, LUT_AMPL_WIDTH),
		26240 => to_signed(19195, LUT_AMPL_WIDTH),
		26241 => to_signed(19192, LUT_AMPL_WIDTH),
		26242 => to_signed(19190, LUT_AMPL_WIDTH),
		26243 => to_signed(19187, LUT_AMPL_WIDTH),
		26244 => to_signed(19185, LUT_AMPL_WIDTH),
		26245 => to_signed(19182, LUT_AMPL_WIDTH),
		26246 => to_signed(19180, LUT_AMPL_WIDTH),
		26247 => to_signed(19177, LUT_AMPL_WIDTH),
		26248 => to_signed(19174, LUT_AMPL_WIDTH),
		26249 => to_signed(19172, LUT_AMPL_WIDTH),
		26250 => to_signed(19169, LUT_AMPL_WIDTH),
		26251 => to_signed(19167, LUT_AMPL_WIDTH),
		26252 => to_signed(19164, LUT_AMPL_WIDTH),
		26253 => to_signed(19162, LUT_AMPL_WIDTH),
		26254 => to_signed(19159, LUT_AMPL_WIDTH),
		26255 => to_signed(19157, LUT_AMPL_WIDTH),
		26256 => to_signed(19154, LUT_AMPL_WIDTH),
		26257 => to_signed(19152, LUT_AMPL_WIDTH),
		26258 => to_signed(19149, LUT_AMPL_WIDTH),
		26259 => to_signed(19146, LUT_AMPL_WIDTH),
		26260 => to_signed(19144, LUT_AMPL_WIDTH),
		26261 => to_signed(19141, LUT_AMPL_WIDTH),
		26262 => to_signed(19139, LUT_AMPL_WIDTH),
		26263 => to_signed(19136, LUT_AMPL_WIDTH),
		26264 => to_signed(19134, LUT_AMPL_WIDTH),
		26265 => to_signed(19131, LUT_AMPL_WIDTH),
		26266 => to_signed(19129, LUT_AMPL_WIDTH),
		26267 => to_signed(19126, LUT_AMPL_WIDTH),
		26268 => to_signed(19123, LUT_AMPL_WIDTH),
		26269 => to_signed(19121, LUT_AMPL_WIDTH),
		26270 => to_signed(19118, LUT_AMPL_WIDTH),
		26271 => to_signed(19116, LUT_AMPL_WIDTH),
		26272 => to_signed(19113, LUT_AMPL_WIDTH),
		26273 => to_signed(19111, LUT_AMPL_WIDTH),
		26274 => to_signed(19108, LUT_AMPL_WIDTH),
		26275 => to_signed(19106, LUT_AMPL_WIDTH),
		26276 => to_signed(19103, LUT_AMPL_WIDTH),
		26277 => to_signed(19101, LUT_AMPL_WIDTH),
		26278 => to_signed(19098, LUT_AMPL_WIDTH),
		26279 => to_signed(19095, LUT_AMPL_WIDTH),
		26280 => to_signed(19093, LUT_AMPL_WIDTH),
		26281 => to_signed(19090, LUT_AMPL_WIDTH),
		26282 => to_signed(19088, LUT_AMPL_WIDTH),
		26283 => to_signed(19085, LUT_AMPL_WIDTH),
		26284 => to_signed(19083, LUT_AMPL_WIDTH),
		26285 => to_signed(19080, LUT_AMPL_WIDTH),
		26286 => to_signed(19078, LUT_AMPL_WIDTH),
		26287 => to_signed(19075, LUT_AMPL_WIDTH),
		26288 => to_signed(19072, LUT_AMPL_WIDTH),
		26289 => to_signed(19070, LUT_AMPL_WIDTH),
		26290 => to_signed(19067, LUT_AMPL_WIDTH),
		26291 => to_signed(19065, LUT_AMPL_WIDTH),
		26292 => to_signed(19062, LUT_AMPL_WIDTH),
		26293 => to_signed(19060, LUT_AMPL_WIDTH),
		26294 => to_signed(19057, LUT_AMPL_WIDTH),
		26295 => to_signed(19055, LUT_AMPL_WIDTH),
		26296 => to_signed(19052, LUT_AMPL_WIDTH),
		26297 => to_signed(19049, LUT_AMPL_WIDTH),
		26298 => to_signed(19047, LUT_AMPL_WIDTH),
		26299 => to_signed(19044, LUT_AMPL_WIDTH),
		26300 => to_signed(19042, LUT_AMPL_WIDTH),
		26301 => to_signed(19039, LUT_AMPL_WIDTH),
		26302 => to_signed(19037, LUT_AMPL_WIDTH),
		26303 => to_signed(19034, LUT_AMPL_WIDTH),
		26304 => to_signed(19032, LUT_AMPL_WIDTH),
		26305 => to_signed(19029, LUT_AMPL_WIDTH),
		26306 => to_signed(19026, LUT_AMPL_WIDTH),
		26307 => to_signed(19024, LUT_AMPL_WIDTH),
		26308 => to_signed(19021, LUT_AMPL_WIDTH),
		26309 => to_signed(19019, LUT_AMPL_WIDTH),
		26310 => to_signed(19016, LUT_AMPL_WIDTH),
		26311 => to_signed(19014, LUT_AMPL_WIDTH),
		26312 => to_signed(19011, LUT_AMPL_WIDTH),
		26313 => to_signed(19009, LUT_AMPL_WIDTH),
		26314 => to_signed(19006, LUT_AMPL_WIDTH),
		26315 => to_signed(19003, LUT_AMPL_WIDTH),
		26316 => to_signed(19001, LUT_AMPL_WIDTH),
		26317 => to_signed(18998, LUT_AMPL_WIDTH),
		26318 => to_signed(18996, LUT_AMPL_WIDTH),
		26319 => to_signed(18993, LUT_AMPL_WIDTH),
		26320 => to_signed(18991, LUT_AMPL_WIDTH),
		26321 => to_signed(18988, LUT_AMPL_WIDTH),
		26322 => to_signed(18985, LUT_AMPL_WIDTH),
		26323 => to_signed(18983, LUT_AMPL_WIDTH),
		26324 => to_signed(18980, LUT_AMPL_WIDTH),
		26325 => to_signed(18978, LUT_AMPL_WIDTH),
		26326 => to_signed(18975, LUT_AMPL_WIDTH),
		26327 => to_signed(18973, LUT_AMPL_WIDTH),
		26328 => to_signed(18970, LUT_AMPL_WIDTH),
		26329 => to_signed(18968, LUT_AMPL_WIDTH),
		26330 => to_signed(18965, LUT_AMPL_WIDTH),
		26331 => to_signed(18962, LUT_AMPL_WIDTH),
		26332 => to_signed(18960, LUT_AMPL_WIDTH),
		26333 => to_signed(18957, LUT_AMPL_WIDTH),
		26334 => to_signed(18955, LUT_AMPL_WIDTH),
		26335 => to_signed(18952, LUT_AMPL_WIDTH),
		26336 => to_signed(18950, LUT_AMPL_WIDTH),
		26337 => to_signed(18947, LUT_AMPL_WIDTH),
		26338 => to_signed(18944, LUT_AMPL_WIDTH),
		26339 => to_signed(18942, LUT_AMPL_WIDTH),
		26340 => to_signed(18939, LUT_AMPL_WIDTH),
		26341 => to_signed(18937, LUT_AMPL_WIDTH),
		26342 => to_signed(18934, LUT_AMPL_WIDTH),
		26343 => to_signed(18932, LUT_AMPL_WIDTH),
		26344 => to_signed(18929, LUT_AMPL_WIDTH),
		26345 => to_signed(18927, LUT_AMPL_WIDTH),
		26346 => to_signed(18924, LUT_AMPL_WIDTH),
		26347 => to_signed(18921, LUT_AMPL_WIDTH),
		26348 => to_signed(18919, LUT_AMPL_WIDTH),
		26349 => to_signed(18916, LUT_AMPL_WIDTH),
		26350 => to_signed(18914, LUT_AMPL_WIDTH),
		26351 => to_signed(18911, LUT_AMPL_WIDTH),
		26352 => to_signed(18909, LUT_AMPL_WIDTH),
		26353 => to_signed(18906, LUT_AMPL_WIDTH),
		26354 => to_signed(18903, LUT_AMPL_WIDTH),
		26355 => to_signed(18901, LUT_AMPL_WIDTH),
		26356 => to_signed(18898, LUT_AMPL_WIDTH),
		26357 => to_signed(18896, LUT_AMPL_WIDTH),
		26358 => to_signed(18893, LUT_AMPL_WIDTH),
		26359 => to_signed(18891, LUT_AMPL_WIDTH),
		26360 => to_signed(18888, LUT_AMPL_WIDTH),
		26361 => to_signed(18885, LUT_AMPL_WIDTH),
		26362 => to_signed(18883, LUT_AMPL_WIDTH),
		26363 => to_signed(18880, LUT_AMPL_WIDTH),
		26364 => to_signed(18878, LUT_AMPL_WIDTH),
		26365 => to_signed(18875, LUT_AMPL_WIDTH),
		26366 => to_signed(18873, LUT_AMPL_WIDTH),
		26367 => to_signed(18870, LUT_AMPL_WIDTH),
		26368 => to_signed(18868, LUT_AMPL_WIDTH),
		26369 => to_signed(18865, LUT_AMPL_WIDTH),
		26370 => to_signed(18862, LUT_AMPL_WIDTH),
		26371 => to_signed(18860, LUT_AMPL_WIDTH),
		26372 => to_signed(18857, LUT_AMPL_WIDTH),
		26373 => to_signed(18855, LUT_AMPL_WIDTH),
		26374 => to_signed(18852, LUT_AMPL_WIDTH),
		26375 => to_signed(18850, LUT_AMPL_WIDTH),
		26376 => to_signed(18847, LUT_AMPL_WIDTH),
		26377 => to_signed(18844, LUT_AMPL_WIDTH),
		26378 => to_signed(18842, LUT_AMPL_WIDTH),
		26379 => to_signed(18839, LUT_AMPL_WIDTH),
		26380 => to_signed(18837, LUT_AMPL_WIDTH),
		26381 => to_signed(18834, LUT_AMPL_WIDTH),
		26382 => to_signed(18832, LUT_AMPL_WIDTH),
		26383 => to_signed(18829, LUT_AMPL_WIDTH),
		26384 => to_signed(18826, LUT_AMPL_WIDTH),
		26385 => to_signed(18824, LUT_AMPL_WIDTH),
		26386 => to_signed(18821, LUT_AMPL_WIDTH),
		26387 => to_signed(18819, LUT_AMPL_WIDTH),
		26388 => to_signed(18816, LUT_AMPL_WIDTH),
		26389 => to_signed(18814, LUT_AMPL_WIDTH),
		26390 => to_signed(18811, LUT_AMPL_WIDTH),
		26391 => to_signed(18808, LUT_AMPL_WIDTH),
		26392 => to_signed(18806, LUT_AMPL_WIDTH),
		26393 => to_signed(18803, LUT_AMPL_WIDTH),
		26394 => to_signed(18801, LUT_AMPL_WIDTH),
		26395 => to_signed(18798, LUT_AMPL_WIDTH),
		26396 => to_signed(18796, LUT_AMPL_WIDTH),
		26397 => to_signed(18793, LUT_AMPL_WIDTH),
		26398 => to_signed(18790, LUT_AMPL_WIDTH),
		26399 => to_signed(18788, LUT_AMPL_WIDTH),
		26400 => to_signed(18785, LUT_AMPL_WIDTH),
		26401 => to_signed(18783, LUT_AMPL_WIDTH),
		26402 => to_signed(18780, LUT_AMPL_WIDTH),
		26403 => to_signed(18778, LUT_AMPL_WIDTH),
		26404 => to_signed(18775, LUT_AMPL_WIDTH),
		26405 => to_signed(18772, LUT_AMPL_WIDTH),
		26406 => to_signed(18770, LUT_AMPL_WIDTH),
		26407 => to_signed(18767, LUT_AMPL_WIDTH),
		26408 => to_signed(18765, LUT_AMPL_WIDTH),
		26409 => to_signed(18762, LUT_AMPL_WIDTH),
		26410 => to_signed(18759, LUT_AMPL_WIDTH),
		26411 => to_signed(18757, LUT_AMPL_WIDTH),
		26412 => to_signed(18754, LUT_AMPL_WIDTH),
		26413 => to_signed(18752, LUT_AMPL_WIDTH),
		26414 => to_signed(18749, LUT_AMPL_WIDTH),
		26415 => to_signed(18747, LUT_AMPL_WIDTH),
		26416 => to_signed(18744, LUT_AMPL_WIDTH),
		26417 => to_signed(18741, LUT_AMPL_WIDTH),
		26418 => to_signed(18739, LUT_AMPL_WIDTH),
		26419 => to_signed(18736, LUT_AMPL_WIDTH),
		26420 => to_signed(18734, LUT_AMPL_WIDTH),
		26421 => to_signed(18731, LUT_AMPL_WIDTH),
		26422 => to_signed(18729, LUT_AMPL_WIDTH),
		26423 => to_signed(18726, LUT_AMPL_WIDTH),
		26424 => to_signed(18723, LUT_AMPL_WIDTH),
		26425 => to_signed(18721, LUT_AMPL_WIDTH),
		26426 => to_signed(18718, LUT_AMPL_WIDTH),
		26427 => to_signed(18716, LUT_AMPL_WIDTH),
		26428 => to_signed(18713, LUT_AMPL_WIDTH),
		26429 => to_signed(18711, LUT_AMPL_WIDTH),
		26430 => to_signed(18708, LUT_AMPL_WIDTH),
		26431 => to_signed(18705, LUT_AMPL_WIDTH),
		26432 => to_signed(18703, LUT_AMPL_WIDTH),
		26433 => to_signed(18700, LUT_AMPL_WIDTH),
		26434 => to_signed(18698, LUT_AMPL_WIDTH),
		26435 => to_signed(18695, LUT_AMPL_WIDTH),
		26436 => to_signed(18692, LUT_AMPL_WIDTH),
		26437 => to_signed(18690, LUT_AMPL_WIDTH),
		26438 => to_signed(18687, LUT_AMPL_WIDTH),
		26439 => to_signed(18685, LUT_AMPL_WIDTH),
		26440 => to_signed(18682, LUT_AMPL_WIDTH),
		26441 => to_signed(18680, LUT_AMPL_WIDTH),
		26442 => to_signed(18677, LUT_AMPL_WIDTH),
		26443 => to_signed(18674, LUT_AMPL_WIDTH),
		26444 => to_signed(18672, LUT_AMPL_WIDTH),
		26445 => to_signed(18669, LUT_AMPL_WIDTH),
		26446 => to_signed(18667, LUT_AMPL_WIDTH),
		26447 => to_signed(18664, LUT_AMPL_WIDTH),
		26448 => to_signed(18661, LUT_AMPL_WIDTH),
		26449 => to_signed(18659, LUT_AMPL_WIDTH),
		26450 => to_signed(18656, LUT_AMPL_WIDTH),
		26451 => to_signed(18654, LUT_AMPL_WIDTH),
		26452 => to_signed(18651, LUT_AMPL_WIDTH),
		26453 => to_signed(18649, LUT_AMPL_WIDTH),
		26454 => to_signed(18646, LUT_AMPL_WIDTH),
		26455 => to_signed(18643, LUT_AMPL_WIDTH),
		26456 => to_signed(18641, LUT_AMPL_WIDTH),
		26457 => to_signed(18638, LUT_AMPL_WIDTH),
		26458 => to_signed(18636, LUT_AMPL_WIDTH),
		26459 => to_signed(18633, LUT_AMPL_WIDTH),
		26460 => to_signed(18630, LUT_AMPL_WIDTH),
		26461 => to_signed(18628, LUT_AMPL_WIDTH),
		26462 => to_signed(18625, LUT_AMPL_WIDTH),
		26463 => to_signed(18623, LUT_AMPL_WIDTH),
		26464 => to_signed(18620, LUT_AMPL_WIDTH),
		26465 => to_signed(18618, LUT_AMPL_WIDTH),
		26466 => to_signed(18615, LUT_AMPL_WIDTH),
		26467 => to_signed(18612, LUT_AMPL_WIDTH),
		26468 => to_signed(18610, LUT_AMPL_WIDTH),
		26469 => to_signed(18607, LUT_AMPL_WIDTH),
		26470 => to_signed(18605, LUT_AMPL_WIDTH),
		26471 => to_signed(18602, LUT_AMPL_WIDTH),
		26472 => to_signed(18599, LUT_AMPL_WIDTH),
		26473 => to_signed(18597, LUT_AMPL_WIDTH),
		26474 => to_signed(18594, LUT_AMPL_WIDTH),
		26475 => to_signed(18592, LUT_AMPL_WIDTH),
		26476 => to_signed(18589, LUT_AMPL_WIDTH),
		26477 => to_signed(18587, LUT_AMPL_WIDTH),
		26478 => to_signed(18584, LUT_AMPL_WIDTH),
		26479 => to_signed(18581, LUT_AMPL_WIDTH),
		26480 => to_signed(18579, LUT_AMPL_WIDTH),
		26481 => to_signed(18576, LUT_AMPL_WIDTH),
		26482 => to_signed(18574, LUT_AMPL_WIDTH),
		26483 => to_signed(18571, LUT_AMPL_WIDTH),
		26484 => to_signed(18568, LUT_AMPL_WIDTH),
		26485 => to_signed(18566, LUT_AMPL_WIDTH),
		26486 => to_signed(18563, LUT_AMPL_WIDTH),
		26487 => to_signed(18561, LUT_AMPL_WIDTH),
		26488 => to_signed(18558, LUT_AMPL_WIDTH),
		26489 => to_signed(18555, LUT_AMPL_WIDTH),
		26490 => to_signed(18553, LUT_AMPL_WIDTH),
		26491 => to_signed(18550, LUT_AMPL_WIDTH),
		26492 => to_signed(18548, LUT_AMPL_WIDTH),
		26493 => to_signed(18545, LUT_AMPL_WIDTH),
		26494 => to_signed(18543, LUT_AMPL_WIDTH),
		26495 => to_signed(18540, LUT_AMPL_WIDTH),
		26496 => to_signed(18537, LUT_AMPL_WIDTH),
		26497 => to_signed(18535, LUT_AMPL_WIDTH),
		26498 => to_signed(18532, LUT_AMPL_WIDTH),
		26499 => to_signed(18530, LUT_AMPL_WIDTH),
		26500 => to_signed(18527, LUT_AMPL_WIDTH),
		26501 => to_signed(18524, LUT_AMPL_WIDTH),
		26502 => to_signed(18522, LUT_AMPL_WIDTH),
		26503 => to_signed(18519, LUT_AMPL_WIDTH),
		26504 => to_signed(18517, LUT_AMPL_WIDTH),
		26505 => to_signed(18514, LUT_AMPL_WIDTH),
		26506 => to_signed(18511, LUT_AMPL_WIDTH),
		26507 => to_signed(18509, LUT_AMPL_WIDTH),
		26508 => to_signed(18506, LUT_AMPL_WIDTH),
		26509 => to_signed(18504, LUT_AMPL_WIDTH),
		26510 => to_signed(18501, LUT_AMPL_WIDTH),
		26511 => to_signed(18498, LUT_AMPL_WIDTH),
		26512 => to_signed(18496, LUT_AMPL_WIDTH),
		26513 => to_signed(18493, LUT_AMPL_WIDTH),
		26514 => to_signed(18491, LUT_AMPL_WIDTH),
		26515 => to_signed(18488, LUT_AMPL_WIDTH),
		26516 => to_signed(18485, LUT_AMPL_WIDTH),
		26517 => to_signed(18483, LUT_AMPL_WIDTH),
		26518 => to_signed(18480, LUT_AMPL_WIDTH),
		26519 => to_signed(18478, LUT_AMPL_WIDTH),
		26520 => to_signed(18475, LUT_AMPL_WIDTH),
		26521 => to_signed(18473, LUT_AMPL_WIDTH),
		26522 => to_signed(18470, LUT_AMPL_WIDTH),
		26523 => to_signed(18467, LUT_AMPL_WIDTH),
		26524 => to_signed(18465, LUT_AMPL_WIDTH),
		26525 => to_signed(18462, LUT_AMPL_WIDTH),
		26526 => to_signed(18460, LUT_AMPL_WIDTH),
		26527 => to_signed(18457, LUT_AMPL_WIDTH),
		26528 => to_signed(18454, LUT_AMPL_WIDTH),
		26529 => to_signed(18452, LUT_AMPL_WIDTH),
		26530 => to_signed(18449, LUT_AMPL_WIDTH),
		26531 => to_signed(18447, LUT_AMPL_WIDTH),
		26532 => to_signed(18444, LUT_AMPL_WIDTH),
		26533 => to_signed(18441, LUT_AMPL_WIDTH),
		26534 => to_signed(18439, LUT_AMPL_WIDTH),
		26535 => to_signed(18436, LUT_AMPL_WIDTH),
		26536 => to_signed(18434, LUT_AMPL_WIDTH),
		26537 => to_signed(18431, LUT_AMPL_WIDTH),
		26538 => to_signed(18428, LUT_AMPL_WIDTH),
		26539 => to_signed(18426, LUT_AMPL_WIDTH),
		26540 => to_signed(18423, LUT_AMPL_WIDTH),
		26541 => to_signed(18421, LUT_AMPL_WIDTH),
		26542 => to_signed(18418, LUT_AMPL_WIDTH),
		26543 => to_signed(18415, LUT_AMPL_WIDTH),
		26544 => to_signed(18413, LUT_AMPL_WIDTH),
		26545 => to_signed(18410, LUT_AMPL_WIDTH),
		26546 => to_signed(18408, LUT_AMPL_WIDTH),
		26547 => to_signed(18405, LUT_AMPL_WIDTH),
		26548 => to_signed(18402, LUT_AMPL_WIDTH),
		26549 => to_signed(18400, LUT_AMPL_WIDTH),
		26550 => to_signed(18397, LUT_AMPL_WIDTH),
		26551 => to_signed(18395, LUT_AMPL_WIDTH),
		26552 => to_signed(18392, LUT_AMPL_WIDTH),
		26553 => to_signed(18389, LUT_AMPL_WIDTH),
		26554 => to_signed(18387, LUT_AMPL_WIDTH),
		26555 => to_signed(18384, LUT_AMPL_WIDTH),
		26556 => to_signed(18382, LUT_AMPL_WIDTH),
		26557 => to_signed(18379, LUT_AMPL_WIDTH),
		26558 => to_signed(18376, LUT_AMPL_WIDTH),
		26559 => to_signed(18374, LUT_AMPL_WIDTH),
		26560 => to_signed(18371, LUT_AMPL_WIDTH),
		26561 => to_signed(18369, LUT_AMPL_WIDTH),
		26562 => to_signed(18366, LUT_AMPL_WIDTH),
		26563 => to_signed(18363, LUT_AMPL_WIDTH),
		26564 => to_signed(18361, LUT_AMPL_WIDTH),
		26565 => to_signed(18358, LUT_AMPL_WIDTH),
		26566 => to_signed(18356, LUT_AMPL_WIDTH),
		26567 => to_signed(18353, LUT_AMPL_WIDTH),
		26568 => to_signed(18350, LUT_AMPL_WIDTH),
		26569 => to_signed(18348, LUT_AMPL_WIDTH),
		26570 => to_signed(18345, LUT_AMPL_WIDTH),
		26571 => to_signed(18343, LUT_AMPL_WIDTH),
		26572 => to_signed(18340, LUT_AMPL_WIDTH),
		26573 => to_signed(18337, LUT_AMPL_WIDTH),
		26574 => to_signed(18335, LUT_AMPL_WIDTH),
		26575 => to_signed(18332, LUT_AMPL_WIDTH),
		26576 => to_signed(18330, LUT_AMPL_WIDTH),
		26577 => to_signed(18327, LUT_AMPL_WIDTH),
		26578 => to_signed(18324, LUT_AMPL_WIDTH),
		26579 => to_signed(18322, LUT_AMPL_WIDTH),
		26580 => to_signed(18319, LUT_AMPL_WIDTH),
		26581 => to_signed(18317, LUT_AMPL_WIDTH),
		26582 => to_signed(18314, LUT_AMPL_WIDTH),
		26583 => to_signed(18311, LUT_AMPL_WIDTH),
		26584 => to_signed(18309, LUT_AMPL_WIDTH),
		26585 => to_signed(18306, LUT_AMPL_WIDTH),
		26586 => to_signed(18304, LUT_AMPL_WIDTH),
		26587 => to_signed(18301, LUT_AMPL_WIDTH),
		26588 => to_signed(18298, LUT_AMPL_WIDTH),
		26589 => to_signed(18296, LUT_AMPL_WIDTH),
		26590 => to_signed(18293, LUT_AMPL_WIDTH),
		26591 => to_signed(18290, LUT_AMPL_WIDTH),
		26592 => to_signed(18288, LUT_AMPL_WIDTH),
		26593 => to_signed(18285, LUT_AMPL_WIDTH),
		26594 => to_signed(18283, LUT_AMPL_WIDTH),
		26595 => to_signed(18280, LUT_AMPL_WIDTH),
		26596 => to_signed(18277, LUT_AMPL_WIDTH),
		26597 => to_signed(18275, LUT_AMPL_WIDTH),
		26598 => to_signed(18272, LUT_AMPL_WIDTH),
		26599 => to_signed(18270, LUT_AMPL_WIDTH),
		26600 => to_signed(18267, LUT_AMPL_WIDTH),
		26601 => to_signed(18264, LUT_AMPL_WIDTH),
		26602 => to_signed(18262, LUT_AMPL_WIDTH),
		26603 => to_signed(18259, LUT_AMPL_WIDTH),
		26604 => to_signed(18257, LUT_AMPL_WIDTH),
		26605 => to_signed(18254, LUT_AMPL_WIDTH),
		26606 => to_signed(18251, LUT_AMPL_WIDTH),
		26607 => to_signed(18249, LUT_AMPL_WIDTH),
		26608 => to_signed(18246, LUT_AMPL_WIDTH),
		26609 => to_signed(18244, LUT_AMPL_WIDTH),
		26610 => to_signed(18241, LUT_AMPL_WIDTH),
		26611 => to_signed(18238, LUT_AMPL_WIDTH),
		26612 => to_signed(18236, LUT_AMPL_WIDTH),
		26613 => to_signed(18233, LUT_AMPL_WIDTH),
		26614 => to_signed(18230, LUT_AMPL_WIDTH),
		26615 => to_signed(18228, LUT_AMPL_WIDTH),
		26616 => to_signed(18225, LUT_AMPL_WIDTH),
		26617 => to_signed(18223, LUT_AMPL_WIDTH),
		26618 => to_signed(18220, LUT_AMPL_WIDTH),
		26619 => to_signed(18217, LUT_AMPL_WIDTH),
		26620 => to_signed(18215, LUT_AMPL_WIDTH),
		26621 => to_signed(18212, LUT_AMPL_WIDTH),
		26622 => to_signed(18210, LUT_AMPL_WIDTH),
		26623 => to_signed(18207, LUT_AMPL_WIDTH),
		26624 => to_signed(18204, LUT_AMPL_WIDTH),
		26625 => to_signed(18202, LUT_AMPL_WIDTH),
		26626 => to_signed(18199, LUT_AMPL_WIDTH),
		26627 => to_signed(18197, LUT_AMPL_WIDTH),
		26628 => to_signed(18194, LUT_AMPL_WIDTH),
		26629 => to_signed(18191, LUT_AMPL_WIDTH),
		26630 => to_signed(18189, LUT_AMPL_WIDTH),
		26631 => to_signed(18186, LUT_AMPL_WIDTH),
		26632 => to_signed(18183, LUT_AMPL_WIDTH),
		26633 => to_signed(18181, LUT_AMPL_WIDTH),
		26634 => to_signed(18178, LUT_AMPL_WIDTH),
		26635 => to_signed(18176, LUT_AMPL_WIDTH),
		26636 => to_signed(18173, LUT_AMPL_WIDTH),
		26637 => to_signed(18170, LUT_AMPL_WIDTH),
		26638 => to_signed(18168, LUT_AMPL_WIDTH),
		26639 => to_signed(18165, LUT_AMPL_WIDTH),
		26640 => to_signed(18163, LUT_AMPL_WIDTH),
		26641 => to_signed(18160, LUT_AMPL_WIDTH),
		26642 => to_signed(18157, LUT_AMPL_WIDTH),
		26643 => to_signed(18155, LUT_AMPL_WIDTH),
		26644 => to_signed(18152, LUT_AMPL_WIDTH),
		26645 => to_signed(18149, LUT_AMPL_WIDTH),
		26646 => to_signed(18147, LUT_AMPL_WIDTH),
		26647 => to_signed(18144, LUT_AMPL_WIDTH),
		26648 => to_signed(18142, LUT_AMPL_WIDTH),
		26649 => to_signed(18139, LUT_AMPL_WIDTH),
		26650 => to_signed(18136, LUT_AMPL_WIDTH),
		26651 => to_signed(18134, LUT_AMPL_WIDTH),
		26652 => to_signed(18131, LUT_AMPL_WIDTH),
		26653 => to_signed(18129, LUT_AMPL_WIDTH),
		26654 => to_signed(18126, LUT_AMPL_WIDTH),
		26655 => to_signed(18123, LUT_AMPL_WIDTH),
		26656 => to_signed(18121, LUT_AMPL_WIDTH),
		26657 => to_signed(18118, LUT_AMPL_WIDTH),
		26658 => to_signed(18115, LUT_AMPL_WIDTH),
		26659 => to_signed(18113, LUT_AMPL_WIDTH),
		26660 => to_signed(18110, LUT_AMPL_WIDTH),
		26661 => to_signed(18108, LUT_AMPL_WIDTH),
		26662 => to_signed(18105, LUT_AMPL_WIDTH),
		26663 => to_signed(18102, LUT_AMPL_WIDTH),
		26664 => to_signed(18100, LUT_AMPL_WIDTH),
		26665 => to_signed(18097, LUT_AMPL_WIDTH),
		26666 => to_signed(18095, LUT_AMPL_WIDTH),
		26667 => to_signed(18092, LUT_AMPL_WIDTH),
		26668 => to_signed(18089, LUT_AMPL_WIDTH),
		26669 => to_signed(18087, LUT_AMPL_WIDTH),
		26670 => to_signed(18084, LUT_AMPL_WIDTH),
		26671 => to_signed(18081, LUT_AMPL_WIDTH),
		26672 => to_signed(18079, LUT_AMPL_WIDTH),
		26673 => to_signed(18076, LUT_AMPL_WIDTH),
		26674 => to_signed(18074, LUT_AMPL_WIDTH),
		26675 => to_signed(18071, LUT_AMPL_WIDTH),
		26676 => to_signed(18068, LUT_AMPL_WIDTH),
		26677 => to_signed(18066, LUT_AMPL_WIDTH),
		26678 => to_signed(18063, LUT_AMPL_WIDTH),
		26679 => to_signed(18060, LUT_AMPL_WIDTH),
		26680 => to_signed(18058, LUT_AMPL_WIDTH),
		26681 => to_signed(18055, LUT_AMPL_WIDTH),
		26682 => to_signed(18053, LUT_AMPL_WIDTH),
		26683 => to_signed(18050, LUT_AMPL_WIDTH),
		26684 => to_signed(18047, LUT_AMPL_WIDTH),
		26685 => to_signed(18045, LUT_AMPL_WIDTH),
		26686 => to_signed(18042, LUT_AMPL_WIDTH),
		26687 => to_signed(18039, LUT_AMPL_WIDTH),
		26688 => to_signed(18037, LUT_AMPL_WIDTH),
		26689 => to_signed(18034, LUT_AMPL_WIDTH),
		26690 => to_signed(18032, LUT_AMPL_WIDTH),
		26691 => to_signed(18029, LUT_AMPL_WIDTH),
		26692 => to_signed(18026, LUT_AMPL_WIDTH),
		26693 => to_signed(18024, LUT_AMPL_WIDTH),
		26694 => to_signed(18021, LUT_AMPL_WIDTH),
		26695 => to_signed(18018, LUT_AMPL_WIDTH),
		26696 => to_signed(18016, LUT_AMPL_WIDTH),
		26697 => to_signed(18013, LUT_AMPL_WIDTH),
		26698 => to_signed(18011, LUT_AMPL_WIDTH),
		26699 => to_signed(18008, LUT_AMPL_WIDTH),
		26700 => to_signed(18005, LUT_AMPL_WIDTH),
		26701 => to_signed(18003, LUT_AMPL_WIDTH),
		26702 => to_signed(18000, LUT_AMPL_WIDTH),
		26703 => to_signed(17997, LUT_AMPL_WIDTH),
		26704 => to_signed(17995, LUT_AMPL_WIDTH),
		26705 => to_signed(17992, LUT_AMPL_WIDTH),
		26706 => to_signed(17990, LUT_AMPL_WIDTH),
		26707 => to_signed(17987, LUT_AMPL_WIDTH),
		26708 => to_signed(17984, LUT_AMPL_WIDTH),
		26709 => to_signed(17982, LUT_AMPL_WIDTH),
		26710 => to_signed(17979, LUT_AMPL_WIDTH),
		26711 => to_signed(17976, LUT_AMPL_WIDTH),
		26712 => to_signed(17974, LUT_AMPL_WIDTH),
		26713 => to_signed(17971, LUT_AMPL_WIDTH),
		26714 => to_signed(17969, LUT_AMPL_WIDTH),
		26715 => to_signed(17966, LUT_AMPL_WIDTH),
		26716 => to_signed(17963, LUT_AMPL_WIDTH),
		26717 => to_signed(17961, LUT_AMPL_WIDTH),
		26718 => to_signed(17958, LUT_AMPL_WIDTH),
		26719 => to_signed(17955, LUT_AMPL_WIDTH),
		26720 => to_signed(17953, LUT_AMPL_WIDTH),
		26721 => to_signed(17950, LUT_AMPL_WIDTH),
		26722 => to_signed(17948, LUT_AMPL_WIDTH),
		26723 => to_signed(17945, LUT_AMPL_WIDTH),
		26724 => to_signed(17942, LUT_AMPL_WIDTH),
		26725 => to_signed(17940, LUT_AMPL_WIDTH),
		26726 => to_signed(17937, LUT_AMPL_WIDTH),
		26727 => to_signed(17934, LUT_AMPL_WIDTH),
		26728 => to_signed(17932, LUT_AMPL_WIDTH),
		26729 => to_signed(17929, LUT_AMPL_WIDTH),
		26730 => to_signed(17927, LUT_AMPL_WIDTH),
		26731 => to_signed(17924, LUT_AMPL_WIDTH),
		26732 => to_signed(17921, LUT_AMPL_WIDTH),
		26733 => to_signed(17919, LUT_AMPL_WIDTH),
		26734 => to_signed(17916, LUT_AMPL_WIDTH),
		26735 => to_signed(17913, LUT_AMPL_WIDTH),
		26736 => to_signed(17911, LUT_AMPL_WIDTH),
		26737 => to_signed(17908, LUT_AMPL_WIDTH),
		26738 => to_signed(17906, LUT_AMPL_WIDTH),
		26739 => to_signed(17903, LUT_AMPL_WIDTH),
		26740 => to_signed(17900, LUT_AMPL_WIDTH),
		26741 => to_signed(17898, LUT_AMPL_WIDTH),
		26742 => to_signed(17895, LUT_AMPL_WIDTH),
		26743 => to_signed(17892, LUT_AMPL_WIDTH),
		26744 => to_signed(17890, LUT_AMPL_WIDTH),
		26745 => to_signed(17887, LUT_AMPL_WIDTH),
		26746 => to_signed(17884, LUT_AMPL_WIDTH),
		26747 => to_signed(17882, LUT_AMPL_WIDTH),
		26748 => to_signed(17879, LUT_AMPL_WIDTH),
		26749 => to_signed(17877, LUT_AMPL_WIDTH),
		26750 => to_signed(17874, LUT_AMPL_WIDTH),
		26751 => to_signed(17871, LUT_AMPL_WIDTH),
		26752 => to_signed(17869, LUT_AMPL_WIDTH),
		26753 => to_signed(17866, LUT_AMPL_WIDTH),
		26754 => to_signed(17863, LUT_AMPL_WIDTH),
		26755 => to_signed(17861, LUT_AMPL_WIDTH),
		26756 => to_signed(17858, LUT_AMPL_WIDTH),
		26757 => to_signed(17855, LUT_AMPL_WIDTH),
		26758 => to_signed(17853, LUT_AMPL_WIDTH),
		26759 => to_signed(17850, LUT_AMPL_WIDTH),
		26760 => to_signed(17848, LUT_AMPL_WIDTH),
		26761 => to_signed(17845, LUT_AMPL_WIDTH),
		26762 => to_signed(17842, LUT_AMPL_WIDTH),
		26763 => to_signed(17840, LUT_AMPL_WIDTH),
		26764 => to_signed(17837, LUT_AMPL_WIDTH),
		26765 => to_signed(17834, LUT_AMPL_WIDTH),
		26766 => to_signed(17832, LUT_AMPL_WIDTH),
		26767 => to_signed(17829, LUT_AMPL_WIDTH),
		26768 => to_signed(17827, LUT_AMPL_WIDTH),
		26769 => to_signed(17824, LUT_AMPL_WIDTH),
		26770 => to_signed(17821, LUT_AMPL_WIDTH),
		26771 => to_signed(17819, LUT_AMPL_WIDTH),
		26772 => to_signed(17816, LUT_AMPL_WIDTH),
		26773 => to_signed(17813, LUT_AMPL_WIDTH),
		26774 => to_signed(17811, LUT_AMPL_WIDTH),
		26775 => to_signed(17808, LUT_AMPL_WIDTH),
		26776 => to_signed(17805, LUT_AMPL_WIDTH),
		26777 => to_signed(17803, LUT_AMPL_WIDTH),
		26778 => to_signed(17800, LUT_AMPL_WIDTH),
		26779 => to_signed(17798, LUT_AMPL_WIDTH),
		26780 => to_signed(17795, LUT_AMPL_WIDTH),
		26781 => to_signed(17792, LUT_AMPL_WIDTH),
		26782 => to_signed(17790, LUT_AMPL_WIDTH),
		26783 => to_signed(17787, LUT_AMPL_WIDTH),
		26784 => to_signed(17784, LUT_AMPL_WIDTH),
		26785 => to_signed(17782, LUT_AMPL_WIDTH),
		26786 => to_signed(17779, LUT_AMPL_WIDTH),
		26787 => to_signed(17776, LUT_AMPL_WIDTH),
		26788 => to_signed(17774, LUT_AMPL_WIDTH),
		26789 => to_signed(17771, LUT_AMPL_WIDTH),
		26790 => to_signed(17768, LUT_AMPL_WIDTH),
		26791 => to_signed(17766, LUT_AMPL_WIDTH),
		26792 => to_signed(17763, LUT_AMPL_WIDTH),
		26793 => to_signed(17761, LUT_AMPL_WIDTH),
		26794 => to_signed(17758, LUT_AMPL_WIDTH),
		26795 => to_signed(17755, LUT_AMPL_WIDTH),
		26796 => to_signed(17753, LUT_AMPL_WIDTH),
		26797 => to_signed(17750, LUT_AMPL_WIDTH),
		26798 => to_signed(17747, LUT_AMPL_WIDTH),
		26799 => to_signed(17745, LUT_AMPL_WIDTH),
		26800 => to_signed(17742, LUT_AMPL_WIDTH),
		26801 => to_signed(17739, LUT_AMPL_WIDTH),
		26802 => to_signed(17737, LUT_AMPL_WIDTH),
		26803 => to_signed(17734, LUT_AMPL_WIDTH),
		26804 => to_signed(17732, LUT_AMPL_WIDTH),
		26805 => to_signed(17729, LUT_AMPL_WIDTH),
		26806 => to_signed(17726, LUT_AMPL_WIDTH),
		26807 => to_signed(17724, LUT_AMPL_WIDTH),
		26808 => to_signed(17721, LUT_AMPL_WIDTH),
		26809 => to_signed(17718, LUT_AMPL_WIDTH),
		26810 => to_signed(17716, LUT_AMPL_WIDTH),
		26811 => to_signed(17713, LUT_AMPL_WIDTH),
		26812 => to_signed(17710, LUT_AMPL_WIDTH),
		26813 => to_signed(17708, LUT_AMPL_WIDTH),
		26814 => to_signed(17705, LUT_AMPL_WIDTH),
		26815 => to_signed(17702, LUT_AMPL_WIDTH),
		26816 => to_signed(17700, LUT_AMPL_WIDTH),
		26817 => to_signed(17697, LUT_AMPL_WIDTH),
		26818 => to_signed(17695, LUT_AMPL_WIDTH),
		26819 => to_signed(17692, LUT_AMPL_WIDTH),
		26820 => to_signed(17689, LUT_AMPL_WIDTH),
		26821 => to_signed(17687, LUT_AMPL_WIDTH),
		26822 => to_signed(17684, LUT_AMPL_WIDTH),
		26823 => to_signed(17681, LUT_AMPL_WIDTH),
		26824 => to_signed(17679, LUT_AMPL_WIDTH),
		26825 => to_signed(17676, LUT_AMPL_WIDTH),
		26826 => to_signed(17673, LUT_AMPL_WIDTH),
		26827 => to_signed(17671, LUT_AMPL_WIDTH),
		26828 => to_signed(17668, LUT_AMPL_WIDTH),
		26829 => to_signed(17665, LUT_AMPL_WIDTH),
		26830 => to_signed(17663, LUT_AMPL_WIDTH),
		26831 => to_signed(17660, LUT_AMPL_WIDTH),
		26832 => to_signed(17657, LUT_AMPL_WIDTH),
		26833 => to_signed(17655, LUT_AMPL_WIDTH),
		26834 => to_signed(17652, LUT_AMPL_WIDTH),
		26835 => to_signed(17650, LUT_AMPL_WIDTH),
		26836 => to_signed(17647, LUT_AMPL_WIDTH),
		26837 => to_signed(17644, LUT_AMPL_WIDTH),
		26838 => to_signed(17642, LUT_AMPL_WIDTH),
		26839 => to_signed(17639, LUT_AMPL_WIDTH),
		26840 => to_signed(17636, LUT_AMPL_WIDTH),
		26841 => to_signed(17634, LUT_AMPL_WIDTH),
		26842 => to_signed(17631, LUT_AMPL_WIDTH),
		26843 => to_signed(17628, LUT_AMPL_WIDTH),
		26844 => to_signed(17626, LUT_AMPL_WIDTH),
		26845 => to_signed(17623, LUT_AMPL_WIDTH),
		26846 => to_signed(17620, LUT_AMPL_WIDTH),
		26847 => to_signed(17618, LUT_AMPL_WIDTH),
		26848 => to_signed(17615, LUT_AMPL_WIDTH),
		26849 => to_signed(17612, LUT_AMPL_WIDTH),
		26850 => to_signed(17610, LUT_AMPL_WIDTH),
		26851 => to_signed(17607, LUT_AMPL_WIDTH),
		26852 => to_signed(17605, LUT_AMPL_WIDTH),
		26853 => to_signed(17602, LUT_AMPL_WIDTH),
		26854 => to_signed(17599, LUT_AMPL_WIDTH),
		26855 => to_signed(17597, LUT_AMPL_WIDTH),
		26856 => to_signed(17594, LUT_AMPL_WIDTH),
		26857 => to_signed(17591, LUT_AMPL_WIDTH),
		26858 => to_signed(17589, LUT_AMPL_WIDTH),
		26859 => to_signed(17586, LUT_AMPL_WIDTH),
		26860 => to_signed(17583, LUT_AMPL_WIDTH),
		26861 => to_signed(17581, LUT_AMPL_WIDTH),
		26862 => to_signed(17578, LUT_AMPL_WIDTH),
		26863 => to_signed(17575, LUT_AMPL_WIDTH),
		26864 => to_signed(17573, LUT_AMPL_WIDTH),
		26865 => to_signed(17570, LUT_AMPL_WIDTH),
		26866 => to_signed(17567, LUT_AMPL_WIDTH),
		26867 => to_signed(17565, LUT_AMPL_WIDTH),
		26868 => to_signed(17562, LUT_AMPL_WIDTH),
		26869 => to_signed(17559, LUT_AMPL_WIDTH),
		26870 => to_signed(17557, LUT_AMPL_WIDTH),
		26871 => to_signed(17554, LUT_AMPL_WIDTH),
		26872 => to_signed(17551, LUT_AMPL_WIDTH),
		26873 => to_signed(17549, LUT_AMPL_WIDTH),
		26874 => to_signed(17546, LUT_AMPL_WIDTH),
		26875 => to_signed(17544, LUT_AMPL_WIDTH),
		26876 => to_signed(17541, LUT_AMPL_WIDTH),
		26877 => to_signed(17538, LUT_AMPL_WIDTH),
		26878 => to_signed(17536, LUT_AMPL_WIDTH),
		26879 => to_signed(17533, LUT_AMPL_WIDTH),
		26880 => to_signed(17530, LUT_AMPL_WIDTH),
		26881 => to_signed(17528, LUT_AMPL_WIDTH),
		26882 => to_signed(17525, LUT_AMPL_WIDTH),
		26883 => to_signed(17522, LUT_AMPL_WIDTH),
		26884 => to_signed(17520, LUT_AMPL_WIDTH),
		26885 => to_signed(17517, LUT_AMPL_WIDTH),
		26886 => to_signed(17514, LUT_AMPL_WIDTH),
		26887 => to_signed(17512, LUT_AMPL_WIDTH),
		26888 => to_signed(17509, LUT_AMPL_WIDTH),
		26889 => to_signed(17506, LUT_AMPL_WIDTH),
		26890 => to_signed(17504, LUT_AMPL_WIDTH),
		26891 => to_signed(17501, LUT_AMPL_WIDTH),
		26892 => to_signed(17498, LUT_AMPL_WIDTH),
		26893 => to_signed(17496, LUT_AMPL_WIDTH),
		26894 => to_signed(17493, LUT_AMPL_WIDTH),
		26895 => to_signed(17490, LUT_AMPL_WIDTH),
		26896 => to_signed(17488, LUT_AMPL_WIDTH),
		26897 => to_signed(17485, LUT_AMPL_WIDTH),
		26898 => to_signed(17482, LUT_AMPL_WIDTH),
		26899 => to_signed(17480, LUT_AMPL_WIDTH),
		26900 => to_signed(17477, LUT_AMPL_WIDTH),
		26901 => to_signed(17474, LUT_AMPL_WIDTH),
		26902 => to_signed(17472, LUT_AMPL_WIDTH),
		26903 => to_signed(17469, LUT_AMPL_WIDTH),
		26904 => to_signed(17467, LUT_AMPL_WIDTH),
		26905 => to_signed(17464, LUT_AMPL_WIDTH),
		26906 => to_signed(17461, LUT_AMPL_WIDTH),
		26907 => to_signed(17459, LUT_AMPL_WIDTH),
		26908 => to_signed(17456, LUT_AMPL_WIDTH),
		26909 => to_signed(17453, LUT_AMPL_WIDTH),
		26910 => to_signed(17451, LUT_AMPL_WIDTH),
		26911 => to_signed(17448, LUT_AMPL_WIDTH),
		26912 => to_signed(17445, LUT_AMPL_WIDTH),
		26913 => to_signed(17443, LUT_AMPL_WIDTH),
		26914 => to_signed(17440, LUT_AMPL_WIDTH),
		26915 => to_signed(17437, LUT_AMPL_WIDTH),
		26916 => to_signed(17435, LUT_AMPL_WIDTH),
		26917 => to_signed(17432, LUT_AMPL_WIDTH),
		26918 => to_signed(17429, LUT_AMPL_WIDTH),
		26919 => to_signed(17427, LUT_AMPL_WIDTH),
		26920 => to_signed(17424, LUT_AMPL_WIDTH),
		26921 => to_signed(17421, LUT_AMPL_WIDTH),
		26922 => to_signed(17419, LUT_AMPL_WIDTH),
		26923 => to_signed(17416, LUT_AMPL_WIDTH),
		26924 => to_signed(17413, LUT_AMPL_WIDTH),
		26925 => to_signed(17411, LUT_AMPL_WIDTH),
		26926 => to_signed(17408, LUT_AMPL_WIDTH),
		26927 => to_signed(17405, LUT_AMPL_WIDTH),
		26928 => to_signed(17403, LUT_AMPL_WIDTH),
		26929 => to_signed(17400, LUT_AMPL_WIDTH),
		26930 => to_signed(17397, LUT_AMPL_WIDTH),
		26931 => to_signed(17395, LUT_AMPL_WIDTH),
		26932 => to_signed(17392, LUT_AMPL_WIDTH),
		26933 => to_signed(17389, LUT_AMPL_WIDTH),
		26934 => to_signed(17387, LUT_AMPL_WIDTH),
		26935 => to_signed(17384, LUT_AMPL_WIDTH),
		26936 => to_signed(17381, LUT_AMPL_WIDTH),
		26937 => to_signed(17379, LUT_AMPL_WIDTH),
		26938 => to_signed(17376, LUT_AMPL_WIDTH),
		26939 => to_signed(17373, LUT_AMPL_WIDTH),
		26940 => to_signed(17371, LUT_AMPL_WIDTH),
		26941 => to_signed(17368, LUT_AMPL_WIDTH),
		26942 => to_signed(17365, LUT_AMPL_WIDTH),
		26943 => to_signed(17363, LUT_AMPL_WIDTH),
		26944 => to_signed(17360, LUT_AMPL_WIDTH),
		26945 => to_signed(17357, LUT_AMPL_WIDTH),
		26946 => to_signed(17355, LUT_AMPL_WIDTH),
		26947 => to_signed(17352, LUT_AMPL_WIDTH),
		26948 => to_signed(17349, LUT_AMPL_WIDTH),
		26949 => to_signed(17347, LUT_AMPL_WIDTH),
		26950 => to_signed(17344, LUT_AMPL_WIDTH),
		26951 => to_signed(17341, LUT_AMPL_WIDTH),
		26952 => to_signed(17339, LUT_AMPL_WIDTH),
		26953 => to_signed(17336, LUT_AMPL_WIDTH),
		26954 => to_signed(17333, LUT_AMPL_WIDTH),
		26955 => to_signed(17331, LUT_AMPL_WIDTH),
		26956 => to_signed(17328, LUT_AMPL_WIDTH),
		26957 => to_signed(17325, LUT_AMPL_WIDTH),
		26958 => to_signed(17323, LUT_AMPL_WIDTH),
		26959 => to_signed(17320, LUT_AMPL_WIDTH),
		26960 => to_signed(17317, LUT_AMPL_WIDTH),
		26961 => to_signed(17315, LUT_AMPL_WIDTH),
		26962 => to_signed(17312, LUT_AMPL_WIDTH),
		26963 => to_signed(17309, LUT_AMPL_WIDTH),
		26964 => to_signed(17307, LUT_AMPL_WIDTH),
		26965 => to_signed(17304, LUT_AMPL_WIDTH),
		26966 => to_signed(17301, LUT_AMPL_WIDTH),
		26967 => to_signed(17299, LUT_AMPL_WIDTH),
		26968 => to_signed(17296, LUT_AMPL_WIDTH),
		26969 => to_signed(17293, LUT_AMPL_WIDTH),
		26970 => to_signed(17291, LUT_AMPL_WIDTH),
		26971 => to_signed(17288, LUT_AMPL_WIDTH),
		26972 => to_signed(17285, LUT_AMPL_WIDTH),
		26973 => to_signed(17283, LUT_AMPL_WIDTH),
		26974 => to_signed(17280, LUT_AMPL_WIDTH),
		26975 => to_signed(17277, LUT_AMPL_WIDTH),
		26976 => to_signed(17275, LUT_AMPL_WIDTH),
		26977 => to_signed(17272, LUT_AMPL_WIDTH),
		26978 => to_signed(17269, LUT_AMPL_WIDTH),
		26979 => to_signed(17267, LUT_AMPL_WIDTH),
		26980 => to_signed(17264, LUT_AMPL_WIDTH),
		26981 => to_signed(17261, LUT_AMPL_WIDTH),
		26982 => to_signed(17259, LUT_AMPL_WIDTH),
		26983 => to_signed(17256, LUT_AMPL_WIDTH),
		26984 => to_signed(17253, LUT_AMPL_WIDTH),
		26985 => to_signed(17251, LUT_AMPL_WIDTH),
		26986 => to_signed(17248, LUT_AMPL_WIDTH),
		26987 => to_signed(17245, LUT_AMPL_WIDTH),
		26988 => to_signed(17243, LUT_AMPL_WIDTH),
		26989 => to_signed(17240, LUT_AMPL_WIDTH),
		26990 => to_signed(17237, LUT_AMPL_WIDTH),
		26991 => to_signed(17235, LUT_AMPL_WIDTH),
		26992 => to_signed(17232, LUT_AMPL_WIDTH),
		26993 => to_signed(17229, LUT_AMPL_WIDTH),
		26994 => to_signed(17227, LUT_AMPL_WIDTH),
		26995 => to_signed(17224, LUT_AMPL_WIDTH),
		26996 => to_signed(17221, LUT_AMPL_WIDTH),
		26997 => to_signed(17219, LUT_AMPL_WIDTH),
		26998 => to_signed(17216, LUT_AMPL_WIDTH),
		26999 => to_signed(17213, LUT_AMPL_WIDTH),
		27000 => to_signed(17211, LUT_AMPL_WIDTH),
		27001 => to_signed(17208, LUT_AMPL_WIDTH),
		27002 => to_signed(17205, LUT_AMPL_WIDTH),
		27003 => to_signed(17203, LUT_AMPL_WIDTH),
		27004 => to_signed(17200, LUT_AMPL_WIDTH),
		27005 => to_signed(17197, LUT_AMPL_WIDTH),
		27006 => to_signed(17195, LUT_AMPL_WIDTH),
		27007 => to_signed(17192, LUT_AMPL_WIDTH),
		27008 => to_signed(17189, LUT_AMPL_WIDTH),
		27009 => to_signed(17187, LUT_AMPL_WIDTH),
		27010 => to_signed(17184, LUT_AMPL_WIDTH),
		27011 => to_signed(17181, LUT_AMPL_WIDTH),
		27012 => to_signed(17179, LUT_AMPL_WIDTH),
		27013 => to_signed(17176, LUT_AMPL_WIDTH),
		27014 => to_signed(17173, LUT_AMPL_WIDTH),
		27015 => to_signed(17171, LUT_AMPL_WIDTH),
		27016 => to_signed(17168, LUT_AMPL_WIDTH),
		27017 => to_signed(17165, LUT_AMPL_WIDTH),
		27018 => to_signed(17162, LUT_AMPL_WIDTH),
		27019 => to_signed(17160, LUT_AMPL_WIDTH),
		27020 => to_signed(17157, LUT_AMPL_WIDTH),
		27021 => to_signed(17154, LUT_AMPL_WIDTH),
		27022 => to_signed(17152, LUT_AMPL_WIDTH),
		27023 => to_signed(17149, LUT_AMPL_WIDTH),
		27024 => to_signed(17146, LUT_AMPL_WIDTH),
		27025 => to_signed(17144, LUT_AMPL_WIDTH),
		27026 => to_signed(17141, LUT_AMPL_WIDTH),
		27027 => to_signed(17138, LUT_AMPL_WIDTH),
		27028 => to_signed(17136, LUT_AMPL_WIDTH),
		27029 => to_signed(17133, LUT_AMPL_WIDTH),
		27030 => to_signed(17130, LUT_AMPL_WIDTH),
		27031 => to_signed(17128, LUT_AMPL_WIDTH),
		27032 => to_signed(17125, LUT_AMPL_WIDTH),
		27033 => to_signed(17122, LUT_AMPL_WIDTH),
		27034 => to_signed(17120, LUT_AMPL_WIDTH),
		27035 => to_signed(17117, LUT_AMPL_WIDTH),
		27036 => to_signed(17114, LUT_AMPL_WIDTH),
		27037 => to_signed(17112, LUT_AMPL_WIDTH),
		27038 => to_signed(17109, LUT_AMPL_WIDTH),
		27039 => to_signed(17106, LUT_AMPL_WIDTH),
		27040 => to_signed(17104, LUT_AMPL_WIDTH),
		27041 => to_signed(17101, LUT_AMPL_WIDTH),
		27042 => to_signed(17098, LUT_AMPL_WIDTH),
		27043 => to_signed(17096, LUT_AMPL_WIDTH),
		27044 => to_signed(17093, LUT_AMPL_WIDTH),
		27045 => to_signed(17090, LUT_AMPL_WIDTH),
		27046 => to_signed(17087, LUT_AMPL_WIDTH),
		27047 => to_signed(17085, LUT_AMPL_WIDTH),
		27048 => to_signed(17082, LUT_AMPL_WIDTH),
		27049 => to_signed(17079, LUT_AMPL_WIDTH),
		27050 => to_signed(17077, LUT_AMPL_WIDTH),
		27051 => to_signed(17074, LUT_AMPL_WIDTH),
		27052 => to_signed(17071, LUT_AMPL_WIDTH),
		27053 => to_signed(17069, LUT_AMPL_WIDTH),
		27054 => to_signed(17066, LUT_AMPL_WIDTH),
		27055 => to_signed(17063, LUT_AMPL_WIDTH),
		27056 => to_signed(17061, LUT_AMPL_WIDTH),
		27057 => to_signed(17058, LUT_AMPL_WIDTH),
		27058 => to_signed(17055, LUT_AMPL_WIDTH),
		27059 => to_signed(17053, LUT_AMPL_WIDTH),
		27060 => to_signed(17050, LUT_AMPL_WIDTH),
		27061 => to_signed(17047, LUT_AMPL_WIDTH),
		27062 => to_signed(17045, LUT_AMPL_WIDTH),
		27063 => to_signed(17042, LUT_AMPL_WIDTH),
		27064 => to_signed(17039, LUT_AMPL_WIDTH),
		27065 => to_signed(17037, LUT_AMPL_WIDTH),
		27066 => to_signed(17034, LUT_AMPL_WIDTH),
		27067 => to_signed(17031, LUT_AMPL_WIDTH),
		27068 => to_signed(17028, LUT_AMPL_WIDTH),
		27069 => to_signed(17026, LUT_AMPL_WIDTH),
		27070 => to_signed(17023, LUT_AMPL_WIDTH),
		27071 => to_signed(17020, LUT_AMPL_WIDTH),
		27072 => to_signed(17018, LUT_AMPL_WIDTH),
		27073 => to_signed(17015, LUT_AMPL_WIDTH),
		27074 => to_signed(17012, LUT_AMPL_WIDTH),
		27075 => to_signed(17010, LUT_AMPL_WIDTH),
		27076 => to_signed(17007, LUT_AMPL_WIDTH),
		27077 => to_signed(17004, LUT_AMPL_WIDTH),
		27078 => to_signed(17002, LUT_AMPL_WIDTH),
		27079 => to_signed(16999, LUT_AMPL_WIDTH),
		27080 => to_signed(16996, LUT_AMPL_WIDTH),
		27081 => to_signed(16994, LUT_AMPL_WIDTH),
		27082 => to_signed(16991, LUT_AMPL_WIDTH),
		27083 => to_signed(16988, LUT_AMPL_WIDTH),
		27084 => to_signed(16986, LUT_AMPL_WIDTH),
		27085 => to_signed(16983, LUT_AMPL_WIDTH),
		27086 => to_signed(16980, LUT_AMPL_WIDTH),
		27087 => to_signed(16977, LUT_AMPL_WIDTH),
		27088 => to_signed(16975, LUT_AMPL_WIDTH),
		27089 => to_signed(16972, LUT_AMPL_WIDTH),
		27090 => to_signed(16969, LUT_AMPL_WIDTH),
		27091 => to_signed(16967, LUT_AMPL_WIDTH),
		27092 => to_signed(16964, LUT_AMPL_WIDTH),
		27093 => to_signed(16961, LUT_AMPL_WIDTH),
		27094 => to_signed(16959, LUT_AMPL_WIDTH),
		27095 => to_signed(16956, LUT_AMPL_WIDTH),
		27096 => to_signed(16953, LUT_AMPL_WIDTH),
		27097 => to_signed(16951, LUT_AMPL_WIDTH),
		27098 => to_signed(16948, LUT_AMPL_WIDTH),
		27099 => to_signed(16945, LUT_AMPL_WIDTH),
		27100 => to_signed(16943, LUT_AMPL_WIDTH),
		27101 => to_signed(16940, LUT_AMPL_WIDTH),
		27102 => to_signed(16937, LUT_AMPL_WIDTH),
		27103 => to_signed(16934, LUT_AMPL_WIDTH),
		27104 => to_signed(16932, LUT_AMPL_WIDTH),
		27105 => to_signed(16929, LUT_AMPL_WIDTH),
		27106 => to_signed(16926, LUT_AMPL_WIDTH),
		27107 => to_signed(16924, LUT_AMPL_WIDTH),
		27108 => to_signed(16921, LUT_AMPL_WIDTH),
		27109 => to_signed(16918, LUT_AMPL_WIDTH),
		27110 => to_signed(16916, LUT_AMPL_WIDTH),
		27111 => to_signed(16913, LUT_AMPL_WIDTH),
		27112 => to_signed(16910, LUT_AMPL_WIDTH),
		27113 => to_signed(16908, LUT_AMPL_WIDTH),
		27114 => to_signed(16905, LUT_AMPL_WIDTH),
		27115 => to_signed(16902, LUT_AMPL_WIDTH),
		27116 => to_signed(16899, LUT_AMPL_WIDTH),
		27117 => to_signed(16897, LUT_AMPL_WIDTH),
		27118 => to_signed(16894, LUT_AMPL_WIDTH),
		27119 => to_signed(16891, LUT_AMPL_WIDTH),
		27120 => to_signed(16889, LUT_AMPL_WIDTH),
		27121 => to_signed(16886, LUT_AMPL_WIDTH),
		27122 => to_signed(16883, LUT_AMPL_WIDTH),
		27123 => to_signed(16881, LUT_AMPL_WIDTH),
		27124 => to_signed(16878, LUT_AMPL_WIDTH),
		27125 => to_signed(16875, LUT_AMPL_WIDTH),
		27126 => to_signed(16873, LUT_AMPL_WIDTH),
		27127 => to_signed(16870, LUT_AMPL_WIDTH),
		27128 => to_signed(16867, LUT_AMPL_WIDTH),
		27129 => to_signed(16864, LUT_AMPL_WIDTH),
		27130 => to_signed(16862, LUT_AMPL_WIDTH),
		27131 => to_signed(16859, LUT_AMPL_WIDTH),
		27132 => to_signed(16856, LUT_AMPL_WIDTH),
		27133 => to_signed(16854, LUT_AMPL_WIDTH),
		27134 => to_signed(16851, LUT_AMPL_WIDTH),
		27135 => to_signed(16848, LUT_AMPL_WIDTH),
		27136 => to_signed(16846, LUT_AMPL_WIDTH),
		27137 => to_signed(16843, LUT_AMPL_WIDTH),
		27138 => to_signed(16840, LUT_AMPL_WIDTH),
		27139 => to_signed(16838, LUT_AMPL_WIDTH),
		27140 => to_signed(16835, LUT_AMPL_WIDTH),
		27141 => to_signed(16832, LUT_AMPL_WIDTH),
		27142 => to_signed(16829, LUT_AMPL_WIDTH),
		27143 => to_signed(16827, LUT_AMPL_WIDTH),
		27144 => to_signed(16824, LUT_AMPL_WIDTH),
		27145 => to_signed(16821, LUT_AMPL_WIDTH),
		27146 => to_signed(16819, LUT_AMPL_WIDTH),
		27147 => to_signed(16816, LUT_AMPL_WIDTH),
		27148 => to_signed(16813, LUT_AMPL_WIDTH),
		27149 => to_signed(16811, LUT_AMPL_WIDTH),
		27150 => to_signed(16808, LUT_AMPL_WIDTH),
		27151 => to_signed(16805, LUT_AMPL_WIDTH),
		27152 => to_signed(16802, LUT_AMPL_WIDTH),
		27153 => to_signed(16800, LUT_AMPL_WIDTH),
		27154 => to_signed(16797, LUT_AMPL_WIDTH),
		27155 => to_signed(16794, LUT_AMPL_WIDTH),
		27156 => to_signed(16792, LUT_AMPL_WIDTH),
		27157 => to_signed(16789, LUT_AMPL_WIDTH),
		27158 => to_signed(16786, LUT_AMPL_WIDTH),
		27159 => to_signed(16784, LUT_AMPL_WIDTH),
		27160 => to_signed(16781, LUT_AMPL_WIDTH),
		27161 => to_signed(16778, LUT_AMPL_WIDTH),
		27162 => to_signed(16775, LUT_AMPL_WIDTH),
		27163 => to_signed(16773, LUT_AMPL_WIDTH),
		27164 => to_signed(16770, LUT_AMPL_WIDTH),
		27165 => to_signed(16767, LUT_AMPL_WIDTH),
		27166 => to_signed(16765, LUT_AMPL_WIDTH),
		27167 => to_signed(16762, LUT_AMPL_WIDTH),
		27168 => to_signed(16759, LUT_AMPL_WIDTH),
		27169 => to_signed(16757, LUT_AMPL_WIDTH),
		27170 => to_signed(16754, LUT_AMPL_WIDTH),
		27171 => to_signed(16751, LUT_AMPL_WIDTH),
		27172 => to_signed(16749, LUT_AMPL_WIDTH),
		27173 => to_signed(16746, LUT_AMPL_WIDTH),
		27174 => to_signed(16743, LUT_AMPL_WIDTH),
		27175 => to_signed(16740, LUT_AMPL_WIDTH),
		27176 => to_signed(16738, LUT_AMPL_WIDTH),
		27177 => to_signed(16735, LUT_AMPL_WIDTH),
		27178 => to_signed(16732, LUT_AMPL_WIDTH),
		27179 => to_signed(16730, LUT_AMPL_WIDTH),
		27180 => to_signed(16727, LUT_AMPL_WIDTH),
		27181 => to_signed(16724, LUT_AMPL_WIDTH),
		27182 => to_signed(16721, LUT_AMPL_WIDTH),
		27183 => to_signed(16719, LUT_AMPL_WIDTH),
		27184 => to_signed(16716, LUT_AMPL_WIDTH),
		27185 => to_signed(16713, LUT_AMPL_WIDTH),
		27186 => to_signed(16711, LUT_AMPL_WIDTH),
		27187 => to_signed(16708, LUT_AMPL_WIDTH),
		27188 => to_signed(16705, LUT_AMPL_WIDTH),
		27189 => to_signed(16703, LUT_AMPL_WIDTH),
		27190 => to_signed(16700, LUT_AMPL_WIDTH),
		27191 => to_signed(16697, LUT_AMPL_WIDTH),
		27192 => to_signed(16694, LUT_AMPL_WIDTH),
		27193 => to_signed(16692, LUT_AMPL_WIDTH),
		27194 => to_signed(16689, LUT_AMPL_WIDTH),
		27195 => to_signed(16686, LUT_AMPL_WIDTH),
		27196 => to_signed(16684, LUT_AMPL_WIDTH),
		27197 => to_signed(16681, LUT_AMPL_WIDTH),
		27198 => to_signed(16678, LUT_AMPL_WIDTH),
		27199 => to_signed(16676, LUT_AMPL_WIDTH),
		27200 => to_signed(16673, LUT_AMPL_WIDTH),
		27201 => to_signed(16670, LUT_AMPL_WIDTH),
		27202 => to_signed(16667, LUT_AMPL_WIDTH),
		27203 => to_signed(16665, LUT_AMPL_WIDTH),
		27204 => to_signed(16662, LUT_AMPL_WIDTH),
		27205 => to_signed(16659, LUT_AMPL_WIDTH),
		27206 => to_signed(16657, LUT_AMPL_WIDTH),
		27207 => to_signed(16654, LUT_AMPL_WIDTH),
		27208 => to_signed(16651, LUT_AMPL_WIDTH),
		27209 => to_signed(16648, LUT_AMPL_WIDTH),
		27210 => to_signed(16646, LUT_AMPL_WIDTH),
		27211 => to_signed(16643, LUT_AMPL_WIDTH),
		27212 => to_signed(16640, LUT_AMPL_WIDTH),
		27213 => to_signed(16638, LUT_AMPL_WIDTH),
		27214 => to_signed(16635, LUT_AMPL_WIDTH),
		27215 => to_signed(16632, LUT_AMPL_WIDTH),
		27216 => to_signed(16630, LUT_AMPL_WIDTH),
		27217 => to_signed(16627, LUT_AMPL_WIDTH),
		27218 => to_signed(16624, LUT_AMPL_WIDTH),
		27219 => to_signed(16621, LUT_AMPL_WIDTH),
		27220 => to_signed(16619, LUT_AMPL_WIDTH),
		27221 => to_signed(16616, LUT_AMPL_WIDTH),
		27222 => to_signed(16613, LUT_AMPL_WIDTH),
		27223 => to_signed(16611, LUT_AMPL_WIDTH),
		27224 => to_signed(16608, LUT_AMPL_WIDTH),
		27225 => to_signed(16605, LUT_AMPL_WIDTH),
		27226 => to_signed(16602, LUT_AMPL_WIDTH),
		27227 => to_signed(16600, LUT_AMPL_WIDTH),
		27228 => to_signed(16597, LUT_AMPL_WIDTH),
		27229 => to_signed(16594, LUT_AMPL_WIDTH),
		27230 => to_signed(16592, LUT_AMPL_WIDTH),
		27231 => to_signed(16589, LUT_AMPL_WIDTH),
		27232 => to_signed(16586, LUT_AMPL_WIDTH),
		27233 => to_signed(16584, LUT_AMPL_WIDTH),
		27234 => to_signed(16581, LUT_AMPL_WIDTH),
		27235 => to_signed(16578, LUT_AMPL_WIDTH),
		27236 => to_signed(16575, LUT_AMPL_WIDTH),
		27237 => to_signed(16573, LUT_AMPL_WIDTH),
		27238 => to_signed(16570, LUT_AMPL_WIDTH),
		27239 => to_signed(16567, LUT_AMPL_WIDTH),
		27240 => to_signed(16565, LUT_AMPL_WIDTH),
		27241 => to_signed(16562, LUT_AMPL_WIDTH),
		27242 => to_signed(16559, LUT_AMPL_WIDTH),
		27243 => to_signed(16556, LUT_AMPL_WIDTH),
		27244 => to_signed(16554, LUT_AMPL_WIDTH),
		27245 => to_signed(16551, LUT_AMPL_WIDTH),
		27246 => to_signed(16548, LUT_AMPL_WIDTH),
		27247 => to_signed(16546, LUT_AMPL_WIDTH),
		27248 => to_signed(16543, LUT_AMPL_WIDTH),
		27249 => to_signed(16540, LUT_AMPL_WIDTH),
		27250 => to_signed(16537, LUT_AMPL_WIDTH),
		27251 => to_signed(16535, LUT_AMPL_WIDTH),
		27252 => to_signed(16532, LUT_AMPL_WIDTH),
		27253 => to_signed(16529, LUT_AMPL_WIDTH),
		27254 => to_signed(16527, LUT_AMPL_WIDTH),
		27255 => to_signed(16524, LUT_AMPL_WIDTH),
		27256 => to_signed(16521, LUT_AMPL_WIDTH),
		27257 => to_signed(16518, LUT_AMPL_WIDTH),
		27258 => to_signed(16516, LUT_AMPL_WIDTH),
		27259 => to_signed(16513, LUT_AMPL_WIDTH),
		27260 => to_signed(16510, LUT_AMPL_WIDTH),
		27261 => to_signed(16508, LUT_AMPL_WIDTH),
		27262 => to_signed(16505, LUT_AMPL_WIDTH),
		27263 => to_signed(16502, LUT_AMPL_WIDTH),
		27264 => to_signed(16499, LUT_AMPL_WIDTH),
		27265 => to_signed(16497, LUT_AMPL_WIDTH),
		27266 => to_signed(16494, LUT_AMPL_WIDTH),
		27267 => to_signed(16491, LUT_AMPL_WIDTH),
		27268 => to_signed(16489, LUT_AMPL_WIDTH),
		27269 => to_signed(16486, LUT_AMPL_WIDTH),
		27270 => to_signed(16483, LUT_AMPL_WIDTH),
		27271 => to_signed(16480, LUT_AMPL_WIDTH),
		27272 => to_signed(16478, LUT_AMPL_WIDTH),
		27273 => to_signed(16475, LUT_AMPL_WIDTH),
		27274 => to_signed(16472, LUT_AMPL_WIDTH),
		27275 => to_signed(16470, LUT_AMPL_WIDTH),
		27276 => to_signed(16467, LUT_AMPL_WIDTH),
		27277 => to_signed(16464, LUT_AMPL_WIDTH),
		27278 => to_signed(16461, LUT_AMPL_WIDTH),
		27279 => to_signed(16459, LUT_AMPL_WIDTH),
		27280 => to_signed(16456, LUT_AMPL_WIDTH),
		27281 => to_signed(16453, LUT_AMPL_WIDTH),
		27282 => to_signed(16451, LUT_AMPL_WIDTH),
		27283 => to_signed(16448, LUT_AMPL_WIDTH),
		27284 => to_signed(16445, LUT_AMPL_WIDTH),
		27285 => to_signed(16442, LUT_AMPL_WIDTH),
		27286 => to_signed(16440, LUT_AMPL_WIDTH),
		27287 => to_signed(16437, LUT_AMPL_WIDTH),
		27288 => to_signed(16434, LUT_AMPL_WIDTH),
		27289 => to_signed(16432, LUT_AMPL_WIDTH),
		27290 => to_signed(16429, LUT_AMPL_WIDTH),
		27291 => to_signed(16426, LUT_AMPL_WIDTH),
		27292 => to_signed(16423, LUT_AMPL_WIDTH),
		27293 => to_signed(16421, LUT_AMPL_WIDTH),
		27294 => to_signed(16418, LUT_AMPL_WIDTH),
		27295 => to_signed(16415, LUT_AMPL_WIDTH),
		27296 => to_signed(16413, LUT_AMPL_WIDTH),
		27297 => to_signed(16410, LUT_AMPL_WIDTH),
		27298 => to_signed(16407, LUT_AMPL_WIDTH),
		27299 => to_signed(16404, LUT_AMPL_WIDTH),
		27300 => to_signed(16402, LUT_AMPL_WIDTH),
		27301 => to_signed(16399, LUT_AMPL_WIDTH),
		27302 => to_signed(16396, LUT_AMPL_WIDTH),
		27303 => to_signed(16393, LUT_AMPL_WIDTH),
		27304 => to_signed(16391, LUT_AMPL_WIDTH),
		27305 => to_signed(16388, LUT_AMPL_WIDTH),
		27306 => to_signed(16385, LUT_AMPL_WIDTH),
		27307 => to_signed(16383, LUT_AMPL_WIDTH),
		27308 => to_signed(16380, LUT_AMPL_WIDTH),
		27309 => to_signed(16377, LUT_AMPL_WIDTH),
		27310 => to_signed(16374, LUT_AMPL_WIDTH),
		27311 => to_signed(16372, LUT_AMPL_WIDTH),
		27312 => to_signed(16369, LUT_AMPL_WIDTH),
		27313 => to_signed(16366, LUT_AMPL_WIDTH),
		27314 => to_signed(16364, LUT_AMPL_WIDTH),
		27315 => to_signed(16361, LUT_AMPL_WIDTH),
		27316 => to_signed(16358, LUT_AMPL_WIDTH),
		27317 => to_signed(16355, LUT_AMPL_WIDTH),
		27318 => to_signed(16353, LUT_AMPL_WIDTH),
		27319 => to_signed(16350, LUT_AMPL_WIDTH),
		27320 => to_signed(16347, LUT_AMPL_WIDTH),
		27321 => to_signed(16344, LUT_AMPL_WIDTH),
		27322 => to_signed(16342, LUT_AMPL_WIDTH),
		27323 => to_signed(16339, LUT_AMPL_WIDTH),
		27324 => to_signed(16336, LUT_AMPL_WIDTH),
		27325 => to_signed(16334, LUT_AMPL_WIDTH),
		27326 => to_signed(16331, LUT_AMPL_WIDTH),
		27327 => to_signed(16328, LUT_AMPL_WIDTH),
		27328 => to_signed(16325, LUT_AMPL_WIDTH),
		27329 => to_signed(16323, LUT_AMPL_WIDTH),
		27330 => to_signed(16320, LUT_AMPL_WIDTH),
		27331 => to_signed(16317, LUT_AMPL_WIDTH),
		27332 => to_signed(16315, LUT_AMPL_WIDTH),
		27333 => to_signed(16312, LUT_AMPL_WIDTH),
		27334 => to_signed(16309, LUT_AMPL_WIDTH),
		27335 => to_signed(16306, LUT_AMPL_WIDTH),
		27336 => to_signed(16304, LUT_AMPL_WIDTH),
		27337 => to_signed(16301, LUT_AMPL_WIDTH),
		27338 => to_signed(16298, LUT_AMPL_WIDTH),
		27339 => to_signed(16295, LUT_AMPL_WIDTH),
		27340 => to_signed(16293, LUT_AMPL_WIDTH),
		27341 => to_signed(16290, LUT_AMPL_WIDTH),
		27342 => to_signed(16287, LUT_AMPL_WIDTH),
		27343 => to_signed(16285, LUT_AMPL_WIDTH),
		27344 => to_signed(16282, LUT_AMPL_WIDTH),
		27345 => to_signed(16279, LUT_AMPL_WIDTH),
		27346 => to_signed(16276, LUT_AMPL_WIDTH),
		27347 => to_signed(16274, LUT_AMPL_WIDTH),
		27348 => to_signed(16271, LUT_AMPL_WIDTH),
		27349 => to_signed(16268, LUT_AMPL_WIDTH),
		27350 => to_signed(16265, LUT_AMPL_WIDTH),
		27351 => to_signed(16263, LUT_AMPL_WIDTH),
		27352 => to_signed(16260, LUT_AMPL_WIDTH),
		27353 => to_signed(16257, LUT_AMPL_WIDTH),
		27354 => to_signed(16255, LUT_AMPL_WIDTH),
		27355 => to_signed(16252, LUT_AMPL_WIDTH),
		27356 => to_signed(16249, LUT_AMPL_WIDTH),
		27357 => to_signed(16246, LUT_AMPL_WIDTH),
		27358 => to_signed(16244, LUT_AMPL_WIDTH),
		27359 => to_signed(16241, LUT_AMPL_WIDTH),
		27360 => to_signed(16238, LUT_AMPL_WIDTH),
		27361 => to_signed(16235, LUT_AMPL_WIDTH),
		27362 => to_signed(16233, LUT_AMPL_WIDTH),
		27363 => to_signed(16230, LUT_AMPL_WIDTH),
		27364 => to_signed(16227, LUT_AMPL_WIDTH),
		27365 => to_signed(16225, LUT_AMPL_WIDTH),
		27366 => to_signed(16222, LUT_AMPL_WIDTH),
		27367 => to_signed(16219, LUT_AMPL_WIDTH),
		27368 => to_signed(16216, LUT_AMPL_WIDTH),
		27369 => to_signed(16214, LUT_AMPL_WIDTH),
		27370 => to_signed(16211, LUT_AMPL_WIDTH),
		27371 => to_signed(16208, LUT_AMPL_WIDTH),
		27372 => to_signed(16205, LUT_AMPL_WIDTH),
		27373 => to_signed(16203, LUT_AMPL_WIDTH),
		27374 => to_signed(16200, LUT_AMPL_WIDTH),
		27375 => to_signed(16197, LUT_AMPL_WIDTH),
		27376 => to_signed(16195, LUT_AMPL_WIDTH),
		27377 => to_signed(16192, LUT_AMPL_WIDTH),
		27378 => to_signed(16189, LUT_AMPL_WIDTH),
		27379 => to_signed(16186, LUT_AMPL_WIDTH),
		27380 => to_signed(16184, LUT_AMPL_WIDTH),
		27381 => to_signed(16181, LUT_AMPL_WIDTH),
		27382 => to_signed(16178, LUT_AMPL_WIDTH),
		27383 => to_signed(16175, LUT_AMPL_WIDTH),
		27384 => to_signed(16173, LUT_AMPL_WIDTH),
		27385 => to_signed(16170, LUT_AMPL_WIDTH),
		27386 => to_signed(16167, LUT_AMPL_WIDTH),
		27387 => to_signed(16164, LUT_AMPL_WIDTH),
		27388 => to_signed(16162, LUT_AMPL_WIDTH),
		27389 => to_signed(16159, LUT_AMPL_WIDTH),
		27390 => to_signed(16156, LUT_AMPL_WIDTH),
		27391 => to_signed(16154, LUT_AMPL_WIDTH),
		27392 => to_signed(16151, LUT_AMPL_WIDTH),
		27393 => to_signed(16148, LUT_AMPL_WIDTH),
		27394 => to_signed(16145, LUT_AMPL_WIDTH),
		27395 => to_signed(16143, LUT_AMPL_WIDTH),
		27396 => to_signed(16140, LUT_AMPL_WIDTH),
		27397 => to_signed(16137, LUT_AMPL_WIDTH),
		27398 => to_signed(16134, LUT_AMPL_WIDTH),
		27399 => to_signed(16132, LUT_AMPL_WIDTH),
		27400 => to_signed(16129, LUT_AMPL_WIDTH),
		27401 => to_signed(16126, LUT_AMPL_WIDTH),
		27402 => to_signed(16123, LUT_AMPL_WIDTH),
		27403 => to_signed(16121, LUT_AMPL_WIDTH),
		27404 => to_signed(16118, LUT_AMPL_WIDTH),
		27405 => to_signed(16115, LUT_AMPL_WIDTH),
		27406 => to_signed(16113, LUT_AMPL_WIDTH),
		27407 => to_signed(16110, LUT_AMPL_WIDTH),
		27408 => to_signed(16107, LUT_AMPL_WIDTH),
		27409 => to_signed(16104, LUT_AMPL_WIDTH),
		27410 => to_signed(16102, LUT_AMPL_WIDTH),
		27411 => to_signed(16099, LUT_AMPL_WIDTH),
		27412 => to_signed(16096, LUT_AMPL_WIDTH),
		27413 => to_signed(16093, LUT_AMPL_WIDTH),
		27414 => to_signed(16091, LUT_AMPL_WIDTH),
		27415 => to_signed(16088, LUT_AMPL_WIDTH),
		27416 => to_signed(16085, LUT_AMPL_WIDTH),
		27417 => to_signed(16082, LUT_AMPL_WIDTH),
		27418 => to_signed(16080, LUT_AMPL_WIDTH),
		27419 => to_signed(16077, LUT_AMPL_WIDTH),
		27420 => to_signed(16074, LUT_AMPL_WIDTH),
		27421 => to_signed(16071, LUT_AMPL_WIDTH),
		27422 => to_signed(16069, LUT_AMPL_WIDTH),
		27423 => to_signed(16066, LUT_AMPL_WIDTH),
		27424 => to_signed(16063, LUT_AMPL_WIDTH),
		27425 => to_signed(16061, LUT_AMPL_WIDTH),
		27426 => to_signed(16058, LUT_AMPL_WIDTH),
		27427 => to_signed(16055, LUT_AMPL_WIDTH),
		27428 => to_signed(16052, LUT_AMPL_WIDTH),
		27429 => to_signed(16050, LUT_AMPL_WIDTH),
		27430 => to_signed(16047, LUT_AMPL_WIDTH),
		27431 => to_signed(16044, LUT_AMPL_WIDTH),
		27432 => to_signed(16041, LUT_AMPL_WIDTH),
		27433 => to_signed(16039, LUT_AMPL_WIDTH),
		27434 => to_signed(16036, LUT_AMPL_WIDTH),
		27435 => to_signed(16033, LUT_AMPL_WIDTH),
		27436 => to_signed(16030, LUT_AMPL_WIDTH),
		27437 => to_signed(16028, LUT_AMPL_WIDTH),
		27438 => to_signed(16025, LUT_AMPL_WIDTH),
		27439 => to_signed(16022, LUT_AMPL_WIDTH),
		27440 => to_signed(16019, LUT_AMPL_WIDTH),
		27441 => to_signed(16017, LUT_AMPL_WIDTH),
		27442 => to_signed(16014, LUT_AMPL_WIDTH),
		27443 => to_signed(16011, LUT_AMPL_WIDTH),
		27444 => to_signed(16008, LUT_AMPL_WIDTH),
		27445 => to_signed(16006, LUT_AMPL_WIDTH),
		27446 => to_signed(16003, LUT_AMPL_WIDTH),
		27447 => to_signed(16000, LUT_AMPL_WIDTH),
		27448 => to_signed(15997, LUT_AMPL_WIDTH),
		27449 => to_signed(15995, LUT_AMPL_WIDTH),
		27450 => to_signed(15992, LUT_AMPL_WIDTH),
		27451 => to_signed(15989, LUT_AMPL_WIDTH),
		27452 => to_signed(15987, LUT_AMPL_WIDTH),
		27453 => to_signed(15984, LUT_AMPL_WIDTH),
		27454 => to_signed(15981, LUT_AMPL_WIDTH),
		27455 => to_signed(15978, LUT_AMPL_WIDTH),
		27456 => to_signed(15976, LUT_AMPL_WIDTH),
		27457 => to_signed(15973, LUT_AMPL_WIDTH),
		27458 => to_signed(15970, LUT_AMPL_WIDTH),
		27459 => to_signed(15967, LUT_AMPL_WIDTH),
		27460 => to_signed(15965, LUT_AMPL_WIDTH),
		27461 => to_signed(15962, LUT_AMPL_WIDTH),
		27462 => to_signed(15959, LUT_AMPL_WIDTH),
		27463 => to_signed(15956, LUT_AMPL_WIDTH),
		27464 => to_signed(15954, LUT_AMPL_WIDTH),
		27465 => to_signed(15951, LUT_AMPL_WIDTH),
		27466 => to_signed(15948, LUT_AMPL_WIDTH),
		27467 => to_signed(15945, LUT_AMPL_WIDTH),
		27468 => to_signed(15943, LUT_AMPL_WIDTH),
		27469 => to_signed(15940, LUT_AMPL_WIDTH),
		27470 => to_signed(15937, LUT_AMPL_WIDTH),
		27471 => to_signed(15934, LUT_AMPL_WIDTH),
		27472 => to_signed(15932, LUT_AMPL_WIDTH),
		27473 => to_signed(15929, LUT_AMPL_WIDTH),
		27474 => to_signed(15926, LUT_AMPL_WIDTH),
		27475 => to_signed(15923, LUT_AMPL_WIDTH),
		27476 => to_signed(15921, LUT_AMPL_WIDTH),
		27477 => to_signed(15918, LUT_AMPL_WIDTH),
		27478 => to_signed(15915, LUT_AMPL_WIDTH),
		27479 => to_signed(15912, LUT_AMPL_WIDTH),
		27480 => to_signed(15910, LUT_AMPL_WIDTH),
		27481 => to_signed(15907, LUT_AMPL_WIDTH),
		27482 => to_signed(15904, LUT_AMPL_WIDTH),
		27483 => to_signed(15901, LUT_AMPL_WIDTH),
		27484 => to_signed(15899, LUT_AMPL_WIDTH),
		27485 => to_signed(15896, LUT_AMPL_WIDTH),
		27486 => to_signed(15893, LUT_AMPL_WIDTH),
		27487 => to_signed(15890, LUT_AMPL_WIDTH),
		27488 => to_signed(15888, LUT_AMPL_WIDTH),
		27489 => to_signed(15885, LUT_AMPL_WIDTH),
		27490 => to_signed(15882, LUT_AMPL_WIDTH),
		27491 => to_signed(15879, LUT_AMPL_WIDTH),
		27492 => to_signed(15877, LUT_AMPL_WIDTH),
		27493 => to_signed(15874, LUT_AMPL_WIDTH),
		27494 => to_signed(15871, LUT_AMPL_WIDTH),
		27495 => to_signed(15868, LUT_AMPL_WIDTH),
		27496 => to_signed(15866, LUT_AMPL_WIDTH),
		27497 => to_signed(15863, LUT_AMPL_WIDTH),
		27498 => to_signed(15860, LUT_AMPL_WIDTH),
		27499 => to_signed(15857, LUT_AMPL_WIDTH),
		27500 => to_signed(15855, LUT_AMPL_WIDTH),
		27501 => to_signed(15852, LUT_AMPL_WIDTH),
		27502 => to_signed(15849, LUT_AMPL_WIDTH),
		27503 => to_signed(15846, LUT_AMPL_WIDTH),
		27504 => to_signed(15844, LUT_AMPL_WIDTH),
		27505 => to_signed(15841, LUT_AMPL_WIDTH),
		27506 => to_signed(15838, LUT_AMPL_WIDTH),
		27507 => to_signed(15835, LUT_AMPL_WIDTH),
		27508 => to_signed(15833, LUT_AMPL_WIDTH),
		27509 => to_signed(15830, LUT_AMPL_WIDTH),
		27510 => to_signed(15827, LUT_AMPL_WIDTH),
		27511 => to_signed(15824, LUT_AMPL_WIDTH),
		27512 => to_signed(15822, LUT_AMPL_WIDTH),
		27513 => to_signed(15819, LUT_AMPL_WIDTH),
		27514 => to_signed(15816, LUT_AMPL_WIDTH),
		27515 => to_signed(15813, LUT_AMPL_WIDTH),
		27516 => to_signed(15811, LUT_AMPL_WIDTH),
		27517 => to_signed(15808, LUT_AMPL_WIDTH),
		27518 => to_signed(15805, LUT_AMPL_WIDTH),
		27519 => to_signed(15802, LUT_AMPL_WIDTH),
		27520 => to_signed(15800, LUT_AMPL_WIDTH),
		27521 => to_signed(15797, LUT_AMPL_WIDTH),
		27522 => to_signed(15794, LUT_AMPL_WIDTH),
		27523 => to_signed(15791, LUT_AMPL_WIDTH),
		27524 => to_signed(15789, LUT_AMPL_WIDTH),
		27525 => to_signed(15786, LUT_AMPL_WIDTH),
		27526 => to_signed(15783, LUT_AMPL_WIDTH),
		27527 => to_signed(15780, LUT_AMPL_WIDTH),
		27528 => to_signed(15778, LUT_AMPL_WIDTH),
		27529 => to_signed(15775, LUT_AMPL_WIDTH),
		27530 => to_signed(15772, LUT_AMPL_WIDTH),
		27531 => to_signed(15769, LUT_AMPL_WIDTH),
		27532 => to_signed(15767, LUT_AMPL_WIDTH),
		27533 => to_signed(15764, LUT_AMPL_WIDTH),
		27534 => to_signed(15761, LUT_AMPL_WIDTH),
		27535 => to_signed(15758, LUT_AMPL_WIDTH),
		27536 => to_signed(15756, LUT_AMPL_WIDTH),
		27537 => to_signed(15753, LUT_AMPL_WIDTH),
		27538 => to_signed(15750, LUT_AMPL_WIDTH),
		27539 => to_signed(15747, LUT_AMPL_WIDTH),
		27540 => to_signed(15745, LUT_AMPL_WIDTH),
		27541 => to_signed(15742, LUT_AMPL_WIDTH),
		27542 => to_signed(15739, LUT_AMPL_WIDTH),
		27543 => to_signed(15736, LUT_AMPL_WIDTH),
		27544 => to_signed(15734, LUT_AMPL_WIDTH),
		27545 => to_signed(15731, LUT_AMPL_WIDTH),
		27546 => to_signed(15728, LUT_AMPL_WIDTH),
		27547 => to_signed(15725, LUT_AMPL_WIDTH),
		27548 => to_signed(15723, LUT_AMPL_WIDTH),
		27549 => to_signed(15720, LUT_AMPL_WIDTH),
		27550 => to_signed(15717, LUT_AMPL_WIDTH),
		27551 => to_signed(15714, LUT_AMPL_WIDTH),
		27552 => to_signed(15712, LUT_AMPL_WIDTH),
		27553 => to_signed(15709, LUT_AMPL_WIDTH),
		27554 => to_signed(15706, LUT_AMPL_WIDTH),
		27555 => to_signed(15703, LUT_AMPL_WIDTH),
		27556 => to_signed(15701, LUT_AMPL_WIDTH),
		27557 => to_signed(15698, LUT_AMPL_WIDTH),
		27558 => to_signed(15695, LUT_AMPL_WIDTH),
		27559 => to_signed(15692, LUT_AMPL_WIDTH),
		27560 => to_signed(15690, LUT_AMPL_WIDTH),
		27561 => to_signed(15687, LUT_AMPL_WIDTH),
		27562 => to_signed(15684, LUT_AMPL_WIDTH),
		27563 => to_signed(15681, LUT_AMPL_WIDTH),
		27564 => to_signed(15678, LUT_AMPL_WIDTH),
		27565 => to_signed(15676, LUT_AMPL_WIDTH),
		27566 => to_signed(15673, LUT_AMPL_WIDTH),
		27567 => to_signed(15670, LUT_AMPL_WIDTH),
		27568 => to_signed(15667, LUT_AMPL_WIDTH),
		27569 => to_signed(15665, LUT_AMPL_WIDTH),
		27570 => to_signed(15662, LUT_AMPL_WIDTH),
		27571 => to_signed(15659, LUT_AMPL_WIDTH),
		27572 => to_signed(15656, LUT_AMPL_WIDTH),
		27573 => to_signed(15654, LUT_AMPL_WIDTH),
		27574 => to_signed(15651, LUT_AMPL_WIDTH),
		27575 => to_signed(15648, LUT_AMPL_WIDTH),
		27576 => to_signed(15645, LUT_AMPL_WIDTH),
		27577 => to_signed(15643, LUT_AMPL_WIDTH),
		27578 => to_signed(15640, LUT_AMPL_WIDTH),
		27579 => to_signed(15637, LUT_AMPL_WIDTH),
		27580 => to_signed(15634, LUT_AMPL_WIDTH),
		27581 => to_signed(15632, LUT_AMPL_WIDTH),
		27582 => to_signed(15629, LUT_AMPL_WIDTH),
		27583 => to_signed(15626, LUT_AMPL_WIDTH),
		27584 => to_signed(15623, LUT_AMPL_WIDTH),
		27585 => to_signed(15621, LUT_AMPL_WIDTH),
		27586 => to_signed(15618, LUT_AMPL_WIDTH),
		27587 => to_signed(15615, LUT_AMPL_WIDTH),
		27588 => to_signed(15612, LUT_AMPL_WIDTH),
		27589 => to_signed(15609, LUT_AMPL_WIDTH),
		27590 => to_signed(15607, LUT_AMPL_WIDTH),
		27591 => to_signed(15604, LUT_AMPL_WIDTH),
		27592 => to_signed(15601, LUT_AMPL_WIDTH),
		27593 => to_signed(15598, LUT_AMPL_WIDTH),
		27594 => to_signed(15596, LUT_AMPL_WIDTH),
		27595 => to_signed(15593, LUT_AMPL_WIDTH),
		27596 => to_signed(15590, LUT_AMPL_WIDTH),
		27597 => to_signed(15587, LUT_AMPL_WIDTH),
		27598 => to_signed(15585, LUT_AMPL_WIDTH),
		27599 => to_signed(15582, LUT_AMPL_WIDTH),
		27600 => to_signed(15579, LUT_AMPL_WIDTH),
		27601 => to_signed(15576, LUT_AMPL_WIDTH),
		27602 => to_signed(15574, LUT_AMPL_WIDTH),
		27603 => to_signed(15571, LUT_AMPL_WIDTH),
		27604 => to_signed(15568, LUT_AMPL_WIDTH),
		27605 => to_signed(15565, LUT_AMPL_WIDTH),
		27606 => to_signed(15562, LUT_AMPL_WIDTH),
		27607 => to_signed(15560, LUT_AMPL_WIDTH),
		27608 => to_signed(15557, LUT_AMPL_WIDTH),
		27609 => to_signed(15554, LUT_AMPL_WIDTH),
		27610 => to_signed(15551, LUT_AMPL_WIDTH),
		27611 => to_signed(15549, LUT_AMPL_WIDTH),
		27612 => to_signed(15546, LUT_AMPL_WIDTH),
		27613 => to_signed(15543, LUT_AMPL_WIDTH),
		27614 => to_signed(15540, LUT_AMPL_WIDTH),
		27615 => to_signed(15538, LUT_AMPL_WIDTH),
		27616 => to_signed(15535, LUT_AMPL_WIDTH),
		27617 => to_signed(15532, LUT_AMPL_WIDTH),
		27618 => to_signed(15529, LUT_AMPL_WIDTH),
		27619 => to_signed(15527, LUT_AMPL_WIDTH),
		27620 => to_signed(15524, LUT_AMPL_WIDTH),
		27621 => to_signed(15521, LUT_AMPL_WIDTH),
		27622 => to_signed(15518, LUT_AMPL_WIDTH),
		27623 => to_signed(15515, LUT_AMPL_WIDTH),
		27624 => to_signed(15513, LUT_AMPL_WIDTH),
		27625 => to_signed(15510, LUT_AMPL_WIDTH),
		27626 => to_signed(15507, LUT_AMPL_WIDTH),
		27627 => to_signed(15504, LUT_AMPL_WIDTH),
		27628 => to_signed(15502, LUT_AMPL_WIDTH),
		27629 => to_signed(15499, LUT_AMPL_WIDTH),
		27630 => to_signed(15496, LUT_AMPL_WIDTH),
		27631 => to_signed(15493, LUT_AMPL_WIDTH),
		27632 => to_signed(15491, LUT_AMPL_WIDTH),
		27633 => to_signed(15488, LUT_AMPL_WIDTH),
		27634 => to_signed(15485, LUT_AMPL_WIDTH),
		27635 => to_signed(15482, LUT_AMPL_WIDTH),
		27636 => to_signed(15479, LUT_AMPL_WIDTH),
		27637 => to_signed(15477, LUT_AMPL_WIDTH),
		27638 => to_signed(15474, LUT_AMPL_WIDTH),
		27639 => to_signed(15471, LUT_AMPL_WIDTH),
		27640 => to_signed(15468, LUT_AMPL_WIDTH),
		27641 => to_signed(15466, LUT_AMPL_WIDTH),
		27642 => to_signed(15463, LUT_AMPL_WIDTH),
		27643 => to_signed(15460, LUT_AMPL_WIDTH),
		27644 => to_signed(15457, LUT_AMPL_WIDTH),
		27645 => to_signed(15455, LUT_AMPL_WIDTH),
		27646 => to_signed(15452, LUT_AMPL_WIDTH),
		27647 => to_signed(15449, LUT_AMPL_WIDTH),
		27648 => to_signed(15446, LUT_AMPL_WIDTH),
		27649 => to_signed(15443, LUT_AMPL_WIDTH),
		27650 => to_signed(15441, LUT_AMPL_WIDTH),
		27651 => to_signed(15438, LUT_AMPL_WIDTH),
		27652 => to_signed(15435, LUT_AMPL_WIDTH),
		27653 => to_signed(15432, LUT_AMPL_WIDTH),
		27654 => to_signed(15430, LUT_AMPL_WIDTH),
		27655 => to_signed(15427, LUT_AMPL_WIDTH),
		27656 => to_signed(15424, LUT_AMPL_WIDTH),
		27657 => to_signed(15421, LUT_AMPL_WIDTH),
		27658 => to_signed(15419, LUT_AMPL_WIDTH),
		27659 => to_signed(15416, LUT_AMPL_WIDTH),
		27660 => to_signed(15413, LUT_AMPL_WIDTH),
		27661 => to_signed(15410, LUT_AMPL_WIDTH),
		27662 => to_signed(15407, LUT_AMPL_WIDTH),
		27663 => to_signed(15405, LUT_AMPL_WIDTH),
		27664 => to_signed(15402, LUT_AMPL_WIDTH),
		27665 => to_signed(15399, LUT_AMPL_WIDTH),
		27666 => to_signed(15396, LUT_AMPL_WIDTH),
		27667 => to_signed(15394, LUT_AMPL_WIDTH),
		27668 => to_signed(15391, LUT_AMPL_WIDTH),
		27669 => to_signed(15388, LUT_AMPL_WIDTH),
		27670 => to_signed(15385, LUT_AMPL_WIDTH),
		27671 => to_signed(15382, LUT_AMPL_WIDTH),
		27672 => to_signed(15380, LUT_AMPL_WIDTH),
		27673 => to_signed(15377, LUT_AMPL_WIDTH),
		27674 => to_signed(15374, LUT_AMPL_WIDTH),
		27675 => to_signed(15371, LUT_AMPL_WIDTH),
		27676 => to_signed(15369, LUT_AMPL_WIDTH),
		27677 => to_signed(15366, LUT_AMPL_WIDTH),
		27678 => to_signed(15363, LUT_AMPL_WIDTH),
		27679 => to_signed(15360, LUT_AMPL_WIDTH),
		27680 => to_signed(15358, LUT_AMPL_WIDTH),
		27681 => to_signed(15355, LUT_AMPL_WIDTH),
		27682 => to_signed(15352, LUT_AMPL_WIDTH),
		27683 => to_signed(15349, LUT_AMPL_WIDTH),
		27684 => to_signed(15346, LUT_AMPL_WIDTH),
		27685 => to_signed(15344, LUT_AMPL_WIDTH),
		27686 => to_signed(15341, LUT_AMPL_WIDTH),
		27687 => to_signed(15338, LUT_AMPL_WIDTH),
		27688 => to_signed(15335, LUT_AMPL_WIDTH),
		27689 => to_signed(15333, LUT_AMPL_WIDTH),
		27690 => to_signed(15330, LUT_AMPL_WIDTH),
		27691 => to_signed(15327, LUT_AMPL_WIDTH),
		27692 => to_signed(15324, LUT_AMPL_WIDTH),
		27693 => to_signed(15321, LUT_AMPL_WIDTH),
		27694 => to_signed(15319, LUT_AMPL_WIDTH),
		27695 => to_signed(15316, LUT_AMPL_WIDTH),
		27696 => to_signed(15313, LUT_AMPL_WIDTH),
		27697 => to_signed(15310, LUT_AMPL_WIDTH),
		27698 => to_signed(15308, LUT_AMPL_WIDTH),
		27699 => to_signed(15305, LUT_AMPL_WIDTH),
		27700 => to_signed(15302, LUT_AMPL_WIDTH),
		27701 => to_signed(15299, LUT_AMPL_WIDTH),
		27702 => to_signed(15296, LUT_AMPL_WIDTH),
		27703 => to_signed(15294, LUT_AMPL_WIDTH),
		27704 => to_signed(15291, LUT_AMPL_WIDTH),
		27705 => to_signed(15288, LUT_AMPL_WIDTH),
		27706 => to_signed(15285, LUT_AMPL_WIDTH),
		27707 => to_signed(15283, LUT_AMPL_WIDTH),
		27708 => to_signed(15280, LUT_AMPL_WIDTH),
		27709 => to_signed(15277, LUT_AMPL_WIDTH),
		27710 => to_signed(15274, LUT_AMPL_WIDTH),
		27711 => to_signed(15271, LUT_AMPL_WIDTH),
		27712 => to_signed(15269, LUT_AMPL_WIDTH),
		27713 => to_signed(15266, LUT_AMPL_WIDTH),
		27714 => to_signed(15263, LUT_AMPL_WIDTH),
		27715 => to_signed(15260, LUT_AMPL_WIDTH),
		27716 => to_signed(15258, LUT_AMPL_WIDTH),
		27717 => to_signed(15255, LUT_AMPL_WIDTH),
		27718 => to_signed(15252, LUT_AMPL_WIDTH),
		27719 => to_signed(15249, LUT_AMPL_WIDTH),
		27720 => to_signed(15246, LUT_AMPL_WIDTH),
		27721 => to_signed(15244, LUT_AMPL_WIDTH),
		27722 => to_signed(15241, LUT_AMPL_WIDTH),
		27723 => to_signed(15238, LUT_AMPL_WIDTH),
		27724 => to_signed(15235, LUT_AMPL_WIDTH),
		27725 => to_signed(15233, LUT_AMPL_WIDTH),
		27726 => to_signed(15230, LUT_AMPL_WIDTH),
		27727 => to_signed(15227, LUT_AMPL_WIDTH),
		27728 => to_signed(15224, LUT_AMPL_WIDTH),
		27729 => to_signed(15221, LUT_AMPL_WIDTH),
		27730 => to_signed(15219, LUT_AMPL_WIDTH),
		27731 => to_signed(15216, LUT_AMPL_WIDTH),
		27732 => to_signed(15213, LUT_AMPL_WIDTH),
		27733 => to_signed(15210, LUT_AMPL_WIDTH),
		27734 => to_signed(15207, LUT_AMPL_WIDTH),
		27735 => to_signed(15205, LUT_AMPL_WIDTH),
		27736 => to_signed(15202, LUT_AMPL_WIDTH),
		27737 => to_signed(15199, LUT_AMPL_WIDTH),
		27738 => to_signed(15196, LUT_AMPL_WIDTH),
		27739 => to_signed(15194, LUT_AMPL_WIDTH),
		27740 => to_signed(15191, LUT_AMPL_WIDTH),
		27741 => to_signed(15188, LUT_AMPL_WIDTH),
		27742 => to_signed(15185, LUT_AMPL_WIDTH),
		27743 => to_signed(15182, LUT_AMPL_WIDTH),
		27744 => to_signed(15180, LUT_AMPL_WIDTH),
		27745 => to_signed(15177, LUT_AMPL_WIDTH),
		27746 => to_signed(15174, LUT_AMPL_WIDTH),
		27747 => to_signed(15171, LUT_AMPL_WIDTH),
		27748 => to_signed(15168, LUT_AMPL_WIDTH),
		27749 => to_signed(15166, LUT_AMPL_WIDTH),
		27750 => to_signed(15163, LUT_AMPL_WIDTH),
		27751 => to_signed(15160, LUT_AMPL_WIDTH),
		27752 => to_signed(15157, LUT_AMPL_WIDTH),
		27753 => to_signed(15155, LUT_AMPL_WIDTH),
		27754 => to_signed(15152, LUT_AMPL_WIDTH),
		27755 => to_signed(15149, LUT_AMPL_WIDTH),
		27756 => to_signed(15146, LUT_AMPL_WIDTH),
		27757 => to_signed(15143, LUT_AMPL_WIDTH),
		27758 => to_signed(15141, LUT_AMPL_WIDTH),
		27759 => to_signed(15138, LUT_AMPL_WIDTH),
		27760 => to_signed(15135, LUT_AMPL_WIDTH),
		27761 => to_signed(15132, LUT_AMPL_WIDTH),
		27762 => to_signed(15129, LUT_AMPL_WIDTH),
		27763 => to_signed(15127, LUT_AMPL_WIDTH),
		27764 => to_signed(15124, LUT_AMPL_WIDTH),
		27765 => to_signed(15121, LUT_AMPL_WIDTH),
		27766 => to_signed(15118, LUT_AMPL_WIDTH),
		27767 => to_signed(15116, LUT_AMPL_WIDTH),
		27768 => to_signed(15113, LUT_AMPL_WIDTH),
		27769 => to_signed(15110, LUT_AMPL_WIDTH),
		27770 => to_signed(15107, LUT_AMPL_WIDTH),
		27771 => to_signed(15104, LUT_AMPL_WIDTH),
		27772 => to_signed(15102, LUT_AMPL_WIDTH),
		27773 => to_signed(15099, LUT_AMPL_WIDTH),
		27774 => to_signed(15096, LUT_AMPL_WIDTH),
		27775 => to_signed(15093, LUT_AMPL_WIDTH),
		27776 => to_signed(15090, LUT_AMPL_WIDTH),
		27777 => to_signed(15088, LUT_AMPL_WIDTH),
		27778 => to_signed(15085, LUT_AMPL_WIDTH),
		27779 => to_signed(15082, LUT_AMPL_WIDTH),
		27780 => to_signed(15079, LUT_AMPL_WIDTH),
		27781 => to_signed(15077, LUT_AMPL_WIDTH),
		27782 => to_signed(15074, LUT_AMPL_WIDTH),
		27783 => to_signed(15071, LUT_AMPL_WIDTH),
		27784 => to_signed(15068, LUT_AMPL_WIDTH),
		27785 => to_signed(15065, LUT_AMPL_WIDTH),
		27786 => to_signed(15063, LUT_AMPL_WIDTH),
		27787 => to_signed(15060, LUT_AMPL_WIDTH),
		27788 => to_signed(15057, LUT_AMPL_WIDTH),
		27789 => to_signed(15054, LUT_AMPL_WIDTH),
		27790 => to_signed(15051, LUT_AMPL_WIDTH),
		27791 => to_signed(15049, LUT_AMPL_WIDTH),
		27792 => to_signed(15046, LUT_AMPL_WIDTH),
		27793 => to_signed(15043, LUT_AMPL_WIDTH),
		27794 => to_signed(15040, LUT_AMPL_WIDTH),
		27795 => to_signed(15037, LUT_AMPL_WIDTH),
		27796 => to_signed(15035, LUT_AMPL_WIDTH),
		27797 => to_signed(15032, LUT_AMPL_WIDTH),
		27798 => to_signed(15029, LUT_AMPL_WIDTH),
		27799 => to_signed(15026, LUT_AMPL_WIDTH),
		27800 => to_signed(15024, LUT_AMPL_WIDTH),
		27801 => to_signed(15021, LUT_AMPL_WIDTH),
		27802 => to_signed(15018, LUT_AMPL_WIDTH),
		27803 => to_signed(15015, LUT_AMPL_WIDTH),
		27804 => to_signed(15012, LUT_AMPL_WIDTH),
		27805 => to_signed(15010, LUT_AMPL_WIDTH),
		27806 => to_signed(15007, LUT_AMPL_WIDTH),
		27807 => to_signed(15004, LUT_AMPL_WIDTH),
		27808 => to_signed(15001, LUT_AMPL_WIDTH),
		27809 => to_signed(14998, LUT_AMPL_WIDTH),
		27810 => to_signed(14996, LUT_AMPL_WIDTH),
		27811 => to_signed(14993, LUT_AMPL_WIDTH),
		27812 => to_signed(14990, LUT_AMPL_WIDTH),
		27813 => to_signed(14987, LUT_AMPL_WIDTH),
		27814 => to_signed(14984, LUT_AMPL_WIDTH),
		27815 => to_signed(14982, LUT_AMPL_WIDTH),
		27816 => to_signed(14979, LUT_AMPL_WIDTH),
		27817 => to_signed(14976, LUT_AMPL_WIDTH),
		27818 => to_signed(14973, LUT_AMPL_WIDTH),
		27819 => to_signed(14970, LUT_AMPL_WIDTH),
		27820 => to_signed(14968, LUT_AMPL_WIDTH),
		27821 => to_signed(14965, LUT_AMPL_WIDTH),
		27822 => to_signed(14962, LUT_AMPL_WIDTH),
		27823 => to_signed(14959, LUT_AMPL_WIDTH),
		27824 => to_signed(14956, LUT_AMPL_WIDTH),
		27825 => to_signed(14954, LUT_AMPL_WIDTH),
		27826 => to_signed(14951, LUT_AMPL_WIDTH),
		27827 => to_signed(14948, LUT_AMPL_WIDTH),
		27828 => to_signed(14945, LUT_AMPL_WIDTH),
		27829 => to_signed(14942, LUT_AMPL_WIDTH),
		27830 => to_signed(14940, LUT_AMPL_WIDTH),
		27831 => to_signed(14937, LUT_AMPL_WIDTH),
		27832 => to_signed(14934, LUT_AMPL_WIDTH),
		27833 => to_signed(14931, LUT_AMPL_WIDTH),
		27834 => to_signed(14929, LUT_AMPL_WIDTH),
		27835 => to_signed(14926, LUT_AMPL_WIDTH),
		27836 => to_signed(14923, LUT_AMPL_WIDTH),
		27837 => to_signed(14920, LUT_AMPL_WIDTH),
		27838 => to_signed(14917, LUT_AMPL_WIDTH),
		27839 => to_signed(14915, LUT_AMPL_WIDTH),
		27840 => to_signed(14912, LUT_AMPL_WIDTH),
		27841 => to_signed(14909, LUT_AMPL_WIDTH),
		27842 => to_signed(14906, LUT_AMPL_WIDTH),
		27843 => to_signed(14903, LUT_AMPL_WIDTH),
		27844 => to_signed(14901, LUT_AMPL_WIDTH),
		27845 => to_signed(14898, LUT_AMPL_WIDTH),
		27846 => to_signed(14895, LUT_AMPL_WIDTH),
		27847 => to_signed(14892, LUT_AMPL_WIDTH),
		27848 => to_signed(14889, LUT_AMPL_WIDTH),
		27849 => to_signed(14887, LUT_AMPL_WIDTH),
		27850 => to_signed(14884, LUT_AMPL_WIDTH),
		27851 => to_signed(14881, LUT_AMPL_WIDTH),
		27852 => to_signed(14878, LUT_AMPL_WIDTH),
		27853 => to_signed(14875, LUT_AMPL_WIDTH),
		27854 => to_signed(14873, LUT_AMPL_WIDTH),
		27855 => to_signed(14870, LUT_AMPL_WIDTH),
		27856 => to_signed(14867, LUT_AMPL_WIDTH),
		27857 => to_signed(14864, LUT_AMPL_WIDTH),
		27858 => to_signed(14861, LUT_AMPL_WIDTH),
		27859 => to_signed(14859, LUT_AMPL_WIDTH),
		27860 => to_signed(14856, LUT_AMPL_WIDTH),
		27861 => to_signed(14853, LUT_AMPL_WIDTH),
		27862 => to_signed(14850, LUT_AMPL_WIDTH),
		27863 => to_signed(14847, LUT_AMPL_WIDTH),
		27864 => to_signed(14845, LUT_AMPL_WIDTH),
		27865 => to_signed(14842, LUT_AMPL_WIDTH),
		27866 => to_signed(14839, LUT_AMPL_WIDTH),
		27867 => to_signed(14836, LUT_AMPL_WIDTH),
		27868 => to_signed(14833, LUT_AMPL_WIDTH),
		27869 => to_signed(14831, LUT_AMPL_WIDTH),
		27870 => to_signed(14828, LUT_AMPL_WIDTH),
		27871 => to_signed(14825, LUT_AMPL_WIDTH),
		27872 => to_signed(14822, LUT_AMPL_WIDTH),
		27873 => to_signed(14819, LUT_AMPL_WIDTH),
		27874 => to_signed(14817, LUT_AMPL_WIDTH),
		27875 => to_signed(14814, LUT_AMPL_WIDTH),
		27876 => to_signed(14811, LUT_AMPL_WIDTH),
		27877 => to_signed(14808, LUT_AMPL_WIDTH),
		27878 => to_signed(14805, LUT_AMPL_WIDTH),
		27879 => to_signed(14803, LUT_AMPL_WIDTH),
		27880 => to_signed(14800, LUT_AMPL_WIDTH),
		27881 => to_signed(14797, LUT_AMPL_WIDTH),
		27882 => to_signed(14794, LUT_AMPL_WIDTH),
		27883 => to_signed(14791, LUT_AMPL_WIDTH),
		27884 => to_signed(14789, LUT_AMPL_WIDTH),
		27885 => to_signed(14786, LUT_AMPL_WIDTH),
		27886 => to_signed(14783, LUT_AMPL_WIDTH),
		27887 => to_signed(14780, LUT_AMPL_WIDTH),
		27888 => to_signed(14777, LUT_AMPL_WIDTH),
		27889 => to_signed(14774, LUT_AMPL_WIDTH),
		27890 => to_signed(14772, LUT_AMPL_WIDTH),
		27891 => to_signed(14769, LUT_AMPL_WIDTH),
		27892 => to_signed(14766, LUT_AMPL_WIDTH),
		27893 => to_signed(14763, LUT_AMPL_WIDTH),
		27894 => to_signed(14760, LUT_AMPL_WIDTH),
		27895 => to_signed(14758, LUT_AMPL_WIDTH),
		27896 => to_signed(14755, LUT_AMPL_WIDTH),
		27897 => to_signed(14752, LUT_AMPL_WIDTH),
		27898 => to_signed(14749, LUT_AMPL_WIDTH),
		27899 => to_signed(14746, LUT_AMPL_WIDTH),
		27900 => to_signed(14744, LUT_AMPL_WIDTH),
		27901 => to_signed(14741, LUT_AMPL_WIDTH),
		27902 => to_signed(14738, LUT_AMPL_WIDTH),
		27903 => to_signed(14735, LUT_AMPL_WIDTH),
		27904 => to_signed(14732, LUT_AMPL_WIDTH),
		27905 => to_signed(14730, LUT_AMPL_WIDTH),
		27906 => to_signed(14727, LUT_AMPL_WIDTH),
		27907 => to_signed(14724, LUT_AMPL_WIDTH),
		27908 => to_signed(14721, LUT_AMPL_WIDTH),
		27909 => to_signed(14718, LUT_AMPL_WIDTH),
		27910 => to_signed(14716, LUT_AMPL_WIDTH),
		27911 => to_signed(14713, LUT_AMPL_WIDTH),
		27912 => to_signed(14710, LUT_AMPL_WIDTH),
		27913 => to_signed(14707, LUT_AMPL_WIDTH),
		27914 => to_signed(14704, LUT_AMPL_WIDTH),
		27915 => to_signed(14702, LUT_AMPL_WIDTH),
		27916 => to_signed(14699, LUT_AMPL_WIDTH),
		27917 => to_signed(14696, LUT_AMPL_WIDTH),
		27918 => to_signed(14693, LUT_AMPL_WIDTH),
		27919 => to_signed(14690, LUT_AMPL_WIDTH),
		27920 => to_signed(14688, LUT_AMPL_WIDTH),
		27921 => to_signed(14685, LUT_AMPL_WIDTH),
		27922 => to_signed(14682, LUT_AMPL_WIDTH),
		27923 => to_signed(14679, LUT_AMPL_WIDTH),
		27924 => to_signed(14676, LUT_AMPL_WIDTH),
		27925 => to_signed(14673, LUT_AMPL_WIDTH),
		27926 => to_signed(14671, LUT_AMPL_WIDTH),
		27927 => to_signed(14668, LUT_AMPL_WIDTH),
		27928 => to_signed(14665, LUT_AMPL_WIDTH),
		27929 => to_signed(14662, LUT_AMPL_WIDTH),
		27930 => to_signed(14659, LUT_AMPL_WIDTH),
		27931 => to_signed(14657, LUT_AMPL_WIDTH),
		27932 => to_signed(14654, LUT_AMPL_WIDTH),
		27933 => to_signed(14651, LUT_AMPL_WIDTH),
		27934 => to_signed(14648, LUT_AMPL_WIDTH),
		27935 => to_signed(14645, LUT_AMPL_WIDTH),
		27936 => to_signed(14643, LUT_AMPL_WIDTH),
		27937 => to_signed(14640, LUT_AMPL_WIDTH),
		27938 => to_signed(14637, LUT_AMPL_WIDTH),
		27939 => to_signed(14634, LUT_AMPL_WIDTH),
		27940 => to_signed(14631, LUT_AMPL_WIDTH),
		27941 => to_signed(14628, LUT_AMPL_WIDTH),
		27942 => to_signed(14626, LUT_AMPL_WIDTH),
		27943 => to_signed(14623, LUT_AMPL_WIDTH),
		27944 => to_signed(14620, LUT_AMPL_WIDTH),
		27945 => to_signed(14617, LUT_AMPL_WIDTH),
		27946 => to_signed(14614, LUT_AMPL_WIDTH),
		27947 => to_signed(14612, LUT_AMPL_WIDTH),
		27948 => to_signed(14609, LUT_AMPL_WIDTH),
		27949 => to_signed(14606, LUT_AMPL_WIDTH),
		27950 => to_signed(14603, LUT_AMPL_WIDTH),
		27951 => to_signed(14600, LUT_AMPL_WIDTH),
		27952 => to_signed(14598, LUT_AMPL_WIDTH),
		27953 => to_signed(14595, LUT_AMPL_WIDTH),
		27954 => to_signed(14592, LUT_AMPL_WIDTH),
		27955 => to_signed(14589, LUT_AMPL_WIDTH),
		27956 => to_signed(14586, LUT_AMPL_WIDTH),
		27957 => to_signed(14584, LUT_AMPL_WIDTH),
		27958 => to_signed(14581, LUT_AMPL_WIDTH),
		27959 => to_signed(14578, LUT_AMPL_WIDTH),
		27960 => to_signed(14575, LUT_AMPL_WIDTH),
		27961 => to_signed(14572, LUT_AMPL_WIDTH),
		27962 => to_signed(14569, LUT_AMPL_WIDTH),
		27963 => to_signed(14567, LUT_AMPL_WIDTH),
		27964 => to_signed(14564, LUT_AMPL_WIDTH),
		27965 => to_signed(14561, LUT_AMPL_WIDTH),
		27966 => to_signed(14558, LUT_AMPL_WIDTH),
		27967 => to_signed(14555, LUT_AMPL_WIDTH),
		27968 => to_signed(14553, LUT_AMPL_WIDTH),
		27969 => to_signed(14550, LUT_AMPL_WIDTH),
		27970 => to_signed(14547, LUT_AMPL_WIDTH),
		27971 => to_signed(14544, LUT_AMPL_WIDTH),
		27972 => to_signed(14541, LUT_AMPL_WIDTH),
		27973 => to_signed(14538, LUT_AMPL_WIDTH),
		27974 => to_signed(14536, LUT_AMPL_WIDTH),
		27975 => to_signed(14533, LUT_AMPL_WIDTH),
		27976 => to_signed(14530, LUT_AMPL_WIDTH),
		27977 => to_signed(14527, LUT_AMPL_WIDTH),
		27978 => to_signed(14524, LUT_AMPL_WIDTH),
		27979 => to_signed(14522, LUT_AMPL_WIDTH),
		27980 => to_signed(14519, LUT_AMPL_WIDTH),
		27981 => to_signed(14516, LUT_AMPL_WIDTH),
		27982 => to_signed(14513, LUT_AMPL_WIDTH),
		27983 => to_signed(14510, LUT_AMPL_WIDTH),
		27984 => to_signed(14507, LUT_AMPL_WIDTH),
		27985 => to_signed(14505, LUT_AMPL_WIDTH),
		27986 => to_signed(14502, LUT_AMPL_WIDTH),
		27987 => to_signed(14499, LUT_AMPL_WIDTH),
		27988 => to_signed(14496, LUT_AMPL_WIDTH),
		27989 => to_signed(14493, LUT_AMPL_WIDTH),
		27990 => to_signed(14491, LUT_AMPL_WIDTH),
		27991 => to_signed(14488, LUT_AMPL_WIDTH),
		27992 => to_signed(14485, LUT_AMPL_WIDTH),
		27993 => to_signed(14482, LUT_AMPL_WIDTH),
		27994 => to_signed(14479, LUT_AMPL_WIDTH),
		27995 => to_signed(14477, LUT_AMPL_WIDTH),
		27996 => to_signed(14474, LUT_AMPL_WIDTH),
		27997 => to_signed(14471, LUT_AMPL_WIDTH),
		27998 => to_signed(14468, LUT_AMPL_WIDTH),
		27999 => to_signed(14465, LUT_AMPL_WIDTH),
		28000 => to_signed(14462, LUT_AMPL_WIDTH),
		28001 => to_signed(14460, LUT_AMPL_WIDTH),
		28002 => to_signed(14457, LUT_AMPL_WIDTH),
		28003 => to_signed(14454, LUT_AMPL_WIDTH),
		28004 => to_signed(14451, LUT_AMPL_WIDTH),
		28005 => to_signed(14448, LUT_AMPL_WIDTH),
		28006 => to_signed(14445, LUT_AMPL_WIDTH),
		28007 => to_signed(14443, LUT_AMPL_WIDTH),
		28008 => to_signed(14440, LUT_AMPL_WIDTH),
		28009 => to_signed(14437, LUT_AMPL_WIDTH),
		28010 => to_signed(14434, LUT_AMPL_WIDTH),
		28011 => to_signed(14431, LUT_AMPL_WIDTH),
		28012 => to_signed(14429, LUT_AMPL_WIDTH),
		28013 => to_signed(14426, LUT_AMPL_WIDTH),
		28014 => to_signed(14423, LUT_AMPL_WIDTH),
		28015 => to_signed(14420, LUT_AMPL_WIDTH),
		28016 => to_signed(14417, LUT_AMPL_WIDTH),
		28017 => to_signed(14414, LUT_AMPL_WIDTH),
		28018 => to_signed(14412, LUT_AMPL_WIDTH),
		28019 => to_signed(14409, LUT_AMPL_WIDTH),
		28020 => to_signed(14406, LUT_AMPL_WIDTH),
		28021 => to_signed(14403, LUT_AMPL_WIDTH),
		28022 => to_signed(14400, LUT_AMPL_WIDTH),
		28023 => to_signed(14398, LUT_AMPL_WIDTH),
		28024 => to_signed(14395, LUT_AMPL_WIDTH),
		28025 => to_signed(14392, LUT_AMPL_WIDTH),
		28026 => to_signed(14389, LUT_AMPL_WIDTH),
		28027 => to_signed(14386, LUT_AMPL_WIDTH),
		28028 => to_signed(14383, LUT_AMPL_WIDTH),
		28029 => to_signed(14381, LUT_AMPL_WIDTH),
		28030 => to_signed(14378, LUT_AMPL_WIDTH),
		28031 => to_signed(14375, LUT_AMPL_WIDTH),
		28032 => to_signed(14372, LUT_AMPL_WIDTH),
		28033 => to_signed(14369, LUT_AMPL_WIDTH),
		28034 => to_signed(14366, LUT_AMPL_WIDTH),
		28035 => to_signed(14364, LUT_AMPL_WIDTH),
		28036 => to_signed(14361, LUT_AMPL_WIDTH),
		28037 => to_signed(14358, LUT_AMPL_WIDTH),
		28038 => to_signed(14355, LUT_AMPL_WIDTH),
		28039 => to_signed(14352, LUT_AMPL_WIDTH),
		28040 => to_signed(14350, LUT_AMPL_WIDTH),
		28041 => to_signed(14347, LUT_AMPL_WIDTH),
		28042 => to_signed(14344, LUT_AMPL_WIDTH),
		28043 => to_signed(14341, LUT_AMPL_WIDTH),
		28044 => to_signed(14338, LUT_AMPL_WIDTH),
		28045 => to_signed(14335, LUT_AMPL_WIDTH),
		28046 => to_signed(14333, LUT_AMPL_WIDTH),
		28047 => to_signed(14330, LUT_AMPL_WIDTH),
		28048 => to_signed(14327, LUT_AMPL_WIDTH),
		28049 => to_signed(14324, LUT_AMPL_WIDTH),
		28050 => to_signed(14321, LUT_AMPL_WIDTH),
		28051 => to_signed(14318, LUT_AMPL_WIDTH),
		28052 => to_signed(14316, LUT_AMPL_WIDTH),
		28053 => to_signed(14313, LUT_AMPL_WIDTH),
		28054 => to_signed(14310, LUT_AMPL_WIDTH),
		28055 => to_signed(14307, LUT_AMPL_WIDTH),
		28056 => to_signed(14304, LUT_AMPL_WIDTH),
		28057 => to_signed(14302, LUT_AMPL_WIDTH),
		28058 => to_signed(14299, LUT_AMPL_WIDTH),
		28059 => to_signed(14296, LUT_AMPL_WIDTH),
		28060 => to_signed(14293, LUT_AMPL_WIDTH),
		28061 => to_signed(14290, LUT_AMPL_WIDTH),
		28062 => to_signed(14287, LUT_AMPL_WIDTH),
		28063 => to_signed(14285, LUT_AMPL_WIDTH),
		28064 => to_signed(14282, LUT_AMPL_WIDTH),
		28065 => to_signed(14279, LUT_AMPL_WIDTH),
		28066 => to_signed(14276, LUT_AMPL_WIDTH),
		28067 => to_signed(14273, LUT_AMPL_WIDTH),
		28068 => to_signed(14270, LUT_AMPL_WIDTH),
		28069 => to_signed(14268, LUT_AMPL_WIDTH),
		28070 => to_signed(14265, LUT_AMPL_WIDTH),
		28071 => to_signed(14262, LUT_AMPL_WIDTH),
		28072 => to_signed(14259, LUT_AMPL_WIDTH),
		28073 => to_signed(14256, LUT_AMPL_WIDTH),
		28074 => to_signed(14253, LUT_AMPL_WIDTH),
		28075 => to_signed(14251, LUT_AMPL_WIDTH),
		28076 => to_signed(14248, LUT_AMPL_WIDTH),
		28077 => to_signed(14245, LUT_AMPL_WIDTH),
		28078 => to_signed(14242, LUT_AMPL_WIDTH),
		28079 => to_signed(14239, LUT_AMPL_WIDTH),
		28080 => to_signed(14236, LUT_AMPL_WIDTH),
		28081 => to_signed(14234, LUT_AMPL_WIDTH),
		28082 => to_signed(14231, LUT_AMPL_WIDTH),
		28083 => to_signed(14228, LUT_AMPL_WIDTH),
		28084 => to_signed(14225, LUT_AMPL_WIDTH),
		28085 => to_signed(14222, LUT_AMPL_WIDTH),
		28086 => to_signed(14219, LUT_AMPL_WIDTH),
		28087 => to_signed(14217, LUT_AMPL_WIDTH),
		28088 => to_signed(14214, LUT_AMPL_WIDTH),
		28089 => to_signed(14211, LUT_AMPL_WIDTH),
		28090 => to_signed(14208, LUT_AMPL_WIDTH),
		28091 => to_signed(14205, LUT_AMPL_WIDTH),
		28092 => to_signed(14203, LUT_AMPL_WIDTH),
		28093 => to_signed(14200, LUT_AMPL_WIDTH),
		28094 => to_signed(14197, LUT_AMPL_WIDTH),
		28095 => to_signed(14194, LUT_AMPL_WIDTH),
		28096 => to_signed(14191, LUT_AMPL_WIDTH),
		28097 => to_signed(14188, LUT_AMPL_WIDTH),
		28098 => to_signed(14186, LUT_AMPL_WIDTH),
		28099 => to_signed(14183, LUT_AMPL_WIDTH),
		28100 => to_signed(14180, LUT_AMPL_WIDTH),
		28101 => to_signed(14177, LUT_AMPL_WIDTH),
		28102 => to_signed(14174, LUT_AMPL_WIDTH),
		28103 => to_signed(14171, LUT_AMPL_WIDTH),
		28104 => to_signed(14169, LUT_AMPL_WIDTH),
		28105 => to_signed(14166, LUT_AMPL_WIDTH),
		28106 => to_signed(14163, LUT_AMPL_WIDTH),
		28107 => to_signed(14160, LUT_AMPL_WIDTH),
		28108 => to_signed(14157, LUT_AMPL_WIDTH),
		28109 => to_signed(14154, LUT_AMPL_WIDTH),
		28110 => to_signed(14152, LUT_AMPL_WIDTH),
		28111 => to_signed(14149, LUT_AMPL_WIDTH),
		28112 => to_signed(14146, LUT_AMPL_WIDTH),
		28113 => to_signed(14143, LUT_AMPL_WIDTH),
		28114 => to_signed(14140, LUT_AMPL_WIDTH),
		28115 => to_signed(14137, LUT_AMPL_WIDTH),
		28116 => to_signed(14135, LUT_AMPL_WIDTH),
		28117 => to_signed(14132, LUT_AMPL_WIDTH),
		28118 => to_signed(14129, LUT_AMPL_WIDTH),
		28119 => to_signed(14126, LUT_AMPL_WIDTH),
		28120 => to_signed(14123, LUT_AMPL_WIDTH),
		28121 => to_signed(14120, LUT_AMPL_WIDTH),
		28122 => to_signed(14118, LUT_AMPL_WIDTH),
		28123 => to_signed(14115, LUT_AMPL_WIDTH),
		28124 => to_signed(14112, LUT_AMPL_WIDTH),
		28125 => to_signed(14109, LUT_AMPL_WIDTH),
		28126 => to_signed(14106, LUT_AMPL_WIDTH),
		28127 => to_signed(14103, LUT_AMPL_WIDTH),
		28128 => to_signed(14101, LUT_AMPL_WIDTH),
		28129 => to_signed(14098, LUT_AMPL_WIDTH),
		28130 => to_signed(14095, LUT_AMPL_WIDTH),
		28131 => to_signed(14092, LUT_AMPL_WIDTH),
		28132 => to_signed(14089, LUT_AMPL_WIDTH),
		28133 => to_signed(14086, LUT_AMPL_WIDTH),
		28134 => to_signed(14083, LUT_AMPL_WIDTH),
		28135 => to_signed(14081, LUT_AMPL_WIDTH),
		28136 => to_signed(14078, LUT_AMPL_WIDTH),
		28137 => to_signed(14075, LUT_AMPL_WIDTH),
		28138 => to_signed(14072, LUT_AMPL_WIDTH),
		28139 => to_signed(14069, LUT_AMPL_WIDTH),
		28140 => to_signed(14066, LUT_AMPL_WIDTH),
		28141 => to_signed(14064, LUT_AMPL_WIDTH),
		28142 => to_signed(14061, LUT_AMPL_WIDTH),
		28143 => to_signed(14058, LUT_AMPL_WIDTH),
		28144 => to_signed(14055, LUT_AMPL_WIDTH),
		28145 => to_signed(14052, LUT_AMPL_WIDTH),
		28146 => to_signed(14049, LUT_AMPL_WIDTH),
		28147 => to_signed(14047, LUT_AMPL_WIDTH),
		28148 => to_signed(14044, LUT_AMPL_WIDTH),
		28149 => to_signed(14041, LUT_AMPL_WIDTH),
		28150 => to_signed(14038, LUT_AMPL_WIDTH),
		28151 => to_signed(14035, LUT_AMPL_WIDTH),
		28152 => to_signed(14032, LUT_AMPL_WIDTH),
		28153 => to_signed(14030, LUT_AMPL_WIDTH),
		28154 => to_signed(14027, LUT_AMPL_WIDTH),
		28155 => to_signed(14024, LUT_AMPL_WIDTH),
		28156 => to_signed(14021, LUT_AMPL_WIDTH),
		28157 => to_signed(14018, LUT_AMPL_WIDTH),
		28158 => to_signed(14015, LUT_AMPL_WIDTH),
		28159 => to_signed(14013, LUT_AMPL_WIDTH),
		28160 => to_signed(14010, LUT_AMPL_WIDTH),
		28161 => to_signed(14007, LUT_AMPL_WIDTH),
		28162 => to_signed(14004, LUT_AMPL_WIDTH),
		28163 => to_signed(14001, LUT_AMPL_WIDTH),
		28164 => to_signed(13998, LUT_AMPL_WIDTH),
		28165 => to_signed(13995, LUT_AMPL_WIDTH),
		28166 => to_signed(13993, LUT_AMPL_WIDTH),
		28167 => to_signed(13990, LUT_AMPL_WIDTH),
		28168 => to_signed(13987, LUT_AMPL_WIDTH),
		28169 => to_signed(13984, LUT_AMPL_WIDTH),
		28170 => to_signed(13981, LUT_AMPL_WIDTH),
		28171 => to_signed(13978, LUT_AMPL_WIDTH),
		28172 => to_signed(13976, LUT_AMPL_WIDTH),
		28173 => to_signed(13973, LUT_AMPL_WIDTH),
		28174 => to_signed(13970, LUT_AMPL_WIDTH),
		28175 => to_signed(13967, LUT_AMPL_WIDTH),
		28176 => to_signed(13964, LUT_AMPL_WIDTH),
		28177 => to_signed(13961, LUT_AMPL_WIDTH),
		28178 => to_signed(13959, LUT_AMPL_WIDTH),
		28179 => to_signed(13956, LUT_AMPL_WIDTH),
		28180 => to_signed(13953, LUT_AMPL_WIDTH),
		28181 => to_signed(13950, LUT_AMPL_WIDTH),
		28182 => to_signed(13947, LUT_AMPL_WIDTH),
		28183 => to_signed(13944, LUT_AMPL_WIDTH),
		28184 => to_signed(13942, LUT_AMPL_WIDTH),
		28185 => to_signed(13939, LUT_AMPL_WIDTH),
		28186 => to_signed(13936, LUT_AMPL_WIDTH),
		28187 => to_signed(13933, LUT_AMPL_WIDTH),
		28188 => to_signed(13930, LUT_AMPL_WIDTH),
		28189 => to_signed(13927, LUT_AMPL_WIDTH),
		28190 => to_signed(13924, LUT_AMPL_WIDTH),
		28191 => to_signed(13922, LUT_AMPL_WIDTH),
		28192 => to_signed(13919, LUT_AMPL_WIDTH),
		28193 => to_signed(13916, LUT_AMPL_WIDTH),
		28194 => to_signed(13913, LUT_AMPL_WIDTH),
		28195 => to_signed(13910, LUT_AMPL_WIDTH),
		28196 => to_signed(13907, LUT_AMPL_WIDTH),
		28197 => to_signed(13905, LUT_AMPL_WIDTH),
		28198 => to_signed(13902, LUT_AMPL_WIDTH),
		28199 => to_signed(13899, LUT_AMPL_WIDTH),
		28200 => to_signed(13896, LUT_AMPL_WIDTH),
		28201 => to_signed(13893, LUT_AMPL_WIDTH),
		28202 => to_signed(13890, LUT_AMPL_WIDTH),
		28203 => to_signed(13887, LUT_AMPL_WIDTH),
		28204 => to_signed(13885, LUT_AMPL_WIDTH),
		28205 => to_signed(13882, LUT_AMPL_WIDTH),
		28206 => to_signed(13879, LUT_AMPL_WIDTH),
		28207 => to_signed(13876, LUT_AMPL_WIDTH),
		28208 => to_signed(13873, LUT_AMPL_WIDTH),
		28209 => to_signed(13870, LUT_AMPL_WIDTH),
		28210 => to_signed(13868, LUT_AMPL_WIDTH),
		28211 => to_signed(13865, LUT_AMPL_WIDTH),
		28212 => to_signed(13862, LUT_AMPL_WIDTH),
		28213 => to_signed(13859, LUT_AMPL_WIDTH),
		28214 => to_signed(13856, LUT_AMPL_WIDTH),
		28215 => to_signed(13853, LUT_AMPL_WIDTH),
		28216 => to_signed(13850, LUT_AMPL_WIDTH),
		28217 => to_signed(13848, LUT_AMPL_WIDTH),
		28218 => to_signed(13845, LUT_AMPL_WIDTH),
		28219 => to_signed(13842, LUT_AMPL_WIDTH),
		28220 => to_signed(13839, LUT_AMPL_WIDTH),
		28221 => to_signed(13836, LUT_AMPL_WIDTH),
		28222 => to_signed(13833, LUT_AMPL_WIDTH),
		28223 => to_signed(13831, LUT_AMPL_WIDTH),
		28224 => to_signed(13828, LUT_AMPL_WIDTH),
		28225 => to_signed(13825, LUT_AMPL_WIDTH),
		28226 => to_signed(13822, LUT_AMPL_WIDTH),
		28227 => to_signed(13819, LUT_AMPL_WIDTH),
		28228 => to_signed(13816, LUT_AMPL_WIDTH),
		28229 => to_signed(13813, LUT_AMPL_WIDTH),
		28230 => to_signed(13811, LUT_AMPL_WIDTH),
		28231 => to_signed(13808, LUT_AMPL_WIDTH),
		28232 => to_signed(13805, LUT_AMPL_WIDTH),
		28233 => to_signed(13802, LUT_AMPL_WIDTH),
		28234 => to_signed(13799, LUT_AMPL_WIDTH),
		28235 => to_signed(13796, LUT_AMPL_WIDTH),
		28236 => to_signed(13793, LUT_AMPL_WIDTH),
		28237 => to_signed(13791, LUT_AMPL_WIDTH),
		28238 => to_signed(13788, LUT_AMPL_WIDTH),
		28239 => to_signed(13785, LUT_AMPL_WIDTH),
		28240 => to_signed(13782, LUT_AMPL_WIDTH),
		28241 => to_signed(13779, LUT_AMPL_WIDTH),
		28242 => to_signed(13776, LUT_AMPL_WIDTH),
		28243 => to_signed(13774, LUT_AMPL_WIDTH),
		28244 => to_signed(13771, LUT_AMPL_WIDTH),
		28245 => to_signed(13768, LUT_AMPL_WIDTH),
		28246 => to_signed(13765, LUT_AMPL_WIDTH),
		28247 => to_signed(13762, LUT_AMPL_WIDTH),
		28248 => to_signed(13759, LUT_AMPL_WIDTH),
		28249 => to_signed(13756, LUT_AMPL_WIDTH),
		28250 => to_signed(13754, LUT_AMPL_WIDTH),
		28251 => to_signed(13751, LUT_AMPL_WIDTH),
		28252 => to_signed(13748, LUT_AMPL_WIDTH),
		28253 => to_signed(13745, LUT_AMPL_WIDTH),
		28254 => to_signed(13742, LUT_AMPL_WIDTH),
		28255 => to_signed(13739, LUT_AMPL_WIDTH),
		28256 => to_signed(13736, LUT_AMPL_WIDTH),
		28257 => to_signed(13734, LUT_AMPL_WIDTH),
		28258 => to_signed(13731, LUT_AMPL_WIDTH),
		28259 => to_signed(13728, LUT_AMPL_WIDTH),
		28260 => to_signed(13725, LUT_AMPL_WIDTH),
		28261 => to_signed(13722, LUT_AMPL_WIDTH),
		28262 => to_signed(13719, LUT_AMPL_WIDTH),
		28263 => to_signed(13717, LUT_AMPL_WIDTH),
		28264 => to_signed(13714, LUT_AMPL_WIDTH),
		28265 => to_signed(13711, LUT_AMPL_WIDTH),
		28266 => to_signed(13708, LUT_AMPL_WIDTH),
		28267 => to_signed(13705, LUT_AMPL_WIDTH),
		28268 => to_signed(13702, LUT_AMPL_WIDTH),
		28269 => to_signed(13699, LUT_AMPL_WIDTH),
		28270 => to_signed(13697, LUT_AMPL_WIDTH),
		28271 => to_signed(13694, LUT_AMPL_WIDTH),
		28272 => to_signed(13691, LUT_AMPL_WIDTH),
		28273 => to_signed(13688, LUT_AMPL_WIDTH),
		28274 => to_signed(13685, LUT_AMPL_WIDTH),
		28275 => to_signed(13682, LUT_AMPL_WIDTH),
		28276 => to_signed(13679, LUT_AMPL_WIDTH),
		28277 => to_signed(13677, LUT_AMPL_WIDTH),
		28278 => to_signed(13674, LUT_AMPL_WIDTH),
		28279 => to_signed(13671, LUT_AMPL_WIDTH),
		28280 => to_signed(13668, LUT_AMPL_WIDTH),
		28281 => to_signed(13665, LUT_AMPL_WIDTH),
		28282 => to_signed(13662, LUT_AMPL_WIDTH),
		28283 => to_signed(13659, LUT_AMPL_WIDTH),
		28284 => to_signed(13657, LUT_AMPL_WIDTH),
		28285 => to_signed(13654, LUT_AMPL_WIDTH),
		28286 => to_signed(13651, LUT_AMPL_WIDTH),
		28287 => to_signed(13648, LUT_AMPL_WIDTH),
		28288 => to_signed(13645, LUT_AMPL_WIDTH),
		28289 => to_signed(13642, LUT_AMPL_WIDTH),
		28290 => to_signed(13639, LUT_AMPL_WIDTH),
		28291 => to_signed(13637, LUT_AMPL_WIDTH),
		28292 => to_signed(13634, LUT_AMPL_WIDTH),
		28293 => to_signed(13631, LUT_AMPL_WIDTH),
		28294 => to_signed(13628, LUT_AMPL_WIDTH),
		28295 => to_signed(13625, LUT_AMPL_WIDTH),
		28296 => to_signed(13622, LUT_AMPL_WIDTH),
		28297 => to_signed(13619, LUT_AMPL_WIDTH),
		28298 => to_signed(13617, LUT_AMPL_WIDTH),
		28299 => to_signed(13614, LUT_AMPL_WIDTH),
		28300 => to_signed(13611, LUT_AMPL_WIDTH),
		28301 => to_signed(13608, LUT_AMPL_WIDTH),
		28302 => to_signed(13605, LUT_AMPL_WIDTH),
		28303 => to_signed(13602, LUT_AMPL_WIDTH),
		28304 => to_signed(13599, LUT_AMPL_WIDTH),
		28305 => to_signed(13597, LUT_AMPL_WIDTH),
		28306 => to_signed(13594, LUT_AMPL_WIDTH),
		28307 => to_signed(13591, LUT_AMPL_WIDTH),
		28308 => to_signed(13588, LUT_AMPL_WIDTH),
		28309 => to_signed(13585, LUT_AMPL_WIDTH),
		28310 => to_signed(13582, LUT_AMPL_WIDTH),
		28311 => to_signed(13579, LUT_AMPL_WIDTH),
		28312 => to_signed(13577, LUT_AMPL_WIDTH),
		28313 => to_signed(13574, LUT_AMPL_WIDTH),
		28314 => to_signed(13571, LUT_AMPL_WIDTH),
		28315 => to_signed(13568, LUT_AMPL_WIDTH),
		28316 => to_signed(13565, LUT_AMPL_WIDTH),
		28317 => to_signed(13562, LUT_AMPL_WIDTH),
		28318 => to_signed(13559, LUT_AMPL_WIDTH),
		28319 => to_signed(13557, LUT_AMPL_WIDTH),
		28320 => to_signed(13554, LUT_AMPL_WIDTH),
		28321 => to_signed(13551, LUT_AMPL_WIDTH),
		28322 => to_signed(13548, LUT_AMPL_WIDTH),
		28323 => to_signed(13545, LUT_AMPL_WIDTH),
		28324 => to_signed(13542, LUT_AMPL_WIDTH),
		28325 => to_signed(13539, LUT_AMPL_WIDTH),
		28326 => to_signed(13537, LUT_AMPL_WIDTH),
		28327 => to_signed(13534, LUT_AMPL_WIDTH),
		28328 => to_signed(13531, LUT_AMPL_WIDTH),
		28329 => to_signed(13528, LUT_AMPL_WIDTH),
		28330 => to_signed(13525, LUT_AMPL_WIDTH),
		28331 => to_signed(13522, LUT_AMPL_WIDTH),
		28332 => to_signed(13519, LUT_AMPL_WIDTH),
		28333 => to_signed(13516, LUT_AMPL_WIDTH),
		28334 => to_signed(13514, LUT_AMPL_WIDTH),
		28335 => to_signed(13511, LUT_AMPL_WIDTH),
		28336 => to_signed(13508, LUT_AMPL_WIDTH),
		28337 => to_signed(13505, LUT_AMPL_WIDTH),
		28338 => to_signed(13502, LUT_AMPL_WIDTH),
		28339 => to_signed(13499, LUT_AMPL_WIDTH),
		28340 => to_signed(13496, LUT_AMPL_WIDTH),
		28341 => to_signed(13494, LUT_AMPL_WIDTH),
		28342 => to_signed(13491, LUT_AMPL_WIDTH),
		28343 => to_signed(13488, LUT_AMPL_WIDTH),
		28344 => to_signed(13485, LUT_AMPL_WIDTH),
		28345 => to_signed(13482, LUT_AMPL_WIDTH),
		28346 => to_signed(13479, LUT_AMPL_WIDTH),
		28347 => to_signed(13476, LUT_AMPL_WIDTH),
		28348 => to_signed(13474, LUT_AMPL_WIDTH),
		28349 => to_signed(13471, LUT_AMPL_WIDTH),
		28350 => to_signed(13468, LUT_AMPL_WIDTH),
		28351 => to_signed(13465, LUT_AMPL_WIDTH),
		28352 => to_signed(13462, LUT_AMPL_WIDTH),
		28353 => to_signed(13459, LUT_AMPL_WIDTH),
		28354 => to_signed(13456, LUT_AMPL_WIDTH),
		28355 => to_signed(13454, LUT_AMPL_WIDTH),
		28356 => to_signed(13451, LUT_AMPL_WIDTH),
		28357 => to_signed(13448, LUT_AMPL_WIDTH),
		28358 => to_signed(13445, LUT_AMPL_WIDTH),
		28359 => to_signed(13442, LUT_AMPL_WIDTH),
		28360 => to_signed(13439, LUT_AMPL_WIDTH),
		28361 => to_signed(13436, LUT_AMPL_WIDTH),
		28362 => to_signed(13433, LUT_AMPL_WIDTH),
		28363 => to_signed(13431, LUT_AMPL_WIDTH),
		28364 => to_signed(13428, LUT_AMPL_WIDTH),
		28365 => to_signed(13425, LUT_AMPL_WIDTH),
		28366 => to_signed(13422, LUT_AMPL_WIDTH),
		28367 => to_signed(13419, LUT_AMPL_WIDTH),
		28368 => to_signed(13416, LUT_AMPL_WIDTH),
		28369 => to_signed(13413, LUT_AMPL_WIDTH),
		28370 => to_signed(13411, LUT_AMPL_WIDTH),
		28371 => to_signed(13408, LUT_AMPL_WIDTH),
		28372 => to_signed(13405, LUT_AMPL_WIDTH),
		28373 => to_signed(13402, LUT_AMPL_WIDTH),
		28374 => to_signed(13399, LUT_AMPL_WIDTH),
		28375 => to_signed(13396, LUT_AMPL_WIDTH),
		28376 => to_signed(13393, LUT_AMPL_WIDTH),
		28377 => to_signed(13390, LUT_AMPL_WIDTH),
		28378 => to_signed(13388, LUT_AMPL_WIDTH),
		28379 => to_signed(13385, LUT_AMPL_WIDTH),
		28380 => to_signed(13382, LUT_AMPL_WIDTH),
		28381 => to_signed(13379, LUT_AMPL_WIDTH),
		28382 => to_signed(13376, LUT_AMPL_WIDTH),
		28383 => to_signed(13373, LUT_AMPL_WIDTH),
		28384 => to_signed(13370, LUT_AMPL_WIDTH),
		28385 => to_signed(13368, LUT_AMPL_WIDTH),
		28386 => to_signed(13365, LUT_AMPL_WIDTH),
		28387 => to_signed(13362, LUT_AMPL_WIDTH),
		28388 => to_signed(13359, LUT_AMPL_WIDTH),
		28389 => to_signed(13356, LUT_AMPL_WIDTH),
		28390 => to_signed(13353, LUT_AMPL_WIDTH),
		28391 => to_signed(13350, LUT_AMPL_WIDTH),
		28392 => to_signed(13347, LUT_AMPL_WIDTH),
		28393 => to_signed(13345, LUT_AMPL_WIDTH),
		28394 => to_signed(13342, LUT_AMPL_WIDTH),
		28395 => to_signed(13339, LUT_AMPL_WIDTH),
		28396 => to_signed(13336, LUT_AMPL_WIDTH),
		28397 => to_signed(13333, LUT_AMPL_WIDTH),
		28398 => to_signed(13330, LUT_AMPL_WIDTH),
		28399 => to_signed(13327, LUT_AMPL_WIDTH),
		28400 => to_signed(13324, LUT_AMPL_WIDTH),
		28401 => to_signed(13322, LUT_AMPL_WIDTH),
		28402 => to_signed(13319, LUT_AMPL_WIDTH),
		28403 => to_signed(13316, LUT_AMPL_WIDTH),
		28404 => to_signed(13313, LUT_AMPL_WIDTH),
		28405 => to_signed(13310, LUT_AMPL_WIDTH),
		28406 => to_signed(13307, LUT_AMPL_WIDTH),
		28407 => to_signed(13304, LUT_AMPL_WIDTH),
		28408 => to_signed(13302, LUT_AMPL_WIDTH),
		28409 => to_signed(13299, LUT_AMPL_WIDTH),
		28410 => to_signed(13296, LUT_AMPL_WIDTH),
		28411 => to_signed(13293, LUT_AMPL_WIDTH),
		28412 => to_signed(13290, LUT_AMPL_WIDTH),
		28413 => to_signed(13287, LUT_AMPL_WIDTH),
		28414 => to_signed(13284, LUT_AMPL_WIDTH),
		28415 => to_signed(13281, LUT_AMPL_WIDTH),
		28416 => to_signed(13279, LUT_AMPL_WIDTH),
		28417 => to_signed(13276, LUT_AMPL_WIDTH),
		28418 => to_signed(13273, LUT_AMPL_WIDTH),
		28419 => to_signed(13270, LUT_AMPL_WIDTH),
		28420 => to_signed(13267, LUT_AMPL_WIDTH),
		28421 => to_signed(13264, LUT_AMPL_WIDTH),
		28422 => to_signed(13261, LUT_AMPL_WIDTH),
		28423 => to_signed(13258, LUT_AMPL_WIDTH),
		28424 => to_signed(13256, LUT_AMPL_WIDTH),
		28425 => to_signed(13253, LUT_AMPL_WIDTH),
		28426 => to_signed(13250, LUT_AMPL_WIDTH),
		28427 => to_signed(13247, LUT_AMPL_WIDTH),
		28428 => to_signed(13244, LUT_AMPL_WIDTH),
		28429 => to_signed(13241, LUT_AMPL_WIDTH),
		28430 => to_signed(13238, LUT_AMPL_WIDTH),
		28431 => to_signed(13235, LUT_AMPL_WIDTH),
		28432 => to_signed(13233, LUT_AMPL_WIDTH),
		28433 => to_signed(13230, LUT_AMPL_WIDTH),
		28434 => to_signed(13227, LUT_AMPL_WIDTH),
		28435 => to_signed(13224, LUT_AMPL_WIDTH),
		28436 => to_signed(13221, LUT_AMPL_WIDTH),
		28437 => to_signed(13218, LUT_AMPL_WIDTH),
		28438 => to_signed(13215, LUT_AMPL_WIDTH),
		28439 => to_signed(13212, LUT_AMPL_WIDTH),
		28440 => to_signed(13210, LUT_AMPL_WIDTH),
		28441 => to_signed(13207, LUT_AMPL_WIDTH),
		28442 => to_signed(13204, LUT_AMPL_WIDTH),
		28443 => to_signed(13201, LUT_AMPL_WIDTH),
		28444 => to_signed(13198, LUT_AMPL_WIDTH),
		28445 => to_signed(13195, LUT_AMPL_WIDTH),
		28446 => to_signed(13192, LUT_AMPL_WIDTH),
		28447 => to_signed(13189, LUT_AMPL_WIDTH),
		28448 => to_signed(13187, LUT_AMPL_WIDTH),
		28449 => to_signed(13184, LUT_AMPL_WIDTH),
		28450 => to_signed(13181, LUT_AMPL_WIDTH),
		28451 => to_signed(13178, LUT_AMPL_WIDTH),
		28452 => to_signed(13175, LUT_AMPL_WIDTH),
		28453 => to_signed(13172, LUT_AMPL_WIDTH),
		28454 => to_signed(13169, LUT_AMPL_WIDTH),
		28455 => to_signed(13166, LUT_AMPL_WIDTH),
		28456 => to_signed(13164, LUT_AMPL_WIDTH),
		28457 => to_signed(13161, LUT_AMPL_WIDTH),
		28458 => to_signed(13158, LUT_AMPL_WIDTH),
		28459 => to_signed(13155, LUT_AMPL_WIDTH),
		28460 => to_signed(13152, LUT_AMPL_WIDTH),
		28461 => to_signed(13149, LUT_AMPL_WIDTH),
		28462 => to_signed(13146, LUT_AMPL_WIDTH),
		28463 => to_signed(13143, LUT_AMPL_WIDTH),
		28464 => to_signed(13141, LUT_AMPL_WIDTH),
		28465 => to_signed(13138, LUT_AMPL_WIDTH),
		28466 => to_signed(13135, LUT_AMPL_WIDTH),
		28467 => to_signed(13132, LUT_AMPL_WIDTH),
		28468 => to_signed(13129, LUT_AMPL_WIDTH),
		28469 => to_signed(13126, LUT_AMPL_WIDTH),
		28470 => to_signed(13123, LUT_AMPL_WIDTH),
		28471 => to_signed(13120, LUT_AMPL_WIDTH),
		28472 => to_signed(13118, LUT_AMPL_WIDTH),
		28473 => to_signed(13115, LUT_AMPL_WIDTH),
		28474 => to_signed(13112, LUT_AMPL_WIDTH),
		28475 => to_signed(13109, LUT_AMPL_WIDTH),
		28476 => to_signed(13106, LUT_AMPL_WIDTH),
		28477 => to_signed(13103, LUT_AMPL_WIDTH),
		28478 => to_signed(13100, LUT_AMPL_WIDTH),
		28479 => to_signed(13097, LUT_AMPL_WIDTH),
		28480 => to_signed(13094, LUT_AMPL_WIDTH),
		28481 => to_signed(13092, LUT_AMPL_WIDTH),
		28482 => to_signed(13089, LUT_AMPL_WIDTH),
		28483 => to_signed(13086, LUT_AMPL_WIDTH),
		28484 => to_signed(13083, LUT_AMPL_WIDTH),
		28485 => to_signed(13080, LUT_AMPL_WIDTH),
		28486 => to_signed(13077, LUT_AMPL_WIDTH),
		28487 => to_signed(13074, LUT_AMPL_WIDTH),
		28488 => to_signed(13071, LUT_AMPL_WIDTH),
		28489 => to_signed(13069, LUT_AMPL_WIDTH),
		28490 => to_signed(13066, LUT_AMPL_WIDTH),
		28491 => to_signed(13063, LUT_AMPL_WIDTH),
		28492 => to_signed(13060, LUT_AMPL_WIDTH),
		28493 => to_signed(13057, LUT_AMPL_WIDTH),
		28494 => to_signed(13054, LUT_AMPL_WIDTH),
		28495 => to_signed(13051, LUT_AMPL_WIDTH),
		28496 => to_signed(13048, LUT_AMPL_WIDTH),
		28497 => to_signed(13046, LUT_AMPL_WIDTH),
		28498 => to_signed(13043, LUT_AMPL_WIDTH),
		28499 => to_signed(13040, LUT_AMPL_WIDTH),
		28500 => to_signed(13037, LUT_AMPL_WIDTH),
		28501 => to_signed(13034, LUT_AMPL_WIDTH),
		28502 => to_signed(13031, LUT_AMPL_WIDTH),
		28503 => to_signed(13028, LUT_AMPL_WIDTH),
		28504 => to_signed(13025, LUT_AMPL_WIDTH),
		28505 => to_signed(13022, LUT_AMPL_WIDTH),
		28506 => to_signed(13020, LUT_AMPL_WIDTH),
		28507 => to_signed(13017, LUT_AMPL_WIDTH),
		28508 => to_signed(13014, LUT_AMPL_WIDTH),
		28509 => to_signed(13011, LUT_AMPL_WIDTH),
		28510 => to_signed(13008, LUT_AMPL_WIDTH),
		28511 => to_signed(13005, LUT_AMPL_WIDTH),
		28512 => to_signed(13002, LUT_AMPL_WIDTH),
		28513 => to_signed(12999, LUT_AMPL_WIDTH),
		28514 => to_signed(12997, LUT_AMPL_WIDTH),
		28515 => to_signed(12994, LUT_AMPL_WIDTH),
		28516 => to_signed(12991, LUT_AMPL_WIDTH),
		28517 => to_signed(12988, LUT_AMPL_WIDTH),
		28518 => to_signed(12985, LUT_AMPL_WIDTH),
		28519 => to_signed(12982, LUT_AMPL_WIDTH),
		28520 => to_signed(12979, LUT_AMPL_WIDTH),
		28521 => to_signed(12976, LUT_AMPL_WIDTH),
		28522 => to_signed(12973, LUT_AMPL_WIDTH),
		28523 => to_signed(12971, LUT_AMPL_WIDTH),
		28524 => to_signed(12968, LUT_AMPL_WIDTH),
		28525 => to_signed(12965, LUT_AMPL_WIDTH),
		28526 => to_signed(12962, LUT_AMPL_WIDTH),
		28527 => to_signed(12959, LUT_AMPL_WIDTH),
		28528 => to_signed(12956, LUT_AMPL_WIDTH),
		28529 => to_signed(12953, LUT_AMPL_WIDTH),
		28530 => to_signed(12950, LUT_AMPL_WIDTH),
		28531 => to_signed(12947, LUT_AMPL_WIDTH),
		28532 => to_signed(12945, LUT_AMPL_WIDTH),
		28533 => to_signed(12942, LUT_AMPL_WIDTH),
		28534 => to_signed(12939, LUT_AMPL_WIDTH),
		28535 => to_signed(12936, LUT_AMPL_WIDTH),
		28536 => to_signed(12933, LUT_AMPL_WIDTH),
		28537 => to_signed(12930, LUT_AMPL_WIDTH),
		28538 => to_signed(12927, LUT_AMPL_WIDTH),
		28539 => to_signed(12924, LUT_AMPL_WIDTH),
		28540 => to_signed(12921, LUT_AMPL_WIDTH),
		28541 => to_signed(12919, LUT_AMPL_WIDTH),
		28542 => to_signed(12916, LUT_AMPL_WIDTH),
		28543 => to_signed(12913, LUT_AMPL_WIDTH),
		28544 => to_signed(12910, LUT_AMPL_WIDTH),
		28545 => to_signed(12907, LUT_AMPL_WIDTH),
		28546 => to_signed(12904, LUT_AMPL_WIDTH),
		28547 => to_signed(12901, LUT_AMPL_WIDTH),
		28548 => to_signed(12898, LUT_AMPL_WIDTH),
		28549 => to_signed(12895, LUT_AMPL_WIDTH),
		28550 => to_signed(12893, LUT_AMPL_WIDTH),
		28551 => to_signed(12890, LUT_AMPL_WIDTH),
		28552 => to_signed(12887, LUT_AMPL_WIDTH),
		28553 => to_signed(12884, LUT_AMPL_WIDTH),
		28554 => to_signed(12881, LUT_AMPL_WIDTH),
		28555 => to_signed(12878, LUT_AMPL_WIDTH),
		28556 => to_signed(12875, LUT_AMPL_WIDTH),
		28557 => to_signed(12872, LUT_AMPL_WIDTH),
		28558 => to_signed(12870, LUT_AMPL_WIDTH),
		28559 => to_signed(12867, LUT_AMPL_WIDTH),
		28560 => to_signed(12864, LUT_AMPL_WIDTH),
		28561 => to_signed(12861, LUT_AMPL_WIDTH),
		28562 => to_signed(12858, LUT_AMPL_WIDTH),
		28563 => to_signed(12855, LUT_AMPL_WIDTH),
		28564 => to_signed(12852, LUT_AMPL_WIDTH),
		28565 => to_signed(12849, LUT_AMPL_WIDTH),
		28566 => to_signed(12846, LUT_AMPL_WIDTH),
		28567 => to_signed(12843, LUT_AMPL_WIDTH),
		28568 => to_signed(12841, LUT_AMPL_WIDTH),
		28569 => to_signed(12838, LUT_AMPL_WIDTH),
		28570 => to_signed(12835, LUT_AMPL_WIDTH),
		28571 => to_signed(12832, LUT_AMPL_WIDTH),
		28572 => to_signed(12829, LUT_AMPL_WIDTH),
		28573 => to_signed(12826, LUT_AMPL_WIDTH),
		28574 => to_signed(12823, LUT_AMPL_WIDTH),
		28575 => to_signed(12820, LUT_AMPL_WIDTH),
		28576 => to_signed(12817, LUT_AMPL_WIDTH),
		28577 => to_signed(12815, LUT_AMPL_WIDTH),
		28578 => to_signed(12812, LUT_AMPL_WIDTH),
		28579 => to_signed(12809, LUT_AMPL_WIDTH),
		28580 => to_signed(12806, LUT_AMPL_WIDTH),
		28581 => to_signed(12803, LUT_AMPL_WIDTH),
		28582 => to_signed(12800, LUT_AMPL_WIDTH),
		28583 => to_signed(12797, LUT_AMPL_WIDTH),
		28584 => to_signed(12794, LUT_AMPL_WIDTH),
		28585 => to_signed(12791, LUT_AMPL_WIDTH),
		28586 => to_signed(12789, LUT_AMPL_WIDTH),
		28587 => to_signed(12786, LUT_AMPL_WIDTH),
		28588 => to_signed(12783, LUT_AMPL_WIDTH),
		28589 => to_signed(12780, LUT_AMPL_WIDTH),
		28590 => to_signed(12777, LUT_AMPL_WIDTH),
		28591 => to_signed(12774, LUT_AMPL_WIDTH),
		28592 => to_signed(12771, LUT_AMPL_WIDTH),
		28593 => to_signed(12768, LUT_AMPL_WIDTH),
		28594 => to_signed(12765, LUT_AMPL_WIDTH),
		28595 => to_signed(12763, LUT_AMPL_WIDTH),
		28596 => to_signed(12760, LUT_AMPL_WIDTH),
		28597 => to_signed(12757, LUT_AMPL_WIDTH),
		28598 => to_signed(12754, LUT_AMPL_WIDTH),
		28599 => to_signed(12751, LUT_AMPL_WIDTH),
		28600 => to_signed(12748, LUT_AMPL_WIDTH),
		28601 => to_signed(12745, LUT_AMPL_WIDTH),
		28602 => to_signed(12742, LUT_AMPL_WIDTH),
		28603 => to_signed(12739, LUT_AMPL_WIDTH),
		28604 => to_signed(12736, LUT_AMPL_WIDTH),
		28605 => to_signed(12734, LUT_AMPL_WIDTH),
		28606 => to_signed(12731, LUT_AMPL_WIDTH),
		28607 => to_signed(12728, LUT_AMPL_WIDTH),
		28608 => to_signed(12725, LUT_AMPL_WIDTH),
		28609 => to_signed(12722, LUT_AMPL_WIDTH),
		28610 => to_signed(12719, LUT_AMPL_WIDTH),
		28611 => to_signed(12716, LUT_AMPL_WIDTH),
		28612 => to_signed(12713, LUT_AMPL_WIDTH),
		28613 => to_signed(12710, LUT_AMPL_WIDTH),
		28614 => to_signed(12708, LUT_AMPL_WIDTH),
		28615 => to_signed(12705, LUT_AMPL_WIDTH),
		28616 => to_signed(12702, LUT_AMPL_WIDTH),
		28617 => to_signed(12699, LUT_AMPL_WIDTH),
		28618 => to_signed(12696, LUT_AMPL_WIDTH),
		28619 => to_signed(12693, LUT_AMPL_WIDTH),
		28620 => to_signed(12690, LUT_AMPL_WIDTH),
		28621 => to_signed(12687, LUT_AMPL_WIDTH),
		28622 => to_signed(12684, LUT_AMPL_WIDTH),
		28623 => to_signed(12681, LUT_AMPL_WIDTH),
		28624 => to_signed(12679, LUT_AMPL_WIDTH),
		28625 => to_signed(12676, LUT_AMPL_WIDTH),
		28626 => to_signed(12673, LUT_AMPL_WIDTH),
		28627 => to_signed(12670, LUT_AMPL_WIDTH),
		28628 => to_signed(12667, LUT_AMPL_WIDTH),
		28629 => to_signed(12664, LUT_AMPL_WIDTH),
		28630 => to_signed(12661, LUT_AMPL_WIDTH),
		28631 => to_signed(12658, LUT_AMPL_WIDTH),
		28632 => to_signed(12655, LUT_AMPL_WIDTH),
		28633 => to_signed(12652, LUT_AMPL_WIDTH),
		28634 => to_signed(12650, LUT_AMPL_WIDTH),
		28635 => to_signed(12647, LUT_AMPL_WIDTH),
		28636 => to_signed(12644, LUT_AMPL_WIDTH),
		28637 => to_signed(12641, LUT_AMPL_WIDTH),
		28638 => to_signed(12638, LUT_AMPL_WIDTH),
		28639 => to_signed(12635, LUT_AMPL_WIDTH),
		28640 => to_signed(12632, LUT_AMPL_WIDTH),
		28641 => to_signed(12629, LUT_AMPL_WIDTH),
		28642 => to_signed(12626, LUT_AMPL_WIDTH),
		28643 => to_signed(12624, LUT_AMPL_WIDTH),
		28644 => to_signed(12621, LUT_AMPL_WIDTH),
		28645 => to_signed(12618, LUT_AMPL_WIDTH),
		28646 => to_signed(12615, LUT_AMPL_WIDTH),
		28647 => to_signed(12612, LUT_AMPL_WIDTH),
		28648 => to_signed(12609, LUT_AMPL_WIDTH),
		28649 => to_signed(12606, LUT_AMPL_WIDTH),
		28650 => to_signed(12603, LUT_AMPL_WIDTH),
		28651 => to_signed(12600, LUT_AMPL_WIDTH),
		28652 => to_signed(12597, LUT_AMPL_WIDTH),
		28653 => to_signed(12595, LUT_AMPL_WIDTH),
		28654 => to_signed(12592, LUT_AMPL_WIDTH),
		28655 => to_signed(12589, LUT_AMPL_WIDTH),
		28656 => to_signed(12586, LUT_AMPL_WIDTH),
		28657 => to_signed(12583, LUT_AMPL_WIDTH),
		28658 => to_signed(12580, LUT_AMPL_WIDTH),
		28659 => to_signed(12577, LUT_AMPL_WIDTH),
		28660 => to_signed(12574, LUT_AMPL_WIDTH),
		28661 => to_signed(12571, LUT_AMPL_WIDTH),
		28662 => to_signed(12568, LUT_AMPL_WIDTH),
		28663 => to_signed(12566, LUT_AMPL_WIDTH),
		28664 => to_signed(12563, LUT_AMPL_WIDTH),
		28665 => to_signed(12560, LUT_AMPL_WIDTH),
		28666 => to_signed(12557, LUT_AMPL_WIDTH),
		28667 => to_signed(12554, LUT_AMPL_WIDTH),
		28668 => to_signed(12551, LUT_AMPL_WIDTH),
		28669 => to_signed(12548, LUT_AMPL_WIDTH),
		28670 => to_signed(12545, LUT_AMPL_WIDTH),
		28671 => to_signed(12542, LUT_AMPL_WIDTH),
		28672 => to_signed(12539, LUT_AMPL_WIDTH),
		28673 => to_signed(12536, LUT_AMPL_WIDTH),
		28674 => to_signed(12534, LUT_AMPL_WIDTH),
		28675 => to_signed(12531, LUT_AMPL_WIDTH),
		28676 => to_signed(12528, LUT_AMPL_WIDTH),
		28677 => to_signed(12525, LUT_AMPL_WIDTH),
		28678 => to_signed(12522, LUT_AMPL_WIDTH),
		28679 => to_signed(12519, LUT_AMPL_WIDTH),
		28680 => to_signed(12516, LUT_AMPL_WIDTH),
		28681 => to_signed(12513, LUT_AMPL_WIDTH),
		28682 => to_signed(12510, LUT_AMPL_WIDTH),
		28683 => to_signed(12507, LUT_AMPL_WIDTH),
		28684 => to_signed(12505, LUT_AMPL_WIDTH),
		28685 => to_signed(12502, LUT_AMPL_WIDTH),
		28686 => to_signed(12499, LUT_AMPL_WIDTH),
		28687 => to_signed(12496, LUT_AMPL_WIDTH),
		28688 => to_signed(12493, LUT_AMPL_WIDTH),
		28689 => to_signed(12490, LUT_AMPL_WIDTH),
		28690 => to_signed(12487, LUT_AMPL_WIDTH),
		28691 => to_signed(12484, LUT_AMPL_WIDTH),
		28692 => to_signed(12481, LUT_AMPL_WIDTH),
		28693 => to_signed(12478, LUT_AMPL_WIDTH),
		28694 => to_signed(12476, LUT_AMPL_WIDTH),
		28695 => to_signed(12473, LUT_AMPL_WIDTH),
		28696 => to_signed(12470, LUT_AMPL_WIDTH),
		28697 => to_signed(12467, LUT_AMPL_WIDTH),
		28698 => to_signed(12464, LUT_AMPL_WIDTH),
		28699 => to_signed(12461, LUT_AMPL_WIDTH),
		28700 => to_signed(12458, LUT_AMPL_WIDTH),
		28701 => to_signed(12455, LUT_AMPL_WIDTH),
		28702 => to_signed(12452, LUT_AMPL_WIDTH),
		28703 => to_signed(12449, LUT_AMPL_WIDTH),
		28704 => to_signed(12446, LUT_AMPL_WIDTH),
		28705 => to_signed(12444, LUT_AMPL_WIDTH),
		28706 => to_signed(12441, LUT_AMPL_WIDTH),
		28707 => to_signed(12438, LUT_AMPL_WIDTH),
		28708 => to_signed(12435, LUT_AMPL_WIDTH),
		28709 => to_signed(12432, LUT_AMPL_WIDTH),
		28710 => to_signed(12429, LUT_AMPL_WIDTH),
		28711 => to_signed(12426, LUT_AMPL_WIDTH),
		28712 => to_signed(12423, LUT_AMPL_WIDTH),
		28713 => to_signed(12420, LUT_AMPL_WIDTH),
		28714 => to_signed(12417, LUT_AMPL_WIDTH),
		28715 => to_signed(12414, LUT_AMPL_WIDTH),
		28716 => to_signed(12412, LUT_AMPL_WIDTH),
		28717 => to_signed(12409, LUT_AMPL_WIDTH),
		28718 => to_signed(12406, LUT_AMPL_WIDTH),
		28719 => to_signed(12403, LUT_AMPL_WIDTH),
		28720 => to_signed(12400, LUT_AMPL_WIDTH),
		28721 => to_signed(12397, LUT_AMPL_WIDTH),
		28722 => to_signed(12394, LUT_AMPL_WIDTH),
		28723 => to_signed(12391, LUT_AMPL_WIDTH),
		28724 => to_signed(12388, LUT_AMPL_WIDTH),
		28725 => to_signed(12385, LUT_AMPL_WIDTH),
		28726 => to_signed(12382, LUT_AMPL_WIDTH),
		28727 => to_signed(12380, LUT_AMPL_WIDTH),
		28728 => to_signed(12377, LUT_AMPL_WIDTH),
		28729 => to_signed(12374, LUT_AMPL_WIDTH),
		28730 => to_signed(12371, LUT_AMPL_WIDTH),
		28731 => to_signed(12368, LUT_AMPL_WIDTH),
		28732 => to_signed(12365, LUT_AMPL_WIDTH),
		28733 => to_signed(12362, LUT_AMPL_WIDTH),
		28734 => to_signed(12359, LUT_AMPL_WIDTH),
		28735 => to_signed(12356, LUT_AMPL_WIDTH),
		28736 => to_signed(12353, LUT_AMPL_WIDTH),
		28737 => to_signed(12350, LUT_AMPL_WIDTH),
		28738 => to_signed(12348, LUT_AMPL_WIDTH),
		28739 => to_signed(12345, LUT_AMPL_WIDTH),
		28740 => to_signed(12342, LUT_AMPL_WIDTH),
		28741 => to_signed(12339, LUT_AMPL_WIDTH),
		28742 => to_signed(12336, LUT_AMPL_WIDTH),
		28743 => to_signed(12333, LUT_AMPL_WIDTH),
		28744 => to_signed(12330, LUT_AMPL_WIDTH),
		28745 => to_signed(12327, LUT_AMPL_WIDTH),
		28746 => to_signed(12324, LUT_AMPL_WIDTH),
		28747 => to_signed(12321, LUT_AMPL_WIDTH),
		28748 => to_signed(12318, LUT_AMPL_WIDTH),
		28749 => to_signed(12316, LUT_AMPL_WIDTH),
		28750 => to_signed(12313, LUT_AMPL_WIDTH),
		28751 => to_signed(12310, LUT_AMPL_WIDTH),
		28752 => to_signed(12307, LUT_AMPL_WIDTH),
		28753 => to_signed(12304, LUT_AMPL_WIDTH),
		28754 => to_signed(12301, LUT_AMPL_WIDTH),
		28755 => to_signed(12298, LUT_AMPL_WIDTH),
		28756 => to_signed(12295, LUT_AMPL_WIDTH),
		28757 => to_signed(12292, LUT_AMPL_WIDTH),
		28758 => to_signed(12289, LUT_AMPL_WIDTH),
		28759 => to_signed(12286, LUT_AMPL_WIDTH),
		28760 => to_signed(12284, LUT_AMPL_WIDTH),
		28761 => to_signed(12281, LUT_AMPL_WIDTH),
		28762 => to_signed(12278, LUT_AMPL_WIDTH),
		28763 => to_signed(12275, LUT_AMPL_WIDTH),
		28764 => to_signed(12272, LUT_AMPL_WIDTH),
		28765 => to_signed(12269, LUT_AMPL_WIDTH),
		28766 => to_signed(12266, LUT_AMPL_WIDTH),
		28767 => to_signed(12263, LUT_AMPL_WIDTH),
		28768 => to_signed(12260, LUT_AMPL_WIDTH),
		28769 => to_signed(12257, LUT_AMPL_WIDTH),
		28770 => to_signed(12254, LUT_AMPL_WIDTH),
		28771 => to_signed(12251, LUT_AMPL_WIDTH),
		28772 => to_signed(12249, LUT_AMPL_WIDTH),
		28773 => to_signed(12246, LUT_AMPL_WIDTH),
		28774 => to_signed(12243, LUT_AMPL_WIDTH),
		28775 => to_signed(12240, LUT_AMPL_WIDTH),
		28776 => to_signed(12237, LUT_AMPL_WIDTH),
		28777 => to_signed(12234, LUT_AMPL_WIDTH),
		28778 => to_signed(12231, LUT_AMPL_WIDTH),
		28779 => to_signed(12228, LUT_AMPL_WIDTH),
		28780 => to_signed(12225, LUT_AMPL_WIDTH),
		28781 => to_signed(12222, LUT_AMPL_WIDTH),
		28782 => to_signed(12219, LUT_AMPL_WIDTH),
		28783 => to_signed(12217, LUT_AMPL_WIDTH),
		28784 => to_signed(12214, LUT_AMPL_WIDTH),
		28785 => to_signed(12211, LUT_AMPL_WIDTH),
		28786 => to_signed(12208, LUT_AMPL_WIDTH),
		28787 => to_signed(12205, LUT_AMPL_WIDTH),
		28788 => to_signed(12202, LUT_AMPL_WIDTH),
		28789 => to_signed(12199, LUT_AMPL_WIDTH),
		28790 => to_signed(12196, LUT_AMPL_WIDTH),
		28791 => to_signed(12193, LUT_AMPL_WIDTH),
		28792 => to_signed(12190, LUT_AMPL_WIDTH),
		28793 => to_signed(12187, LUT_AMPL_WIDTH),
		28794 => to_signed(12184, LUT_AMPL_WIDTH),
		28795 => to_signed(12182, LUT_AMPL_WIDTH),
		28796 => to_signed(12179, LUT_AMPL_WIDTH),
		28797 => to_signed(12176, LUT_AMPL_WIDTH),
		28798 => to_signed(12173, LUT_AMPL_WIDTH),
		28799 => to_signed(12170, LUT_AMPL_WIDTH),
		28800 => to_signed(12167, LUT_AMPL_WIDTH),
		28801 => to_signed(12164, LUT_AMPL_WIDTH),
		28802 => to_signed(12161, LUT_AMPL_WIDTH),
		28803 => to_signed(12158, LUT_AMPL_WIDTH),
		28804 => to_signed(12155, LUT_AMPL_WIDTH),
		28805 => to_signed(12152, LUT_AMPL_WIDTH),
		28806 => to_signed(12149, LUT_AMPL_WIDTH),
		28807 => to_signed(12147, LUT_AMPL_WIDTH),
		28808 => to_signed(12144, LUT_AMPL_WIDTH),
		28809 => to_signed(12141, LUT_AMPL_WIDTH),
		28810 => to_signed(12138, LUT_AMPL_WIDTH),
		28811 => to_signed(12135, LUT_AMPL_WIDTH),
		28812 => to_signed(12132, LUT_AMPL_WIDTH),
		28813 => to_signed(12129, LUT_AMPL_WIDTH),
		28814 => to_signed(12126, LUT_AMPL_WIDTH),
		28815 => to_signed(12123, LUT_AMPL_WIDTH),
		28816 => to_signed(12120, LUT_AMPL_WIDTH),
		28817 => to_signed(12117, LUT_AMPL_WIDTH),
		28818 => to_signed(12114, LUT_AMPL_WIDTH),
		28819 => to_signed(12112, LUT_AMPL_WIDTH),
		28820 => to_signed(12109, LUT_AMPL_WIDTH),
		28821 => to_signed(12106, LUT_AMPL_WIDTH),
		28822 => to_signed(12103, LUT_AMPL_WIDTH),
		28823 => to_signed(12100, LUT_AMPL_WIDTH),
		28824 => to_signed(12097, LUT_AMPL_WIDTH),
		28825 => to_signed(12094, LUT_AMPL_WIDTH),
		28826 => to_signed(12091, LUT_AMPL_WIDTH),
		28827 => to_signed(12088, LUT_AMPL_WIDTH),
		28828 => to_signed(12085, LUT_AMPL_WIDTH),
		28829 => to_signed(12082, LUT_AMPL_WIDTH),
		28830 => to_signed(12079, LUT_AMPL_WIDTH),
		28831 => to_signed(12076, LUT_AMPL_WIDTH),
		28832 => to_signed(12074, LUT_AMPL_WIDTH),
		28833 => to_signed(12071, LUT_AMPL_WIDTH),
		28834 => to_signed(12068, LUT_AMPL_WIDTH),
		28835 => to_signed(12065, LUT_AMPL_WIDTH),
		28836 => to_signed(12062, LUT_AMPL_WIDTH),
		28837 => to_signed(12059, LUT_AMPL_WIDTH),
		28838 => to_signed(12056, LUT_AMPL_WIDTH),
		28839 => to_signed(12053, LUT_AMPL_WIDTH),
		28840 => to_signed(12050, LUT_AMPL_WIDTH),
		28841 => to_signed(12047, LUT_AMPL_WIDTH),
		28842 => to_signed(12044, LUT_AMPL_WIDTH),
		28843 => to_signed(12041, LUT_AMPL_WIDTH),
		28844 => to_signed(12038, LUT_AMPL_WIDTH),
		28845 => to_signed(12036, LUT_AMPL_WIDTH),
		28846 => to_signed(12033, LUT_AMPL_WIDTH),
		28847 => to_signed(12030, LUT_AMPL_WIDTH),
		28848 => to_signed(12027, LUT_AMPL_WIDTH),
		28849 => to_signed(12024, LUT_AMPL_WIDTH),
		28850 => to_signed(12021, LUT_AMPL_WIDTH),
		28851 => to_signed(12018, LUT_AMPL_WIDTH),
		28852 => to_signed(12015, LUT_AMPL_WIDTH),
		28853 => to_signed(12012, LUT_AMPL_WIDTH),
		28854 => to_signed(12009, LUT_AMPL_WIDTH),
		28855 => to_signed(12006, LUT_AMPL_WIDTH),
		28856 => to_signed(12003, LUT_AMPL_WIDTH),
		28857 => to_signed(12001, LUT_AMPL_WIDTH),
		28858 => to_signed(11998, LUT_AMPL_WIDTH),
		28859 => to_signed(11995, LUT_AMPL_WIDTH),
		28860 => to_signed(11992, LUT_AMPL_WIDTH),
		28861 => to_signed(11989, LUT_AMPL_WIDTH),
		28862 => to_signed(11986, LUT_AMPL_WIDTH),
		28863 => to_signed(11983, LUT_AMPL_WIDTH),
		28864 => to_signed(11980, LUT_AMPL_WIDTH),
		28865 => to_signed(11977, LUT_AMPL_WIDTH),
		28866 => to_signed(11974, LUT_AMPL_WIDTH),
		28867 => to_signed(11971, LUT_AMPL_WIDTH),
		28868 => to_signed(11968, LUT_AMPL_WIDTH),
		28869 => to_signed(11965, LUT_AMPL_WIDTH),
		28870 => to_signed(11962, LUT_AMPL_WIDTH),
		28871 => to_signed(11960, LUT_AMPL_WIDTH),
		28872 => to_signed(11957, LUT_AMPL_WIDTH),
		28873 => to_signed(11954, LUT_AMPL_WIDTH),
		28874 => to_signed(11951, LUT_AMPL_WIDTH),
		28875 => to_signed(11948, LUT_AMPL_WIDTH),
		28876 => to_signed(11945, LUT_AMPL_WIDTH),
		28877 => to_signed(11942, LUT_AMPL_WIDTH),
		28878 => to_signed(11939, LUT_AMPL_WIDTH),
		28879 => to_signed(11936, LUT_AMPL_WIDTH),
		28880 => to_signed(11933, LUT_AMPL_WIDTH),
		28881 => to_signed(11930, LUT_AMPL_WIDTH),
		28882 => to_signed(11927, LUT_AMPL_WIDTH),
		28883 => to_signed(11924, LUT_AMPL_WIDTH),
		28884 => to_signed(11922, LUT_AMPL_WIDTH),
		28885 => to_signed(11919, LUT_AMPL_WIDTH),
		28886 => to_signed(11916, LUT_AMPL_WIDTH),
		28887 => to_signed(11913, LUT_AMPL_WIDTH),
		28888 => to_signed(11910, LUT_AMPL_WIDTH),
		28889 => to_signed(11907, LUT_AMPL_WIDTH),
		28890 => to_signed(11904, LUT_AMPL_WIDTH),
		28891 => to_signed(11901, LUT_AMPL_WIDTH),
		28892 => to_signed(11898, LUT_AMPL_WIDTH),
		28893 => to_signed(11895, LUT_AMPL_WIDTH),
		28894 => to_signed(11892, LUT_AMPL_WIDTH),
		28895 => to_signed(11889, LUT_AMPL_WIDTH),
		28896 => to_signed(11886, LUT_AMPL_WIDTH),
		28897 => to_signed(11883, LUT_AMPL_WIDTH),
		28898 => to_signed(11881, LUT_AMPL_WIDTH),
		28899 => to_signed(11878, LUT_AMPL_WIDTH),
		28900 => to_signed(11875, LUT_AMPL_WIDTH),
		28901 => to_signed(11872, LUT_AMPL_WIDTH),
		28902 => to_signed(11869, LUT_AMPL_WIDTH),
		28903 => to_signed(11866, LUT_AMPL_WIDTH),
		28904 => to_signed(11863, LUT_AMPL_WIDTH),
		28905 => to_signed(11860, LUT_AMPL_WIDTH),
		28906 => to_signed(11857, LUT_AMPL_WIDTH),
		28907 => to_signed(11854, LUT_AMPL_WIDTH),
		28908 => to_signed(11851, LUT_AMPL_WIDTH),
		28909 => to_signed(11848, LUT_AMPL_WIDTH),
		28910 => to_signed(11845, LUT_AMPL_WIDTH),
		28911 => to_signed(11842, LUT_AMPL_WIDTH),
		28912 => to_signed(11840, LUT_AMPL_WIDTH),
		28913 => to_signed(11837, LUT_AMPL_WIDTH),
		28914 => to_signed(11834, LUT_AMPL_WIDTH),
		28915 => to_signed(11831, LUT_AMPL_WIDTH),
		28916 => to_signed(11828, LUT_AMPL_WIDTH),
		28917 => to_signed(11825, LUT_AMPL_WIDTH),
		28918 => to_signed(11822, LUT_AMPL_WIDTH),
		28919 => to_signed(11819, LUT_AMPL_WIDTH),
		28920 => to_signed(11816, LUT_AMPL_WIDTH),
		28921 => to_signed(11813, LUT_AMPL_WIDTH),
		28922 => to_signed(11810, LUT_AMPL_WIDTH),
		28923 => to_signed(11807, LUT_AMPL_WIDTH),
		28924 => to_signed(11804, LUT_AMPL_WIDTH),
		28925 => to_signed(11801, LUT_AMPL_WIDTH),
		28926 => to_signed(11799, LUT_AMPL_WIDTH),
		28927 => to_signed(11796, LUT_AMPL_WIDTH),
		28928 => to_signed(11793, LUT_AMPL_WIDTH),
		28929 => to_signed(11790, LUT_AMPL_WIDTH),
		28930 => to_signed(11787, LUT_AMPL_WIDTH),
		28931 => to_signed(11784, LUT_AMPL_WIDTH),
		28932 => to_signed(11781, LUT_AMPL_WIDTH),
		28933 => to_signed(11778, LUT_AMPL_WIDTH),
		28934 => to_signed(11775, LUT_AMPL_WIDTH),
		28935 => to_signed(11772, LUT_AMPL_WIDTH),
		28936 => to_signed(11769, LUT_AMPL_WIDTH),
		28937 => to_signed(11766, LUT_AMPL_WIDTH),
		28938 => to_signed(11763, LUT_AMPL_WIDTH),
		28939 => to_signed(11760, LUT_AMPL_WIDTH),
		28940 => to_signed(11758, LUT_AMPL_WIDTH),
		28941 => to_signed(11755, LUT_AMPL_WIDTH),
		28942 => to_signed(11752, LUT_AMPL_WIDTH),
		28943 => to_signed(11749, LUT_AMPL_WIDTH),
		28944 => to_signed(11746, LUT_AMPL_WIDTH),
		28945 => to_signed(11743, LUT_AMPL_WIDTH),
		28946 => to_signed(11740, LUT_AMPL_WIDTH),
		28947 => to_signed(11737, LUT_AMPL_WIDTH),
		28948 => to_signed(11734, LUT_AMPL_WIDTH),
		28949 => to_signed(11731, LUT_AMPL_WIDTH),
		28950 => to_signed(11728, LUT_AMPL_WIDTH),
		28951 => to_signed(11725, LUT_AMPL_WIDTH),
		28952 => to_signed(11722, LUT_AMPL_WIDTH),
		28953 => to_signed(11719, LUT_AMPL_WIDTH),
		28954 => to_signed(11716, LUT_AMPL_WIDTH),
		28955 => to_signed(11714, LUT_AMPL_WIDTH),
		28956 => to_signed(11711, LUT_AMPL_WIDTH),
		28957 => to_signed(11708, LUT_AMPL_WIDTH),
		28958 => to_signed(11705, LUT_AMPL_WIDTH),
		28959 => to_signed(11702, LUT_AMPL_WIDTH),
		28960 => to_signed(11699, LUT_AMPL_WIDTH),
		28961 => to_signed(11696, LUT_AMPL_WIDTH),
		28962 => to_signed(11693, LUT_AMPL_WIDTH),
		28963 => to_signed(11690, LUT_AMPL_WIDTH),
		28964 => to_signed(11687, LUT_AMPL_WIDTH),
		28965 => to_signed(11684, LUT_AMPL_WIDTH),
		28966 => to_signed(11681, LUT_AMPL_WIDTH),
		28967 => to_signed(11678, LUT_AMPL_WIDTH),
		28968 => to_signed(11675, LUT_AMPL_WIDTH),
		28969 => to_signed(11672, LUT_AMPL_WIDTH),
		28970 => to_signed(11669, LUT_AMPL_WIDTH),
		28971 => to_signed(11667, LUT_AMPL_WIDTH),
		28972 => to_signed(11664, LUT_AMPL_WIDTH),
		28973 => to_signed(11661, LUT_AMPL_WIDTH),
		28974 => to_signed(11658, LUT_AMPL_WIDTH),
		28975 => to_signed(11655, LUT_AMPL_WIDTH),
		28976 => to_signed(11652, LUT_AMPL_WIDTH),
		28977 => to_signed(11649, LUT_AMPL_WIDTH),
		28978 => to_signed(11646, LUT_AMPL_WIDTH),
		28979 => to_signed(11643, LUT_AMPL_WIDTH),
		28980 => to_signed(11640, LUT_AMPL_WIDTH),
		28981 => to_signed(11637, LUT_AMPL_WIDTH),
		28982 => to_signed(11634, LUT_AMPL_WIDTH),
		28983 => to_signed(11631, LUT_AMPL_WIDTH),
		28984 => to_signed(11628, LUT_AMPL_WIDTH),
		28985 => to_signed(11625, LUT_AMPL_WIDTH),
		28986 => to_signed(11623, LUT_AMPL_WIDTH),
		28987 => to_signed(11620, LUT_AMPL_WIDTH),
		28988 => to_signed(11617, LUT_AMPL_WIDTH),
		28989 => to_signed(11614, LUT_AMPL_WIDTH),
		28990 => to_signed(11611, LUT_AMPL_WIDTH),
		28991 => to_signed(11608, LUT_AMPL_WIDTH),
		28992 => to_signed(11605, LUT_AMPL_WIDTH),
		28993 => to_signed(11602, LUT_AMPL_WIDTH),
		28994 => to_signed(11599, LUT_AMPL_WIDTH),
		28995 => to_signed(11596, LUT_AMPL_WIDTH),
		28996 => to_signed(11593, LUT_AMPL_WIDTH),
		28997 => to_signed(11590, LUT_AMPL_WIDTH),
		28998 => to_signed(11587, LUT_AMPL_WIDTH),
		28999 => to_signed(11584, LUT_AMPL_WIDTH),
		29000 => to_signed(11581, LUT_AMPL_WIDTH),
		29001 => to_signed(11578, LUT_AMPL_WIDTH),
		29002 => to_signed(11575, LUT_AMPL_WIDTH),
		29003 => to_signed(11573, LUT_AMPL_WIDTH),
		29004 => to_signed(11570, LUT_AMPL_WIDTH),
		29005 => to_signed(11567, LUT_AMPL_WIDTH),
		29006 => to_signed(11564, LUT_AMPL_WIDTH),
		29007 => to_signed(11561, LUT_AMPL_WIDTH),
		29008 => to_signed(11558, LUT_AMPL_WIDTH),
		29009 => to_signed(11555, LUT_AMPL_WIDTH),
		29010 => to_signed(11552, LUT_AMPL_WIDTH),
		29011 => to_signed(11549, LUT_AMPL_WIDTH),
		29012 => to_signed(11546, LUT_AMPL_WIDTH),
		29013 => to_signed(11543, LUT_AMPL_WIDTH),
		29014 => to_signed(11540, LUT_AMPL_WIDTH),
		29015 => to_signed(11537, LUT_AMPL_WIDTH),
		29016 => to_signed(11534, LUT_AMPL_WIDTH),
		29017 => to_signed(11531, LUT_AMPL_WIDTH),
		29018 => to_signed(11528, LUT_AMPL_WIDTH),
		29019 => to_signed(11526, LUT_AMPL_WIDTH),
		29020 => to_signed(11523, LUT_AMPL_WIDTH),
		29021 => to_signed(11520, LUT_AMPL_WIDTH),
		29022 => to_signed(11517, LUT_AMPL_WIDTH),
		29023 => to_signed(11514, LUT_AMPL_WIDTH),
		29024 => to_signed(11511, LUT_AMPL_WIDTH),
		29025 => to_signed(11508, LUT_AMPL_WIDTH),
		29026 => to_signed(11505, LUT_AMPL_WIDTH),
		29027 => to_signed(11502, LUT_AMPL_WIDTH),
		29028 => to_signed(11499, LUT_AMPL_WIDTH),
		29029 => to_signed(11496, LUT_AMPL_WIDTH),
		29030 => to_signed(11493, LUT_AMPL_WIDTH),
		29031 => to_signed(11490, LUT_AMPL_WIDTH),
		29032 => to_signed(11487, LUT_AMPL_WIDTH),
		29033 => to_signed(11484, LUT_AMPL_WIDTH),
		29034 => to_signed(11481, LUT_AMPL_WIDTH),
		29035 => to_signed(11478, LUT_AMPL_WIDTH),
		29036 => to_signed(11476, LUT_AMPL_WIDTH),
		29037 => to_signed(11473, LUT_AMPL_WIDTH),
		29038 => to_signed(11470, LUT_AMPL_WIDTH),
		29039 => to_signed(11467, LUT_AMPL_WIDTH),
		29040 => to_signed(11464, LUT_AMPL_WIDTH),
		29041 => to_signed(11461, LUT_AMPL_WIDTH),
		29042 => to_signed(11458, LUT_AMPL_WIDTH),
		29043 => to_signed(11455, LUT_AMPL_WIDTH),
		29044 => to_signed(11452, LUT_AMPL_WIDTH),
		29045 => to_signed(11449, LUT_AMPL_WIDTH),
		29046 => to_signed(11446, LUT_AMPL_WIDTH),
		29047 => to_signed(11443, LUT_AMPL_WIDTH),
		29048 => to_signed(11440, LUT_AMPL_WIDTH),
		29049 => to_signed(11437, LUT_AMPL_WIDTH),
		29050 => to_signed(11434, LUT_AMPL_WIDTH),
		29051 => to_signed(11431, LUT_AMPL_WIDTH),
		29052 => to_signed(11428, LUT_AMPL_WIDTH),
		29053 => to_signed(11425, LUT_AMPL_WIDTH),
		29054 => to_signed(11423, LUT_AMPL_WIDTH),
		29055 => to_signed(11420, LUT_AMPL_WIDTH),
		29056 => to_signed(11417, LUT_AMPL_WIDTH),
		29057 => to_signed(11414, LUT_AMPL_WIDTH),
		29058 => to_signed(11411, LUT_AMPL_WIDTH),
		29059 => to_signed(11408, LUT_AMPL_WIDTH),
		29060 => to_signed(11405, LUT_AMPL_WIDTH),
		29061 => to_signed(11402, LUT_AMPL_WIDTH),
		29062 => to_signed(11399, LUT_AMPL_WIDTH),
		29063 => to_signed(11396, LUT_AMPL_WIDTH),
		29064 => to_signed(11393, LUT_AMPL_WIDTH),
		29065 => to_signed(11390, LUT_AMPL_WIDTH),
		29066 => to_signed(11387, LUT_AMPL_WIDTH),
		29067 => to_signed(11384, LUT_AMPL_WIDTH),
		29068 => to_signed(11381, LUT_AMPL_WIDTH),
		29069 => to_signed(11378, LUT_AMPL_WIDTH),
		29070 => to_signed(11375, LUT_AMPL_WIDTH),
		29071 => to_signed(11372, LUT_AMPL_WIDTH),
		29072 => to_signed(11370, LUT_AMPL_WIDTH),
		29073 => to_signed(11367, LUT_AMPL_WIDTH),
		29074 => to_signed(11364, LUT_AMPL_WIDTH),
		29075 => to_signed(11361, LUT_AMPL_WIDTH),
		29076 => to_signed(11358, LUT_AMPL_WIDTH),
		29077 => to_signed(11355, LUT_AMPL_WIDTH),
		29078 => to_signed(11352, LUT_AMPL_WIDTH),
		29079 => to_signed(11349, LUT_AMPL_WIDTH),
		29080 => to_signed(11346, LUT_AMPL_WIDTH),
		29081 => to_signed(11343, LUT_AMPL_WIDTH),
		29082 => to_signed(11340, LUT_AMPL_WIDTH),
		29083 => to_signed(11337, LUT_AMPL_WIDTH),
		29084 => to_signed(11334, LUT_AMPL_WIDTH),
		29085 => to_signed(11331, LUT_AMPL_WIDTH),
		29086 => to_signed(11328, LUT_AMPL_WIDTH),
		29087 => to_signed(11325, LUT_AMPL_WIDTH),
		29088 => to_signed(11322, LUT_AMPL_WIDTH),
		29089 => to_signed(11319, LUT_AMPL_WIDTH),
		29090 => to_signed(11316, LUT_AMPL_WIDTH),
		29091 => to_signed(11314, LUT_AMPL_WIDTH),
		29092 => to_signed(11311, LUT_AMPL_WIDTH),
		29093 => to_signed(11308, LUT_AMPL_WIDTH),
		29094 => to_signed(11305, LUT_AMPL_WIDTH),
		29095 => to_signed(11302, LUT_AMPL_WIDTH),
		29096 => to_signed(11299, LUT_AMPL_WIDTH),
		29097 => to_signed(11296, LUT_AMPL_WIDTH),
		29098 => to_signed(11293, LUT_AMPL_WIDTH),
		29099 => to_signed(11290, LUT_AMPL_WIDTH),
		29100 => to_signed(11287, LUT_AMPL_WIDTH),
		29101 => to_signed(11284, LUT_AMPL_WIDTH),
		29102 => to_signed(11281, LUT_AMPL_WIDTH),
		29103 => to_signed(11278, LUT_AMPL_WIDTH),
		29104 => to_signed(11275, LUT_AMPL_WIDTH),
		29105 => to_signed(11272, LUT_AMPL_WIDTH),
		29106 => to_signed(11269, LUT_AMPL_WIDTH),
		29107 => to_signed(11266, LUT_AMPL_WIDTH),
		29108 => to_signed(11263, LUT_AMPL_WIDTH),
		29109 => to_signed(11260, LUT_AMPL_WIDTH),
		29110 => to_signed(11257, LUT_AMPL_WIDTH),
		29111 => to_signed(11255, LUT_AMPL_WIDTH),
		29112 => to_signed(11252, LUT_AMPL_WIDTH),
		29113 => to_signed(11249, LUT_AMPL_WIDTH),
		29114 => to_signed(11246, LUT_AMPL_WIDTH),
		29115 => to_signed(11243, LUT_AMPL_WIDTH),
		29116 => to_signed(11240, LUT_AMPL_WIDTH),
		29117 => to_signed(11237, LUT_AMPL_WIDTH),
		29118 => to_signed(11234, LUT_AMPL_WIDTH),
		29119 => to_signed(11231, LUT_AMPL_WIDTH),
		29120 => to_signed(11228, LUT_AMPL_WIDTH),
		29121 => to_signed(11225, LUT_AMPL_WIDTH),
		29122 => to_signed(11222, LUT_AMPL_WIDTH),
		29123 => to_signed(11219, LUT_AMPL_WIDTH),
		29124 => to_signed(11216, LUT_AMPL_WIDTH),
		29125 => to_signed(11213, LUT_AMPL_WIDTH),
		29126 => to_signed(11210, LUT_AMPL_WIDTH),
		29127 => to_signed(11207, LUT_AMPL_WIDTH),
		29128 => to_signed(11204, LUT_AMPL_WIDTH),
		29129 => to_signed(11201, LUT_AMPL_WIDTH),
		29130 => to_signed(11198, LUT_AMPL_WIDTH),
		29131 => to_signed(11195, LUT_AMPL_WIDTH),
		29132 => to_signed(11193, LUT_AMPL_WIDTH),
		29133 => to_signed(11190, LUT_AMPL_WIDTH),
		29134 => to_signed(11187, LUT_AMPL_WIDTH),
		29135 => to_signed(11184, LUT_AMPL_WIDTH),
		29136 => to_signed(11181, LUT_AMPL_WIDTH),
		29137 => to_signed(11178, LUT_AMPL_WIDTH),
		29138 => to_signed(11175, LUT_AMPL_WIDTH),
		29139 => to_signed(11172, LUT_AMPL_WIDTH),
		29140 => to_signed(11169, LUT_AMPL_WIDTH),
		29141 => to_signed(11166, LUT_AMPL_WIDTH),
		29142 => to_signed(11163, LUT_AMPL_WIDTH),
		29143 => to_signed(11160, LUT_AMPL_WIDTH),
		29144 => to_signed(11157, LUT_AMPL_WIDTH),
		29145 => to_signed(11154, LUT_AMPL_WIDTH),
		29146 => to_signed(11151, LUT_AMPL_WIDTH),
		29147 => to_signed(11148, LUT_AMPL_WIDTH),
		29148 => to_signed(11145, LUT_AMPL_WIDTH),
		29149 => to_signed(11142, LUT_AMPL_WIDTH),
		29150 => to_signed(11139, LUT_AMPL_WIDTH),
		29151 => to_signed(11136, LUT_AMPL_WIDTH),
		29152 => to_signed(11133, LUT_AMPL_WIDTH),
		29153 => to_signed(11131, LUT_AMPL_WIDTH),
		29154 => to_signed(11128, LUT_AMPL_WIDTH),
		29155 => to_signed(11125, LUT_AMPL_WIDTH),
		29156 => to_signed(11122, LUT_AMPL_WIDTH),
		29157 => to_signed(11119, LUT_AMPL_WIDTH),
		29158 => to_signed(11116, LUT_AMPL_WIDTH),
		29159 => to_signed(11113, LUT_AMPL_WIDTH),
		29160 => to_signed(11110, LUT_AMPL_WIDTH),
		29161 => to_signed(11107, LUT_AMPL_WIDTH),
		29162 => to_signed(11104, LUT_AMPL_WIDTH),
		29163 => to_signed(11101, LUT_AMPL_WIDTH),
		29164 => to_signed(11098, LUT_AMPL_WIDTH),
		29165 => to_signed(11095, LUT_AMPL_WIDTH),
		29166 => to_signed(11092, LUT_AMPL_WIDTH),
		29167 => to_signed(11089, LUT_AMPL_WIDTH),
		29168 => to_signed(11086, LUT_AMPL_WIDTH),
		29169 => to_signed(11083, LUT_AMPL_WIDTH),
		29170 => to_signed(11080, LUT_AMPL_WIDTH),
		29171 => to_signed(11077, LUT_AMPL_WIDTH),
		29172 => to_signed(11074, LUT_AMPL_WIDTH),
		29173 => to_signed(11071, LUT_AMPL_WIDTH),
		29174 => to_signed(11068, LUT_AMPL_WIDTH),
		29175 => to_signed(11065, LUT_AMPL_WIDTH),
		29176 => to_signed(11063, LUT_AMPL_WIDTH),
		29177 => to_signed(11060, LUT_AMPL_WIDTH),
		29178 => to_signed(11057, LUT_AMPL_WIDTH),
		29179 => to_signed(11054, LUT_AMPL_WIDTH),
		29180 => to_signed(11051, LUT_AMPL_WIDTH),
		29181 => to_signed(11048, LUT_AMPL_WIDTH),
		29182 => to_signed(11045, LUT_AMPL_WIDTH),
		29183 => to_signed(11042, LUT_AMPL_WIDTH),
		29184 => to_signed(11039, LUT_AMPL_WIDTH),
		29185 => to_signed(11036, LUT_AMPL_WIDTH),
		29186 => to_signed(11033, LUT_AMPL_WIDTH),
		29187 => to_signed(11030, LUT_AMPL_WIDTH),
		29188 => to_signed(11027, LUT_AMPL_WIDTH),
		29189 => to_signed(11024, LUT_AMPL_WIDTH),
		29190 => to_signed(11021, LUT_AMPL_WIDTH),
		29191 => to_signed(11018, LUT_AMPL_WIDTH),
		29192 => to_signed(11015, LUT_AMPL_WIDTH),
		29193 => to_signed(11012, LUT_AMPL_WIDTH),
		29194 => to_signed(11009, LUT_AMPL_WIDTH),
		29195 => to_signed(11006, LUT_AMPL_WIDTH),
		29196 => to_signed(11003, LUT_AMPL_WIDTH),
		29197 => to_signed(11000, LUT_AMPL_WIDTH),
		29198 => to_signed(10997, LUT_AMPL_WIDTH),
		29199 => to_signed(10994, LUT_AMPL_WIDTH),
		29200 => to_signed(10992, LUT_AMPL_WIDTH),
		29201 => to_signed(10989, LUT_AMPL_WIDTH),
		29202 => to_signed(10986, LUT_AMPL_WIDTH),
		29203 => to_signed(10983, LUT_AMPL_WIDTH),
		29204 => to_signed(10980, LUT_AMPL_WIDTH),
		29205 => to_signed(10977, LUT_AMPL_WIDTH),
		29206 => to_signed(10974, LUT_AMPL_WIDTH),
		29207 => to_signed(10971, LUT_AMPL_WIDTH),
		29208 => to_signed(10968, LUT_AMPL_WIDTH),
		29209 => to_signed(10965, LUT_AMPL_WIDTH),
		29210 => to_signed(10962, LUT_AMPL_WIDTH),
		29211 => to_signed(10959, LUT_AMPL_WIDTH),
		29212 => to_signed(10956, LUT_AMPL_WIDTH),
		29213 => to_signed(10953, LUT_AMPL_WIDTH),
		29214 => to_signed(10950, LUT_AMPL_WIDTH),
		29215 => to_signed(10947, LUT_AMPL_WIDTH),
		29216 => to_signed(10944, LUT_AMPL_WIDTH),
		29217 => to_signed(10941, LUT_AMPL_WIDTH),
		29218 => to_signed(10938, LUT_AMPL_WIDTH),
		29219 => to_signed(10935, LUT_AMPL_WIDTH),
		29220 => to_signed(10932, LUT_AMPL_WIDTH),
		29221 => to_signed(10929, LUT_AMPL_WIDTH),
		29222 => to_signed(10926, LUT_AMPL_WIDTH),
		29223 => to_signed(10923, LUT_AMPL_WIDTH),
		29224 => to_signed(10920, LUT_AMPL_WIDTH),
		29225 => to_signed(10918, LUT_AMPL_WIDTH),
		29226 => to_signed(10915, LUT_AMPL_WIDTH),
		29227 => to_signed(10912, LUT_AMPL_WIDTH),
		29228 => to_signed(10909, LUT_AMPL_WIDTH),
		29229 => to_signed(10906, LUT_AMPL_WIDTH),
		29230 => to_signed(10903, LUT_AMPL_WIDTH),
		29231 => to_signed(10900, LUT_AMPL_WIDTH),
		29232 => to_signed(10897, LUT_AMPL_WIDTH),
		29233 => to_signed(10894, LUT_AMPL_WIDTH),
		29234 => to_signed(10891, LUT_AMPL_WIDTH),
		29235 => to_signed(10888, LUT_AMPL_WIDTH),
		29236 => to_signed(10885, LUT_AMPL_WIDTH),
		29237 => to_signed(10882, LUT_AMPL_WIDTH),
		29238 => to_signed(10879, LUT_AMPL_WIDTH),
		29239 => to_signed(10876, LUT_AMPL_WIDTH),
		29240 => to_signed(10873, LUT_AMPL_WIDTH),
		29241 => to_signed(10870, LUT_AMPL_WIDTH),
		29242 => to_signed(10867, LUT_AMPL_WIDTH),
		29243 => to_signed(10864, LUT_AMPL_WIDTH),
		29244 => to_signed(10861, LUT_AMPL_WIDTH),
		29245 => to_signed(10858, LUT_AMPL_WIDTH),
		29246 => to_signed(10855, LUT_AMPL_WIDTH),
		29247 => to_signed(10852, LUT_AMPL_WIDTH),
		29248 => to_signed(10849, LUT_AMPL_WIDTH),
		29249 => to_signed(10846, LUT_AMPL_WIDTH),
		29250 => to_signed(10843, LUT_AMPL_WIDTH),
		29251 => to_signed(10840, LUT_AMPL_WIDTH),
		29252 => to_signed(10838, LUT_AMPL_WIDTH),
		29253 => to_signed(10835, LUT_AMPL_WIDTH),
		29254 => to_signed(10832, LUT_AMPL_WIDTH),
		29255 => to_signed(10829, LUT_AMPL_WIDTH),
		29256 => to_signed(10826, LUT_AMPL_WIDTH),
		29257 => to_signed(10823, LUT_AMPL_WIDTH),
		29258 => to_signed(10820, LUT_AMPL_WIDTH),
		29259 => to_signed(10817, LUT_AMPL_WIDTH),
		29260 => to_signed(10814, LUT_AMPL_WIDTH),
		29261 => to_signed(10811, LUT_AMPL_WIDTH),
		29262 => to_signed(10808, LUT_AMPL_WIDTH),
		29263 => to_signed(10805, LUT_AMPL_WIDTH),
		29264 => to_signed(10802, LUT_AMPL_WIDTH),
		29265 => to_signed(10799, LUT_AMPL_WIDTH),
		29266 => to_signed(10796, LUT_AMPL_WIDTH),
		29267 => to_signed(10793, LUT_AMPL_WIDTH),
		29268 => to_signed(10790, LUT_AMPL_WIDTH),
		29269 => to_signed(10787, LUT_AMPL_WIDTH),
		29270 => to_signed(10784, LUT_AMPL_WIDTH),
		29271 => to_signed(10781, LUT_AMPL_WIDTH),
		29272 => to_signed(10778, LUT_AMPL_WIDTH),
		29273 => to_signed(10775, LUT_AMPL_WIDTH),
		29274 => to_signed(10772, LUT_AMPL_WIDTH),
		29275 => to_signed(10769, LUT_AMPL_WIDTH),
		29276 => to_signed(10766, LUT_AMPL_WIDTH),
		29277 => to_signed(10763, LUT_AMPL_WIDTH),
		29278 => to_signed(10760, LUT_AMPL_WIDTH),
		29279 => to_signed(10757, LUT_AMPL_WIDTH),
		29280 => to_signed(10754, LUT_AMPL_WIDTH),
		29281 => to_signed(10751, LUT_AMPL_WIDTH),
		29282 => to_signed(10749, LUT_AMPL_WIDTH),
		29283 => to_signed(10746, LUT_AMPL_WIDTH),
		29284 => to_signed(10743, LUT_AMPL_WIDTH),
		29285 => to_signed(10740, LUT_AMPL_WIDTH),
		29286 => to_signed(10737, LUT_AMPL_WIDTH),
		29287 => to_signed(10734, LUT_AMPL_WIDTH),
		29288 => to_signed(10731, LUT_AMPL_WIDTH),
		29289 => to_signed(10728, LUT_AMPL_WIDTH),
		29290 => to_signed(10725, LUT_AMPL_WIDTH),
		29291 => to_signed(10722, LUT_AMPL_WIDTH),
		29292 => to_signed(10719, LUT_AMPL_WIDTH),
		29293 => to_signed(10716, LUT_AMPL_WIDTH),
		29294 => to_signed(10713, LUT_AMPL_WIDTH),
		29295 => to_signed(10710, LUT_AMPL_WIDTH),
		29296 => to_signed(10707, LUT_AMPL_WIDTH),
		29297 => to_signed(10704, LUT_AMPL_WIDTH),
		29298 => to_signed(10701, LUT_AMPL_WIDTH),
		29299 => to_signed(10698, LUT_AMPL_WIDTH),
		29300 => to_signed(10695, LUT_AMPL_WIDTH),
		29301 => to_signed(10692, LUT_AMPL_WIDTH),
		29302 => to_signed(10689, LUT_AMPL_WIDTH),
		29303 => to_signed(10686, LUT_AMPL_WIDTH),
		29304 => to_signed(10683, LUT_AMPL_WIDTH),
		29305 => to_signed(10680, LUT_AMPL_WIDTH),
		29306 => to_signed(10677, LUT_AMPL_WIDTH),
		29307 => to_signed(10674, LUT_AMPL_WIDTH),
		29308 => to_signed(10671, LUT_AMPL_WIDTH),
		29309 => to_signed(10668, LUT_AMPL_WIDTH),
		29310 => to_signed(10665, LUT_AMPL_WIDTH),
		29311 => to_signed(10662, LUT_AMPL_WIDTH),
		29312 => to_signed(10659, LUT_AMPL_WIDTH),
		29313 => to_signed(10656, LUT_AMPL_WIDTH),
		29314 => to_signed(10654, LUT_AMPL_WIDTH),
		29315 => to_signed(10651, LUT_AMPL_WIDTH),
		29316 => to_signed(10648, LUT_AMPL_WIDTH),
		29317 => to_signed(10645, LUT_AMPL_WIDTH),
		29318 => to_signed(10642, LUT_AMPL_WIDTH),
		29319 => to_signed(10639, LUT_AMPL_WIDTH),
		29320 => to_signed(10636, LUT_AMPL_WIDTH),
		29321 => to_signed(10633, LUT_AMPL_WIDTH),
		29322 => to_signed(10630, LUT_AMPL_WIDTH),
		29323 => to_signed(10627, LUT_AMPL_WIDTH),
		29324 => to_signed(10624, LUT_AMPL_WIDTH),
		29325 => to_signed(10621, LUT_AMPL_WIDTH),
		29326 => to_signed(10618, LUT_AMPL_WIDTH),
		29327 => to_signed(10615, LUT_AMPL_WIDTH),
		29328 => to_signed(10612, LUT_AMPL_WIDTH),
		29329 => to_signed(10609, LUT_AMPL_WIDTH),
		29330 => to_signed(10606, LUT_AMPL_WIDTH),
		29331 => to_signed(10603, LUT_AMPL_WIDTH),
		29332 => to_signed(10600, LUT_AMPL_WIDTH),
		29333 => to_signed(10597, LUT_AMPL_WIDTH),
		29334 => to_signed(10594, LUT_AMPL_WIDTH),
		29335 => to_signed(10591, LUT_AMPL_WIDTH),
		29336 => to_signed(10588, LUT_AMPL_WIDTH),
		29337 => to_signed(10585, LUT_AMPL_WIDTH),
		29338 => to_signed(10582, LUT_AMPL_WIDTH),
		29339 => to_signed(10579, LUT_AMPL_WIDTH),
		29340 => to_signed(10576, LUT_AMPL_WIDTH),
		29341 => to_signed(10573, LUT_AMPL_WIDTH),
		29342 => to_signed(10570, LUT_AMPL_WIDTH),
		29343 => to_signed(10567, LUT_AMPL_WIDTH),
		29344 => to_signed(10564, LUT_AMPL_WIDTH),
		29345 => to_signed(10561, LUT_AMPL_WIDTH),
		29346 => to_signed(10558, LUT_AMPL_WIDTH),
		29347 => to_signed(10555, LUT_AMPL_WIDTH),
		29348 => to_signed(10552, LUT_AMPL_WIDTH),
		29349 => to_signed(10549, LUT_AMPL_WIDTH),
		29350 => to_signed(10546, LUT_AMPL_WIDTH),
		29351 => to_signed(10544, LUT_AMPL_WIDTH),
		29352 => to_signed(10541, LUT_AMPL_WIDTH),
		29353 => to_signed(10538, LUT_AMPL_WIDTH),
		29354 => to_signed(10535, LUT_AMPL_WIDTH),
		29355 => to_signed(10532, LUT_AMPL_WIDTH),
		29356 => to_signed(10529, LUT_AMPL_WIDTH),
		29357 => to_signed(10526, LUT_AMPL_WIDTH),
		29358 => to_signed(10523, LUT_AMPL_WIDTH),
		29359 => to_signed(10520, LUT_AMPL_WIDTH),
		29360 => to_signed(10517, LUT_AMPL_WIDTH),
		29361 => to_signed(10514, LUT_AMPL_WIDTH),
		29362 => to_signed(10511, LUT_AMPL_WIDTH),
		29363 => to_signed(10508, LUT_AMPL_WIDTH),
		29364 => to_signed(10505, LUT_AMPL_WIDTH),
		29365 => to_signed(10502, LUT_AMPL_WIDTH),
		29366 => to_signed(10499, LUT_AMPL_WIDTH),
		29367 => to_signed(10496, LUT_AMPL_WIDTH),
		29368 => to_signed(10493, LUT_AMPL_WIDTH),
		29369 => to_signed(10490, LUT_AMPL_WIDTH),
		29370 => to_signed(10487, LUT_AMPL_WIDTH),
		29371 => to_signed(10484, LUT_AMPL_WIDTH),
		29372 => to_signed(10481, LUT_AMPL_WIDTH),
		29373 => to_signed(10478, LUT_AMPL_WIDTH),
		29374 => to_signed(10475, LUT_AMPL_WIDTH),
		29375 => to_signed(10472, LUT_AMPL_WIDTH),
		29376 => to_signed(10469, LUT_AMPL_WIDTH),
		29377 => to_signed(10466, LUT_AMPL_WIDTH),
		29378 => to_signed(10463, LUT_AMPL_WIDTH),
		29379 => to_signed(10460, LUT_AMPL_WIDTH),
		29380 => to_signed(10457, LUT_AMPL_WIDTH),
		29381 => to_signed(10454, LUT_AMPL_WIDTH),
		29382 => to_signed(10451, LUT_AMPL_WIDTH),
		29383 => to_signed(10448, LUT_AMPL_WIDTH),
		29384 => to_signed(10445, LUT_AMPL_WIDTH),
		29385 => to_signed(10442, LUT_AMPL_WIDTH),
		29386 => to_signed(10439, LUT_AMPL_WIDTH),
		29387 => to_signed(10436, LUT_AMPL_WIDTH),
		29388 => to_signed(10433, LUT_AMPL_WIDTH),
		29389 => to_signed(10430, LUT_AMPL_WIDTH),
		29390 => to_signed(10427, LUT_AMPL_WIDTH),
		29391 => to_signed(10424, LUT_AMPL_WIDTH),
		29392 => to_signed(10421, LUT_AMPL_WIDTH),
		29393 => to_signed(10419, LUT_AMPL_WIDTH),
		29394 => to_signed(10416, LUT_AMPL_WIDTH),
		29395 => to_signed(10413, LUT_AMPL_WIDTH),
		29396 => to_signed(10410, LUT_AMPL_WIDTH),
		29397 => to_signed(10407, LUT_AMPL_WIDTH),
		29398 => to_signed(10404, LUT_AMPL_WIDTH),
		29399 => to_signed(10401, LUT_AMPL_WIDTH),
		29400 => to_signed(10398, LUT_AMPL_WIDTH),
		29401 => to_signed(10395, LUT_AMPL_WIDTH),
		29402 => to_signed(10392, LUT_AMPL_WIDTH),
		29403 => to_signed(10389, LUT_AMPL_WIDTH),
		29404 => to_signed(10386, LUT_AMPL_WIDTH),
		29405 => to_signed(10383, LUT_AMPL_WIDTH),
		29406 => to_signed(10380, LUT_AMPL_WIDTH),
		29407 => to_signed(10377, LUT_AMPL_WIDTH),
		29408 => to_signed(10374, LUT_AMPL_WIDTH),
		29409 => to_signed(10371, LUT_AMPL_WIDTH),
		29410 => to_signed(10368, LUT_AMPL_WIDTH),
		29411 => to_signed(10365, LUT_AMPL_WIDTH),
		29412 => to_signed(10362, LUT_AMPL_WIDTH),
		29413 => to_signed(10359, LUT_AMPL_WIDTH),
		29414 => to_signed(10356, LUT_AMPL_WIDTH),
		29415 => to_signed(10353, LUT_AMPL_WIDTH),
		29416 => to_signed(10350, LUT_AMPL_WIDTH),
		29417 => to_signed(10347, LUT_AMPL_WIDTH),
		29418 => to_signed(10344, LUT_AMPL_WIDTH),
		29419 => to_signed(10341, LUT_AMPL_WIDTH),
		29420 => to_signed(10338, LUT_AMPL_WIDTH),
		29421 => to_signed(10335, LUT_AMPL_WIDTH),
		29422 => to_signed(10332, LUT_AMPL_WIDTH),
		29423 => to_signed(10329, LUT_AMPL_WIDTH),
		29424 => to_signed(10326, LUT_AMPL_WIDTH),
		29425 => to_signed(10323, LUT_AMPL_WIDTH),
		29426 => to_signed(10320, LUT_AMPL_WIDTH),
		29427 => to_signed(10317, LUT_AMPL_WIDTH),
		29428 => to_signed(10314, LUT_AMPL_WIDTH),
		29429 => to_signed(10311, LUT_AMPL_WIDTH),
		29430 => to_signed(10308, LUT_AMPL_WIDTH),
		29431 => to_signed(10305, LUT_AMPL_WIDTH),
		29432 => to_signed(10302, LUT_AMPL_WIDTH),
		29433 => to_signed(10299, LUT_AMPL_WIDTH),
		29434 => to_signed(10296, LUT_AMPL_WIDTH),
		29435 => to_signed(10293, LUT_AMPL_WIDTH),
		29436 => to_signed(10290, LUT_AMPL_WIDTH),
		29437 => to_signed(10287, LUT_AMPL_WIDTH),
		29438 => to_signed(10284, LUT_AMPL_WIDTH),
		29439 => to_signed(10281, LUT_AMPL_WIDTH),
		29440 => to_signed(10278, LUT_AMPL_WIDTH),
		29441 => to_signed(10275, LUT_AMPL_WIDTH),
		29442 => to_signed(10272, LUT_AMPL_WIDTH),
		29443 => to_signed(10269, LUT_AMPL_WIDTH),
		29444 => to_signed(10266, LUT_AMPL_WIDTH),
		29445 => to_signed(10263, LUT_AMPL_WIDTH),
		29446 => to_signed(10261, LUT_AMPL_WIDTH),
		29447 => to_signed(10258, LUT_AMPL_WIDTH),
		29448 => to_signed(10255, LUT_AMPL_WIDTH),
		29449 => to_signed(10252, LUT_AMPL_WIDTH),
		29450 => to_signed(10249, LUT_AMPL_WIDTH),
		29451 => to_signed(10246, LUT_AMPL_WIDTH),
		29452 => to_signed(10243, LUT_AMPL_WIDTH),
		29453 => to_signed(10240, LUT_AMPL_WIDTH),
		29454 => to_signed(10237, LUT_AMPL_WIDTH),
		29455 => to_signed(10234, LUT_AMPL_WIDTH),
		29456 => to_signed(10231, LUT_AMPL_WIDTH),
		29457 => to_signed(10228, LUT_AMPL_WIDTH),
		29458 => to_signed(10225, LUT_AMPL_WIDTH),
		29459 => to_signed(10222, LUT_AMPL_WIDTH),
		29460 => to_signed(10219, LUT_AMPL_WIDTH),
		29461 => to_signed(10216, LUT_AMPL_WIDTH),
		29462 => to_signed(10213, LUT_AMPL_WIDTH),
		29463 => to_signed(10210, LUT_AMPL_WIDTH),
		29464 => to_signed(10207, LUT_AMPL_WIDTH),
		29465 => to_signed(10204, LUT_AMPL_WIDTH),
		29466 => to_signed(10201, LUT_AMPL_WIDTH),
		29467 => to_signed(10198, LUT_AMPL_WIDTH),
		29468 => to_signed(10195, LUT_AMPL_WIDTH),
		29469 => to_signed(10192, LUT_AMPL_WIDTH),
		29470 => to_signed(10189, LUT_AMPL_WIDTH),
		29471 => to_signed(10186, LUT_AMPL_WIDTH),
		29472 => to_signed(10183, LUT_AMPL_WIDTH),
		29473 => to_signed(10180, LUT_AMPL_WIDTH),
		29474 => to_signed(10177, LUT_AMPL_WIDTH),
		29475 => to_signed(10174, LUT_AMPL_WIDTH),
		29476 => to_signed(10171, LUT_AMPL_WIDTH),
		29477 => to_signed(10168, LUT_AMPL_WIDTH),
		29478 => to_signed(10165, LUT_AMPL_WIDTH),
		29479 => to_signed(10162, LUT_AMPL_WIDTH),
		29480 => to_signed(10159, LUT_AMPL_WIDTH),
		29481 => to_signed(10156, LUT_AMPL_WIDTH),
		29482 => to_signed(10153, LUT_AMPL_WIDTH),
		29483 => to_signed(10150, LUT_AMPL_WIDTH),
		29484 => to_signed(10147, LUT_AMPL_WIDTH),
		29485 => to_signed(10144, LUT_AMPL_WIDTH),
		29486 => to_signed(10141, LUT_AMPL_WIDTH),
		29487 => to_signed(10138, LUT_AMPL_WIDTH),
		29488 => to_signed(10135, LUT_AMPL_WIDTH),
		29489 => to_signed(10132, LUT_AMPL_WIDTH),
		29490 => to_signed(10129, LUT_AMPL_WIDTH),
		29491 => to_signed(10126, LUT_AMPL_WIDTH),
		29492 => to_signed(10123, LUT_AMPL_WIDTH),
		29493 => to_signed(10120, LUT_AMPL_WIDTH),
		29494 => to_signed(10117, LUT_AMPL_WIDTH),
		29495 => to_signed(10114, LUT_AMPL_WIDTH),
		29496 => to_signed(10111, LUT_AMPL_WIDTH),
		29497 => to_signed(10108, LUT_AMPL_WIDTH),
		29498 => to_signed(10105, LUT_AMPL_WIDTH),
		29499 => to_signed(10102, LUT_AMPL_WIDTH),
		29500 => to_signed(10099, LUT_AMPL_WIDTH),
		29501 => to_signed(10096, LUT_AMPL_WIDTH),
		29502 => to_signed(10093, LUT_AMPL_WIDTH),
		29503 => to_signed(10090, LUT_AMPL_WIDTH),
		29504 => to_signed(10087, LUT_AMPL_WIDTH),
		29505 => to_signed(10084, LUT_AMPL_WIDTH),
		29506 => to_signed(10081, LUT_AMPL_WIDTH),
		29507 => to_signed(10078, LUT_AMPL_WIDTH),
		29508 => to_signed(10075, LUT_AMPL_WIDTH),
		29509 => to_signed(10072, LUT_AMPL_WIDTH),
		29510 => to_signed(10069, LUT_AMPL_WIDTH),
		29511 => to_signed(10066, LUT_AMPL_WIDTH),
		29512 => to_signed(10063, LUT_AMPL_WIDTH),
		29513 => to_signed(10060, LUT_AMPL_WIDTH),
		29514 => to_signed(10057, LUT_AMPL_WIDTH),
		29515 => to_signed(10054, LUT_AMPL_WIDTH),
		29516 => to_signed(10051, LUT_AMPL_WIDTH),
		29517 => to_signed(10048, LUT_AMPL_WIDTH),
		29518 => to_signed(10045, LUT_AMPL_WIDTH),
		29519 => to_signed(10042, LUT_AMPL_WIDTH),
		29520 => to_signed(10039, LUT_AMPL_WIDTH),
		29521 => to_signed(10036, LUT_AMPL_WIDTH),
		29522 => to_signed(10033, LUT_AMPL_WIDTH),
		29523 => to_signed(10031, LUT_AMPL_WIDTH),
		29524 => to_signed(10028, LUT_AMPL_WIDTH),
		29525 => to_signed(10025, LUT_AMPL_WIDTH),
		29526 => to_signed(10022, LUT_AMPL_WIDTH),
		29527 => to_signed(10019, LUT_AMPL_WIDTH),
		29528 => to_signed(10016, LUT_AMPL_WIDTH),
		29529 => to_signed(10013, LUT_AMPL_WIDTH),
		29530 => to_signed(10010, LUT_AMPL_WIDTH),
		29531 => to_signed(10007, LUT_AMPL_WIDTH),
		29532 => to_signed(10004, LUT_AMPL_WIDTH),
		29533 => to_signed(10001, LUT_AMPL_WIDTH),
		29534 => to_signed(9998, LUT_AMPL_WIDTH),
		29535 => to_signed(9995, LUT_AMPL_WIDTH),
		29536 => to_signed(9992, LUT_AMPL_WIDTH),
		29537 => to_signed(9989, LUT_AMPL_WIDTH),
		29538 => to_signed(9986, LUT_AMPL_WIDTH),
		29539 => to_signed(9983, LUT_AMPL_WIDTH),
		29540 => to_signed(9980, LUT_AMPL_WIDTH),
		29541 => to_signed(9977, LUT_AMPL_WIDTH),
		29542 => to_signed(9974, LUT_AMPL_WIDTH),
		29543 => to_signed(9971, LUT_AMPL_WIDTH),
		29544 => to_signed(9968, LUT_AMPL_WIDTH),
		29545 => to_signed(9965, LUT_AMPL_WIDTH),
		29546 => to_signed(9962, LUT_AMPL_WIDTH),
		29547 => to_signed(9959, LUT_AMPL_WIDTH),
		29548 => to_signed(9956, LUT_AMPL_WIDTH),
		29549 => to_signed(9953, LUT_AMPL_WIDTH),
		29550 => to_signed(9950, LUT_AMPL_WIDTH),
		29551 => to_signed(9947, LUT_AMPL_WIDTH),
		29552 => to_signed(9944, LUT_AMPL_WIDTH),
		29553 => to_signed(9941, LUT_AMPL_WIDTH),
		29554 => to_signed(9938, LUT_AMPL_WIDTH),
		29555 => to_signed(9935, LUT_AMPL_WIDTH),
		29556 => to_signed(9932, LUT_AMPL_WIDTH),
		29557 => to_signed(9929, LUT_AMPL_WIDTH),
		29558 => to_signed(9926, LUT_AMPL_WIDTH),
		29559 => to_signed(9923, LUT_AMPL_WIDTH),
		29560 => to_signed(9920, LUT_AMPL_WIDTH),
		29561 => to_signed(9917, LUT_AMPL_WIDTH),
		29562 => to_signed(9914, LUT_AMPL_WIDTH),
		29563 => to_signed(9911, LUT_AMPL_WIDTH),
		29564 => to_signed(9908, LUT_AMPL_WIDTH),
		29565 => to_signed(9905, LUT_AMPL_WIDTH),
		29566 => to_signed(9902, LUT_AMPL_WIDTH),
		29567 => to_signed(9899, LUT_AMPL_WIDTH),
		29568 => to_signed(9896, LUT_AMPL_WIDTH),
		29569 => to_signed(9893, LUT_AMPL_WIDTH),
		29570 => to_signed(9890, LUT_AMPL_WIDTH),
		29571 => to_signed(9887, LUT_AMPL_WIDTH),
		29572 => to_signed(9884, LUT_AMPL_WIDTH),
		29573 => to_signed(9881, LUT_AMPL_WIDTH),
		29574 => to_signed(9878, LUT_AMPL_WIDTH),
		29575 => to_signed(9875, LUT_AMPL_WIDTH),
		29576 => to_signed(9872, LUT_AMPL_WIDTH),
		29577 => to_signed(9869, LUT_AMPL_WIDTH),
		29578 => to_signed(9866, LUT_AMPL_WIDTH),
		29579 => to_signed(9863, LUT_AMPL_WIDTH),
		29580 => to_signed(9860, LUT_AMPL_WIDTH),
		29581 => to_signed(9857, LUT_AMPL_WIDTH),
		29582 => to_signed(9854, LUT_AMPL_WIDTH),
		29583 => to_signed(9851, LUT_AMPL_WIDTH),
		29584 => to_signed(9848, LUT_AMPL_WIDTH),
		29585 => to_signed(9845, LUT_AMPL_WIDTH),
		29586 => to_signed(9842, LUT_AMPL_WIDTH),
		29587 => to_signed(9839, LUT_AMPL_WIDTH),
		29588 => to_signed(9836, LUT_AMPL_WIDTH),
		29589 => to_signed(9833, LUT_AMPL_WIDTH),
		29590 => to_signed(9830, LUT_AMPL_WIDTH),
		29591 => to_signed(9827, LUT_AMPL_WIDTH),
		29592 => to_signed(9824, LUT_AMPL_WIDTH),
		29593 => to_signed(9821, LUT_AMPL_WIDTH),
		29594 => to_signed(9818, LUT_AMPL_WIDTH),
		29595 => to_signed(9815, LUT_AMPL_WIDTH),
		29596 => to_signed(9812, LUT_AMPL_WIDTH),
		29597 => to_signed(9809, LUT_AMPL_WIDTH),
		29598 => to_signed(9806, LUT_AMPL_WIDTH),
		29599 => to_signed(9803, LUT_AMPL_WIDTH),
		29600 => to_signed(9800, LUT_AMPL_WIDTH),
		29601 => to_signed(9797, LUT_AMPL_WIDTH),
		29602 => to_signed(9794, LUT_AMPL_WIDTH),
		29603 => to_signed(9791, LUT_AMPL_WIDTH),
		29604 => to_signed(9788, LUT_AMPL_WIDTH),
		29605 => to_signed(9785, LUT_AMPL_WIDTH),
		29606 => to_signed(9782, LUT_AMPL_WIDTH),
		29607 => to_signed(9779, LUT_AMPL_WIDTH),
		29608 => to_signed(9776, LUT_AMPL_WIDTH),
		29609 => to_signed(9773, LUT_AMPL_WIDTH),
		29610 => to_signed(9770, LUT_AMPL_WIDTH),
		29611 => to_signed(9767, LUT_AMPL_WIDTH),
		29612 => to_signed(9764, LUT_AMPL_WIDTH),
		29613 => to_signed(9761, LUT_AMPL_WIDTH),
		29614 => to_signed(9758, LUT_AMPL_WIDTH),
		29615 => to_signed(9755, LUT_AMPL_WIDTH),
		29616 => to_signed(9752, LUT_AMPL_WIDTH),
		29617 => to_signed(9749, LUT_AMPL_WIDTH),
		29618 => to_signed(9746, LUT_AMPL_WIDTH),
		29619 => to_signed(9743, LUT_AMPL_WIDTH),
		29620 => to_signed(9740, LUT_AMPL_WIDTH),
		29621 => to_signed(9737, LUT_AMPL_WIDTH),
		29622 => to_signed(9734, LUT_AMPL_WIDTH),
		29623 => to_signed(9731, LUT_AMPL_WIDTH),
		29624 => to_signed(9728, LUT_AMPL_WIDTH),
		29625 => to_signed(9725, LUT_AMPL_WIDTH),
		29626 => to_signed(9722, LUT_AMPL_WIDTH),
		29627 => to_signed(9719, LUT_AMPL_WIDTH),
		29628 => to_signed(9716, LUT_AMPL_WIDTH),
		29629 => to_signed(9713, LUT_AMPL_WIDTH),
		29630 => to_signed(9710, LUT_AMPL_WIDTH),
		29631 => to_signed(9707, LUT_AMPL_WIDTH),
		29632 => to_signed(9704, LUT_AMPL_WIDTH),
		29633 => to_signed(9701, LUT_AMPL_WIDTH),
		29634 => to_signed(9698, LUT_AMPL_WIDTH),
		29635 => to_signed(9695, LUT_AMPL_WIDTH),
		29636 => to_signed(9692, LUT_AMPL_WIDTH),
		29637 => to_signed(9689, LUT_AMPL_WIDTH),
		29638 => to_signed(9686, LUT_AMPL_WIDTH),
		29639 => to_signed(9683, LUT_AMPL_WIDTH),
		29640 => to_signed(9680, LUT_AMPL_WIDTH),
		29641 => to_signed(9677, LUT_AMPL_WIDTH),
		29642 => to_signed(9674, LUT_AMPL_WIDTH),
		29643 => to_signed(9671, LUT_AMPL_WIDTH),
		29644 => to_signed(9668, LUT_AMPL_WIDTH),
		29645 => to_signed(9665, LUT_AMPL_WIDTH),
		29646 => to_signed(9662, LUT_AMPL_WIDTH),
		29647 => to_signed(9659, LUT_AMPL_WIDTH),
		29648 => to_signed(9656, LUT_AMPL_WIDTH),
		29649 => to_signed(9653, LUT_AMPL_WIDTH),
		29650 => to_signed(9650, LUT_AMPL_WIDTH),
		29651 => to_signed(9647, LUT_AMPL_WIDTH),
		29652 => to_signed(9644, LUT_AMPL_WIDTH),
		29653 => to_signed(9641, LUT_AMPL_WIDTH),
		29654 => to_signed(9638, LUT_AMPL_WIDTH),
		29655 => to_signed(9635, LUT_AMPL_WIDTH),
		29656 => to_signed(9632, LUT_AMPL_WIDTH),
		29657 => to_signed(9629, LUT_AMPL_WIDTH),
		29658 => to_signed(9626, LUT_AMPL_WIDTH),
		29659 => to_signed(9623, LUT_AMPL_WIDTH),
		29660 => to_signed(9620, LUT_AMPL_WIDTH),
		29661 => to_signed(9617, LUT_AMPL_WIDTH),
		29662 => to_signed(9614, LUT_AMPL_WIDTH),
		29663 => to_signed(9611, LUT_AMPL_WIDTH),
		29664 => to_signed(9608, LUT_AMPL_WIDTH),
		29665 => to_signed(9605, LUT_AMPL_WIDTH),
		29666 => to_signed(9602, LUT_AMPL_WIDTH),
		29667 => to_signed(9599, LUT_AMPL_WIDTH),
		29668 => to_signed(9596, LUT_AMPL_WIDTH),
		29669 => to_signed(9593, LUT_AMPL_WIDTH),
		29670 => to_signed(9590, LUT_AMPL_WIDTH),
		29671 => to_signed(9587, LUT_AMPL_WIDTH),
		29672 => to_signed(9584, LUT_AMPL_WIDTH),
		29673 => to_signed(9581, LUT_AMPL_WIDTH),
		29674 => to_signed(9578, LUT_AMPL_WIDTH),
		29675 => to_signed(9575, LUT_AMPL_WIDTH),
		29676 => to_signed(9572, LUT_AMPL_WIDTH),
		29677 => to_signed(9569, LUT_AMPL_WIDTH),
		29678 => to_signed(9566, LUT_AMPL_WIDTH),
		29679 => to_signed(9563, LUT_AMPL_WIDTH),
		29680 => to_signed(9560, LUT_AMPL_WIDTH),
		29681 => to_signed(9557, LUT_AMPL_WIDTH),
		29682 => to_signed(9554, LUT_AMPL_WIDTH),
		29683 => to_signed(9551, LUT_AMPL_WIDTH),
		29684 => to_signed(9548, LUT_AMPL_WIDTH),
		29685 => to_signed(9545, LUT_AMPL_WIDTH),
		29686 => to_signed(9542, LUT_AMPL_WIDTH),
		29687 => to_signed(9539, LUT_AMPL_WIDTH),
		29688 => to_signed(9536, LUT_AMPL_WIDTH),
		29689 => to_signed(9533, LUT_AMPL_WIDTH),
		29690 => to_signed(9530, LUT_AMPL_WIDTH),
		29691 => to_signed(9527, LUT_AMPL_WIDTH),
		29692 => to_signed(9524, LUT_AMPL_WIDTH),
		29693 => to_signed(9521, LUT_AMPL_WIDTH),
		29694 => to_signed(9518, LUT_AMPL_WIDTH),
		29695 => to_signed(9515, LUT_AMPL_WIDTH),
		29696 => to_signed(9512, LUT_AMPL_WIDTH),
		29697 => to_signed(9509, LUT_AMPL_WIDTH),
		29698 => to_signed(9506, LUT_AMPL_WIDTH),
		29699 => to_signed(9503, LUT_AMPL_WIDTH),
		29700 => to_signed(9500, LUT_AMPL_WIDTH),
		29701 => to_signed(9497, LUT_AMPL_WIDTH),
		29702 => to_signed(9494, LUT_AMPL_WIDTH),
		29703 => to_signed(9491, LUT_AMPL_WIDTH),
		29704 => to_signed(9488, LUT_AMPL_WIDTH),
		29705 => to_signed(9485, LUT_AMPL_WIDTH),
		29706 => to_signed(9482, LUT_AMPL_WIDTH),
		29707 => to_signed(9479, LUT_AMPL_WIDTH),
		29708 => to_signed(9476, LUT_AMPL_WIDTH),
		29709 => to_signed(9473, LUT_AMPL_WIDTH),
		29710 => to_signed(9470, LUT_AMPL_WIDTH),
		29711 => to_signed(9467, LUT_AMPL_WIDTH),
		29712 => to_signed(9464, LUT_AMPL_WIDTH),
		29713 => to_signed(9461, LUT_AMPL_WIDTH),
		29714 => to_signed(9458, LUT_AMPL_WIDTH),
		29715 => to_signed(9455, LUT_AMPL_WIDTH),
		29716 => to_signed(9452, LUT_AMPL_WIDTH),
		29717 => to_signed(9449, LUT_AMPL_WIDTH),
		29718 => to_signed(9446, LUT_AMPL_WIDTH),
		29719 => to_signed(9443, LUT_AMPL_WIDTH),
		29720 => to_signed(9440, LUT_AMPL_WIDTH),
		29721 => to_signed(9437, LUT_AMPL_WIDTH),
		29722 => to_signed(9434, LUT_AMPL_WIDTH),
		29723 => to_signed(9431, LUT_AMPL_WIDTH),
		29724 => to_signed(9428, LUT_AMPL_WIDTH),
		29725 => to_signed(9425, LUT_AMPL_WIDTH),
		29726 => to_signed(9422, LUT_AMPL_WIDTH),
		29727 => to_signed(9419, LUT_AMPL_WIDTH),
		29728 => to_signed(9416, LUT_AMPL_WIDTH),
		29729 => to_signed(9413, LUT_AMPL_WIDTH),
		29730 => to_signed(9409, LUT_AMPL_WIDTH),
		29731 => to_signed(9406, LUT_AMPL_WIDTH),
		29732 => to_signed(9403, LUT_AMPL_WIDTH),
		29733 => to_signed(9400, LUT_AMPL_WIDTH),
		29734 => to_signed(9397, LUT_AMPL_WIDTH),
		29735 => to_signed(9394, LUT_AMPL_WIDTH),
		29736 => to_signed(9391, LUT_AMPL_WIDTH),
		29737 => to_signed(9388, LUT_AMPL_WIDTH),
		29738 => to_signed(9385, LUT_AMPL_WIDTH),
		29739 => to_signed(9382, LUT_AMPL_WIDTH),
		29740 => to_signed(9379, LUT_AMPL_WIDTH),
		29741 => to_signed(9376, LUT_AMPL_WIDTH),
		29742 => to_signed(9373, LUT_AMPL_WIDTH),
		29743 => to_signed(9370, LUT_AMPL_WIDTH),
		29744 => to_signed(9367, LUT_AMPL_WIDTH),
		29745 => to_signed(9364, LUT_AMPL_WIDTH),
		29746 => to_signed(9361, LUT_AMPL_WIDTH),
		29747 => to_signed(9358, LUT_AMPL_WIDTH),
		29748 => to_signed(9355, LUT_AMPL_WIDTH),
		29749 => to_signed(9352, LUT_AMPL_WIDTH),
		29750 => to_signed(9349, LUT_AMPL_WIDTH),
		29751 => to_signed(9346, LUT_AMPL_WIDTH),
		29752 => to_signed(9343, LUT_AMPL_WIDTH),
		29753 => to_signed(9340, LUT_AMPL_WIDTH),
		29754 => to_signed(9337, LUT_AMPL_WIDTH),
		29755 => to_signed(9334, LUT_AMPL_WIDTH),
		29756 => to_signed(9331, LUT_AMPL_WIDTH),
		29757 => to_signed(9328, LUT_AMPL_WIDTH),
		29758 => to_signed(9325, LUT_AMPL_WIDTH),
		29759 => to_signed(9322, LUT_AMPL_WIDTH),
		29760 => to_signed(9319, LUT_AMPL_WIDTH),
		29761 => to_signed(9316, LUT_AMPL_WIDTH),
		29762 => to_signed(9313, LUT_AMPL_WIDTH),
		29763 => to_signed(9310, LUT_AMPL_WIDTH),
		29764 => to_signed(9307, LUT_AMPL_WIDTH),
		29765 => to_signed(9304, LUT_AMPL_WIDTH),
		29766 => to_signed(9301, LUT_AMPL_WIDTH),
		29767 => to_signed(9298, LUT_AMPL_WIDTH),
		29768 => to_signed(9295, LUT_AMPL_WIDTH),
		29769 => to_signed(9292, LUT_AMPL_WIDTH),
		29770 => to_signed(9289, LUT_AMPL_WIDTH),
		29771 => to_signed(9286, LUT_AMPL_WIDTH),
		29772 => to_signed(9283, LUT_AMPL_WIDTH),
		29773 => to_signed(9280, LUT_AMPL_WIDTH),
		29774 => to_signed(9277, LUT_AMPL_WIDTH),
		29775 => to_signed(9274, LUT_AMPL_WIDTH),
		29776 => to_signed(9271, LUT_AMPL_WIDTH),
		29777 => to_signed(9268, LUT_AMPL_WIDTH),
		29778 => to_signed(9265, LUT_AMPL_WIDTH),
		29779 => to_signed(9262, LUT_AMPL_WIDTH),
		29780 => to_signed(9259, LUT_AMPL_WIDTH),
		29781 => to_signed(9256, LUT_AMPL_WIDTH),
		29782 => to_signed(9253, LUT_AMPL_WIDTH),
		29783 => to_signed(9250, LUT_AMPL_WIDTH),
		29784 => to_signed(9247, LUT_AMPL_WIDTH),
		29785 => to_signed(9244, LUT_AMPL_WIDTH),
		29786 => to_signed(9241, LUT_AMPL_WIDTH),
		29787 => to_signed(9238, LUT_AMPL_WIDTH),
		29788 => to_signed(9235, LUT_AMPL_WIDTH),
		29789 => to_signed(9232, LUT_AMPL_WIDTH),
		29790 => to_signed(9229, LUT_AMPL_WIDTH),
		29791 => to_signed(9226, LUT_AMPL_WIDTH),
		29792 => to_signed(9223, LUT_AMPL_WIDTH),
		29793 => to_signed(9220, LUT_AMPL_WIDTH),
		29794 => to_signed(9217, LUT_AMPL_WIDTH),
		29795 => to_signed(9214, LUT_AMPL_WIDTH),
		29796 => to_signed(9211, LUT_AMPL_WIDTH),
		29797 => to_signed(9208, LUT_AMPL_WIDTH),
		29798 => to_signed(9205, LUT_AMPL_WIDTH),
		29799 => to_signed(9202, LUT_AMPL_WIDTH),
		29800 => to_signed(9199, LUT_AMPL_WIDTH),
		29801 => to_signed(9196, LUT_AMPL_WIDTH),
		29802 => to_signed(9193, LUT_AMPL_WIDTH),
		29803 => to_signed(9190, LUT_AMPL_WIDTH),
		29804 => to_signed(9187, LUT_AMPL_WIDTH),
		29805 => to_signed(9184, LUT_AMPL_WIDTH),
		29806 => to_signed(9181, LUT_AMPL_WIDTH),
		29807 => to_signed(9178, LUT_AMPL_WIDTH),
		29808 => to_signed(9175, LUT_AMPL_WIDTH),
		29809 => to_signed(9172, LUT_AMPL_WIDTH),
		29810 => to_signed(9168, LUT_AMPL_WIDTH),
		29811 => to_signed(9165, LUT_AMPL_WIDTH),
		29812 => to_signed(9162, LUT_AMPL_WIDTH),
		29813 => to_signed(9159, LUT_AMPL_WIDTH),
		29814 => to_signed(9156, LUT_AMPL_WIDTH),
		29815 => to_signed(9153, LUT_AMPL_WIDTH),
		29816 => to_signed(9150, LUT_AMPL_WIDTH),
		29817 => to_signed(9147, LUT_AMPL_WIDTH),
		29818 => to_signed(9144, LUT_AMPL_WIDTH),
		29819 => to_signed(9141, LUT_AMPL_WIDTH),
		29820 => to_signed(9138, LUT_AMPL_WIDTH),
		29821 => to_signed(9135, LUT_AMPL_WIDTH),
		29822 => to_signed(9132, LUT_AMPL_WIDTH),
		29823 => to_signed(9129, LUT_AMPL_WIDTH),
		29824 => to_signed(9126, LUT_AMPL_WIDTH),
		29825 => to_signed(9123, LUT_AMPL_WIDTH),
		29826 => to_signed(9120, LUT_AMPL_WIDTH),
		29827 => to_signed(9117, LUT_AMPL_WIDTH),
		29828 => to_signed(9114, LUT_AMPL_WIDTH),
		29829 => to_signed(9111, LUT_AMPL_WIDTH),
		29830 => to_signed(9108, LUT_AMPL_WIDTH),
		29831 => to_signed(9105, LUT_AMPL_WIDTH),
		29832 => to_signed(9102, LUT_AMPL_WIDTH),
		29833 => to_signed(9099, LUT_AMPL_WIDTH),
		29834 => to_signed(9096, LUT_AMPL_WIDTH),
		29835 => to_signed(9093, LUT_AMPL_WIDTH),
		29836 => to_signed(9090, LUT_AMPL_WIDTH),
		29837 => to_signed(9087, LUT_AMPL_WIDTH),
		29838 => to_signed(9084, LUT_AMPL_WIDTH),
		29839 => to_signed(9081, LUT_AMPL_WIDTH),
		29840 => to_signed(9078, LUT_AMPL_WIDTH),
		29841 => to_signed(9075, LUT_AMPL_WIDTH),
		29842 => to_signed(9072, LUT_AMPL_WIDTH),
		29843 => to_signed(9069, LUT_AMPL_WIDTH),
		29844 => to_signed(9066, LUT_AMPL_WIDTH),
		29845 => to_signed(9063, LUT_AMPL_WIDTH),
		29846 => to_signed(9060, LUT_AMPL_WIDTH),
		29847 => to_signed(9057, LUT_AMPL_WIDTH),
		29848 => to_signed(9054, LUT_AMPL_WIDTH),
		29849 => to_signed(9051, LUT_AMPL_WIDTH),
		29850 => to_signed(9048, LUT_AMPL_WIDTH),
		29851 => to_signed(9045, LUT_AMPL_WIDTH),
		29852 => to_signed(9042, LUT_AMPL_WIDTH),
		29853 => to_signed(9039, LUT_AMPL_WIDTH),
		29854 => to_signed(9036, LUT_AMPL_WIDTH),
		29855 => to_signed(9033, LUT_AMPL_WIDTH),
		29856 => to_signed(9030, LUT_AMPL_WIDTH),
		29857 => to_signed(9027, LUT_AMPL_WIDTH),
		29858 => to_signed(9024, LUT_AMPL_WIDTH),
		29859 => to_signed(9021, LUT_AMPL_WIDTH),
		29860 => to_signed(9018, LUT_AMPL_WIDTH),
		29861 => to_signed(9015, LUT_AMPL_WIDTH),
		29862 => to_signed(9012, LUT_AMPL_WIDTH),
		29863 => to_signed(9009, LUT_AMPL_WIDTH),
		29864 => to_signed(9006, LUT_AMPL_WIDTH),
		29865 => to_signed(9002, LUT_AMPL_WIDTH),
		29866 => to_signed(8999, LUT_AMPL_WIDTH),
		29867 => to_signed(8996, LUT_AMPL_WIDTH),
		29868 => to_signed(8993, LUT_AMPL_WIDTH),
		29869 => to_signed(8990, LUT_AMPL_WIDTH),
		29870 => to_signed(8987, LUT_AMPL_WIDTH),
		29871 => to_signed(8984, LUT_AMPL_WIDTH),
		29872 => to_signed(8981, LUT_AMPL_WIDTH),
		29873 => to_signed(8978, LUT_AMPL_WIDTH),
		29874 => to_signed(8975, LUT_AMPL_WIDTH),
		29875 => to_signed(8972, LUT_AMPL_WIDTH),
		29876 => to_signed(8969, LUT_AMPL_WIDTH),
		29877 => to_signed(8966, LUT_AMPL_WIDTH),
		29878 => to_signed(8963, LUT_AMPL_WIDTH),
		29879 => to_signed(8960, LUT_AMPL_WIDTH),
		29880 => to_signed(8957, LUT_AMPL_WIDTH),
		29881 => to_signed(8954, LUT_AMPL_WIDTH),
		29882 => to_signed(8951, LUT_AMPL_WIDTH),
		29883 => to_signed(8948, LUT_AMPL_WIDTH),
		29884 => to_signed(8945, LUT_AMPL_WIDTH),
		29885 => to_signed(8942, LUT_AMPL_WIDTH),
		29886 => to_signed(8939, LUT_AMPL_WIDTH),
		29887 => to_signed(8936, LUT_AMPL_WIDTH),
		29888 => to_signed(8933, LUT_AMPL_WIDTH),
		29889 => to_signed(8930, LUT_AMPL_WIDTH),
		29890 => to_signed(8927, LUT_AMPL_WIDTH),
		29891 => to_signed(8924, LUT_AMPL_WIDTH),
		29892 => to_signed(8921, LUT_AMPL_WIDTH),
		29893 => to_signed(8918, LUT_AMPL_WIDTH),
		29894 => to_signed(8915, LUT_AMPL_WIDTH),
		29895 => to_signed(8912, LUT_AMPL_WIDTH),
		29896 => to_signed(8909, LUT_AMPL_WIDTH),
		29897 => to_signed(8906, LUT_AMPL_WIDTH),
		29898 => to_signed(8903, LUT_AMPL_WIDTH),
		29899 => to_signed(8900, LUT_AMPL_WIDTH),
		29900 => to_signed(8897, LUT_AMPL_WIDTH),
		29901 => to_signed(8894, LUT_AMPL_WIDTH),
		29902 => to_signed(8891, LUT_AMPL_WIDTH),
		29903 => to_signed(8888, LUT_AMPL_WIDTH),
		29904 => to_signed(8885, LUT_AMPL_WIDTH),
		29905 => to_signed(8882, LUT_AMPL_WIDTH),
		29906 => to_signed(8879, LUT_AMPL_WIDTH),
		29907 => to_signed(8876, LUT_AMPL_WIDTH),
		29908 => to_signed(8873, LUT_AMPL_WIDTH),
		29909 => to_signed(8869, LUT_AMPL_WIDTH),
		29910 => to_signed(8866, LUT_AMPL_WIDTH),
		29911 => to_signed(8863, LUT_AMPL_WIDTH),
		29912 => to_signed(8860, LUT_AMPL_WIDTH),
		29913 => to_signed(8857, LUT_AMPL_WIDTH),
		29914 => to_signed(8854, LUT_AMPL_WIDTH),
		29915 => to_signed(8851, LUT_AMPL_WIDTH),
		29916 => to_signed(8848, LUT_AMPL_WIDTH),
		29917 => to_signed(8845, LUT_AMPL_WIDTH),
		29918 => to_signed(8842, LUT_AMPL_WIDTH),
		29919 => to_signed(8839, LUT_AMPL_WIDTH),
		29920 => to_signed(8836, LUT_AMPL_WIDTH),
		29921 => to_signed(8833, LUT_AMPL_WIDTH),
		29922 => to_signed(8830, LUT_AMPL_WIDTH),
		29923 => to_signed(8827, LUT_AMPL_WIDTH),
		29924 => to_signed(8824, LUT_AMPL_WIDTH),
		29925 => to_signed(8821, LUT_AMPL_WIDTH),
		29926 => to_signed(8818, LUT_AMPL_WIDTH),
		29927 => to_signed(8815, LUT_AMPL_WIDTH),
		29928 => to_signed(8812, LUT_AMPL_WIDTH),
		29929 => to_signed(8809, LUT_AMPL_WIDTH),
		29930 => to_signed(8806, LUT_AMPL_WIDTH),
		29931 => to_signed(8803, LUT_AMPL_WIDTH),
		29932 => to_signed(8800, LUT_AMPL_WIDTH),
		29933 => to_signed(8797, LUT_AMPL_WIDTH),
		29934 => to_signed(8794, LUT_AMPL_WIDTH),
		29935 => to_signed(8791, LUT_AMPL_WIDTH),
		29936 => to_signed(8788, LUT_AMPL_WIDTH),
		29937 => to_signed(8785, LUT_AMPL_WIDTH),
		29938 => to_signed(8782, LUT_AMPL_WIDTH),
		29939 => to_signed(8779, LUT_AMPL_WIDTH),
		29940 => to_signed(8776, LUT_AMPL_WIDTH),
		29941 => to_signed(8773, LUT_AMPL_WIDTH),
		29942 => to_signed(8770, LUT_AMPL_WIDTH),
		29943 => to_signed(8767, LUT_AMPL_WIDTH),
		29944 => to_signed(8764, LUT_AMPL_WIDTH),
		29945 => to_signed(8761, LUT_AMPL_WIDTH),
		29946 => to_signed(8758, LUT_AMPL_WIDTH),
		29947 => to_signed(8755, LUT_AMPL_WIDTH),
		29948 => to_signed(8751, LUT_AMPL_WIDTH),
		29949 => to_signed(8748, LUT_AMPL_WIDTH),
		29950 => to_signed(8745, LUT_AMPL_WIDTH),
		29951 => to_signed(8742, LUT_AMPL_WIDTH),
		29952 => to_signed(8739, LUT_AMPL_WIDTH),
		29953 => to_signed(8736, LUT_AMPL_WIDTH),
		29954 => to_signed(8733, LUT_AMPL_WIDTH),
		29955 => to_signed(8730, LUT_AMPL_WIDTH),
		29956 => to_signed(8727, LUT_AMPL_WIDTH),
		29957 => to_signed(8724, LUT_AMPL_WIDTH),
		29958 => to_signed(8721, LUT_AMPL_WIDTH),
		29959 => to_signed(8718, LUT_AMPL_WIDTH),
		29960 => to_signed(8715, LUT_AMPL_WIDTH),
		29961 => to_signed(8712, LUT_AMPL_WIDTH),
		29962 => to_signed(8709, LUT_AMPL_WIDTH),
		29963 => to_signed(8706, LUT_AMPL_WIDTH),
		29964 => to_signed(8703, LUT_AMPL_WIDTH),
		29965 => to_signed(8700, LUT_AMPL_WIDTH),
		29966 => to_signed(8697, LUT_AMPL_WIDTH),
		29967 => to_signed(8694, LUT_AMPL_WIDTH),
		29968 => to_signed(8691, LUT_AMPL_WIDTH),
		29969 => to_signed(8688, LUT_AMPL_WIDTH),
		29970 => to_signed(8685, LUT_AMPL_WIDTH),
		29971 => to_signed(8682, LUT_AMPL_WIDTH),
		29972 => to_signed(8679, LUT_AMPL_WIDTH),
		29973 => to_signed(8676, LUT_AMPL_WIDTH),
		29974 => to_signed(8673, LUT_AMPL_WIDTH),
		29975 => to_signed(8670, LUT_AMPL_WIDTH),
		29976 => to_signed(8667, LUT_AMPL_WIDTH),
		29977 => to_signed(8664, LUT_AMPL_WIDTH),
		29978 => to_signed(8661, LUT_AMPL_WIDTH),
		29979 => to_signed(8658, LUT_AMPL_WIDTH),
		29980 => to_signed(8655, LUT_AMPL_WIDTH),
		29981 => to_signed(8652, LUT_AMPL_WIDTH),
		29982 => to_signed(8649, LUT_AMPL_WIDTH),
		29983 => to_signed(8645, LUT_AMPL_WIDTH),
		29984 => to_signed(8642, LUT_AMPL_WIDTH),
		29985 => to_signed(8639, LUT_AMPL_WIDTH),
		29986 => to_signed(8636, LUT_AMPL_WIDTH),
		29987 => to_signed(8633, LUT_AMPL_WIDTH),
		29988 => to_signed(8630, LUT_AMPL_WIDTH),
		29989 => to_signed(8627, LUT_AMPL_WIDTH),
		29990 => to_signed(8624, LUT_AMPL_WIDTH),
		29991 => to_signed(8621, LUT_AMPL_WIDTH),
		29992 => to_signed(8618, LUT_AMPL_WIDTH),
		29993 => to_signed(8615, LUT_AMPL_WIDTH),
		29994 => to_signed(8612, LUT_AMPL_WIDTH),
		29995 => to_signed(8609, LUT_AMPL_WIDTH),
		29996 => to_signed(8606, LUT_AMPL_WIDTH),
		29997 => to_signed(8603, LUT_AMPL_WIDTH),
		29998 => to_signed(8600, LUT_AMPL_WIDTH),
		29999 => to_signed(8597, LUT_AMPL_WIDTH),
		30000 => to_signed(8594, LUT_AMPL_WIDTH),
		30001 => to_signed(8591, LUT_AMPL_WIDTH),
		30002 => to_signed(8588, LUT_AMPL_WIDTH),
		30003 => to_signed(8585, LUT_AMPL_WIDTH),
		30004 => to_signed(8582, LUT_AMPL_WIDTH),
		30005 => to_signed(8579, LUT_AMPL_WIDTH),
		30006 => to_signed(8576, LUT_AMPL_WIDTH),
		30007 => to_signed(8573, LUT_AMPL_WIDTH),
		30008 => to_signed(8570, LUT_AMPL_WIDTH),
		30009 => to_signed(8567, LUT_AMPL_WIDTH),
		30010 => to_signed(8564, LUT_AMPL_WIDTH),
		30011 => to_signed(8561, LUT_AMPL_WIDTH),
		30012 => to_signed(8558, LUT_AMPL_WIDTH),
		30013 => to_signed(8555, LUT_AMPL_WIDTH),
		30014 => to_signed(8552, LUT_AMPL_WIDTH),
		30015 => to_signed(8548, LUT_AMPL_WIDTH),
		30016 => to_signed(8545, LUT_AMPL_WIDTH),
		30017 => to_signed(8542, LUT_AMPL_WIDTH),
		30018 => to_signed(8539, LUT_AMPL_WIDTH),
		30019 => to_signed(8536, LUT_AMPL_WIDTH),
		30020 => to_signed(8533, LUT_AMPL_WIDTH),
		30021 => to_signed(8530, LUT_AMPL_WIDTH),
		30022 => to_signed(8527, LUT_AMPL_WIDTH),
		30023 => to_signed(8524, LUT_AMPL_WIDTH),
		30024 => to_signed(8521, LUT_AMPL_WIDTH),
		30025 => to_signed(8518, LUT_AMPL_WIDTH),
		30026 => to_signed(8515, LUT_AMPL_WIDTH),
		30027 => to_signed(8512, LUT_AMPL_WIDTH),
		30028 => to_signed(8509, LUT_AMPL_WIDTH),
		30029 => to_signed(8506, LUT_AMPL_WIDTH),
		30030 => to_signed(8503, LUT_AMPL_WIDTH),
		30031 => to_signed(8500, LUT_AMPL_WIDTH),
		30032 => to_signed(8497, LUT_AMPL_WIDTH),
		30033 => to_signed(8494, LUT_AMPL_WIDTH),
		30034 => to_signed(8491, LUT_AMPL_WIDTH),
		30035 => to_signed(8488, LUT_AMPL_WIDTH),
		30036 => to_signed(8485, LUT_AMPL_WIDTH),
		30037 => to_signed(8482, LUT_AMPL_WIDTH),
		30038 => to_signed(8479, LUT_AMPL_WIDTH),
		30039 => to_signed(8476, LUT_AMPL_WIDTH),
		30040 => to_signed(8473, LUT_AMPL_WIDTH),
		30041 => to_signed(8470, LUT_AMPL_WIDTH),
		30042 => to_signed(8467, LUT_AMPL_WIDTH),
		30043 => to_signed(8464, LUT_AMPL_WIDTH),
		30044 => to_signed(8460, LUT_AMPL_WIDTH),
		30045 => to_signed(8457, LUT_AMPL_WIDTH),
		30046 => to_signed(8454, LUT_AMPL_WIDTH),
		30047 => to_signed(8451, LUT_AMPL_WIDTH),
		30048 => to_signed(8448, LUT_AMPL_WIDTH),
		30049 => to_signed(8445, LUT_AMPL_WIDTH),
		30050 => to_signed(8442, LUT_AMPL_WIDTH),
		30051 => to_signed(8439, LUT_AMPL_WIDTH),
		30052 => to_signed(8436, LUT_AMPL_WIDTH),
		30053 => to_signed(8433, LUT_AMPL_WIDTH),
		30054 => to_signed(8430, LUT_AMPL_WIDTH),
		30055 => to_signed(8427, LUT_AMPL_WIDTH),
		30056 => to_signed(8424, LUT_AMPL_WIDTH),
		30057 => to_signed(8421, LUT_AMPL_WIDTH),
		30058 => to_signed(8418, LUT_AMPL_WIDTH),
		30059 => to_signed(8415, LUT_AMPL_WIDTH),
		30060 => to_signed(8412, LUT_AMPL_WIDTH),
		30061 => to_signed(8409, LUT_AMPL_WIDTH),
		30062 => to_signed(8406, LUT_AMPL_WIDTH),
		30063 => to_signed(8403, LUT_AMPL_WIDTH),
		30064 => to_signed(8400, LUT_AMPL_WIDTH),
		30065 => to_signed(8397, LUT_AMPL_WIDTH),
		30066 => to_signed(8394, LUT_AMPL_WIDTH),
		30067 => to_signed(8391, LUT_AMPL_WIDTH),
		30068 => to_signed(8388, LUT_AMPL_WIDTH),
		30069 => to_signed(8385, LUT_AMPL_WIDTH),
		30070 => to_signed(8382, LUT_AMPL_WIDTH),
		30071 => to_signed(8379, LUT_AMPL_WIDTH),
		30072 => to_signed(8375, LUT_AMPL_WIDTH),
		30073 => to_signed(8372, LUT_AMPL_WIDTH),
		30074 => to_signed(8369, LUT_AMPL_WIDTH),
		30075 => to_signed(8366, LUT_AMPL_WIDTH),
		30076 => to_signed(8363, LUT_AMPL_WIDTH),
		30077 => to_signed(8360, LUT_AMPL_WIDTH),
		30078 => to_signed(8357, LUT_AMPL_WIDTH),
		30079 => to_signed(8354, LUT_AMPL_WIDTH),
		30080 => to_signed(8351, LUT_AMPL_WIDTH),
		30081 => to_signed(8348, LUT_AMPL_WIDTH),
		30082 => to_signed(8345, LUT_AMPL_WIDTH),
		30083 => to_signed(8342, LUT_AMPL_WIDTH),
		30084 => to_signed(8339, LUT_AMPL_WIDTH),
		30085 => to_signed(8336, LUT_AMPL_WIDTH),
		30086 => to_signed(8333, LUT_AMPL_WIDTH),
		30087 => to_signed(8330, LUT_AMPL_WIDTH),
		30088 => to_signed(8327, LUT_AMPL_WIDTH),
		30089 => to_signed(8324, LUT_AMPL_WIDTH),
		30090 => to_signed(8321, LUT_AMPL_WIDTH),
		30091 => to_signed(8318, LUT_AMPL_WIDTH),
		30092 => to_signed(8315, LUT_AMPL_WIDTH),
		30093 => to_signed(8312, LUT_AMPL_WIDTH),
		30094 => to_signed(8309, LUT_AMPL_WIDTH),
		30095 => to_signed(8306, LUT_AMPL_WIDTH),
		30096 => to_signed(8303, LUT_AMPL_WIDTH),
		30097 => to_signed(8300, LUT_AMPL_WIDTH),
		30098 => to_signed(8296, LUT_AMPL_WIDTH),
		30099 => to_signed(8293, LUT_AMPL_WIDTH),
		30100 => to_signed(8290, LUT_AMPL_WIDTH),
		30101 => to_signed(8287, LUT_AMPL_WIDTH),
		30102 => to_signed(8284, LUT_AMPL_WIDTH),
		30103 => to_signed(8281, LUT_AMPL_WIDTH),
		30104 => to_signed(8278, LUT_AMPL_WIDTH),
		30105 => to_signed(8275, LUT_AMPL_WIDTH),
		30106 => to_signed(8272, LUT_AMPL_WIDTH),
		30107 => to_signed(8269, LUT_AMPL_WIDTH),
		30108 => to_signed(8266, LUT_AMPL_WIDTH),
		30109 => to_signed(8263, LUT_AMPL_WIDTH),
		30110 => to_signed(8260, LUT_AMPL_WIDTH),
		30111 => to_signed(8257, LUT_AMPL_WIDTH),
		30112 => to_signed(8254, LUT_AMPL_WIDTH),
		30113 => to_signed(8251, LUT_AMPL_WIDTH),
		30114 => to_signed(8248, LUT_AMPL_WIDTH),
		30115 => to_signed(8245, LUT_AMPL_WIDTH),
		30116 => to_signed(8242, LUT_AMPL_WIDTH),
		30117 => to_signed(8239, LUT_AMPL_WIDTH),
		30118 => to_signed(8236, LUT_AMPL_WIDTH),
		30119 => to_signed(8233, LUT_AMPL_WIDTH),
		30120 => to_signed(8230, LUT_AMPL_WIDTH),
		30121 => to_signed(8227, LUT_AMPL_WIDTH),
		30122 => to_signed(8224, LUT_AMPL_WIDTH),
		30123 => to_signed(8220, LUT_AMPL_WIDTH),
		30124 => to_signed(8217, LUT_AMPL_WIDTH),
		30125 => to_signed(8214, LUT_AMPL_WIDTH),
		30126 => to_signed(8211, LUT_AMPL_WIDTH),
		30127 => to_signed(8208, LUT_AMPL_WIDTH),
		30128 => to_signed(8205, LUT_AMPL_WIDTH),
		30129 => to_signed(8202, LUT_AMPL_WIDTH),
		30130 => to_signed(8199, LUT_AMPL_WIDTH),
		30131 => to_signed(8196, LUT_AMPL_WIDTH),
		30132 => to_signed(8193, LUT_AMPL_WIDTH),
		30133 => to_signed(8190, LUT_AMPL_WIDTH),
		30134 => to_signed(8187, LUT_AMPL_WIDTH),
		30135 => to_signed(8184, LUT_AMPL_WIDTH),
		30136 => to_signed(8181, LUT_AMPL_WIDTH),
		30137 => to_signed(8178, LUT_AMPL_WIDTH),
		30138 => to_signed(8175, LUT_AMPL_WIDTH),
		30139 => to_signed(8172, LUT_AMPL_WIDTH),
		30140 => to_signed(8169, LUT_AMPL_WIDTH),
		30141 => to_signed(8166, LUT_AMPL_WIDTH),
		30142 => to_signed(8163, LUT_AMPL_WIDTH),
		30143 => to_signed(8160, LUT_AMPL_WIDTH),
		30144 => to_signed(8157, LUT_AMPL_WIDTH),
		30145 => to_signed(8154, LUT_AMPL_WIDTH),
		30146 => to_signed(8151, LUT_AMPL_WIDTH),
		30147 => to_signed(8147, LUT_AMPL_WIDTH),
		30148 => to_signed(8144, LUT_AMPL_WIDTH),
		30149 => to_signed(8141, LUT_AMPL_WIDTH),
		30150 => to_signed(8138, LUT_AMPL_WIDTH),
		30151 => to_signed(8135, LUT_AMPL_WIDTH),
		30152 => to_signed(8132, LUT_AMPL_WIDTH),
		30153 => to_signed(8129, LUT_AMPL_WIDTH),
		30154 => to_signed(8126, LUT_AMPL_WIDTH),
		30155 => to_signed(8123, LUT_AMPL_WIDTH),
		30156 => to_signed(8120, LUT_AMPL_WIDTH),
		30157 => to_signed(8117, LUT_AMPL_WIDTH),
		30158 => to_signed(8114, LUT_AMPL_WIDTH),
		30159 => to_signed(8111, LUT_AMPL_WIDTH),
		30160 => to_signed(8108, LUT_AMPL_WIDTH),
		30161 => to_signed(8105, LUT_AMPL_WIDTH),
		30162 => to_signed(8102, LUT_AMPL_WIDTH),
		30163 => to_signed(8099, LUT_AMPL_WIDTH),
		30164 => to_signed(8096, LUT_AMPL_WIDTH),
		30165 => to_signed(8093, LUT_AMPL_WIDTH),
		30166 => to_signed(8090, LUT_AMPL_WIDTH),
		30167 => to_signed(8087, LUT_AMPL_WIDTH),
		30168 => to_signed(8084, LUT_AMPL_WIDTH),
		30169 => to_signed(8081, LUT_AMPL_WIDTH),
		30170 => to_signed(8077, LUT_AMPL_WIDTH),
		30171 => to_signed(8074, LUT_AMPL_WIDTH),
		30172 => to_signed(8071, LUT_AMPL_WIDTH),
		30173 => to_signed(8068, LUT_AMPL_WIDTH),
		30174 => to_signed(8065, LUT_AMPL_WIDTH),
		30175 => to_signed(8062, LUT_AMPL_WIDTH),
		30176 => to_signed(8059, LUT_AMPL_WIDTH),
		30177 => to_signed(8056, LUT_AMPL_WIDTH),
		30178 => to_signed(8053, LUT_AMPL_WIDTH),
		30179 => to_signed(8050, LUT_AMPL_WIDTH),
		30180 => to_signed(8047, LUT_AMPL_WIDTH),
		30181 => to_signed(8044, LUT_AMPL_WIDTH),
		30182 => to_signed(8041, LUT_AMPL_WIDTH),
		30183 => to_signed(8038, LUT_AMPL_WIDTH),
		30184 => to_signed(8035, LUT_AMPL_WIDTH),
		30185 => to_signed(8032, LUT_AMPL_WIDTH),
		30186 => to_signed(8029, LUT_AMPL_WIDTH),
		30187 => to_signed(8026, LUT_AMPL_WIDTH),
		30188 => to_signed(8023, LUT_AMPL_WIDTH),
		30189 => to_signed(8020, LUT_AMPL_WIDTH),
		30190 => to_signed(8017, LUT_AMPL_WIDTH),
		30191 => to_signed(8014, LUT_AMPL_WIDTH),
		30192 => to_signed(8010, LUT_AMPL_WIDTH),
		30193 => to_signed(8007, LUT_AMPL_WIDTH),
		30194 => to_signed(8004, LUT_AMPL_WIDTH),
		30195 => to_signed(8001, LUT_AMPL_WIDTH),
		30196 => to_signed(7998, LUT_AMPL_WIDTH),
		30197 => to_signed(7995, LUT_AMPL_WIDTH),
		30198 => to_signed(7992, LUT_AMPL_WIDTH),
		30199 => to_signed(7989, LUT_AMPL_WIDTH),
		30200 => to_signed(7986, LUT_AMPL_WIDTH),
		30201 => to_signed(7983, LUT_AMPL_WIDTH),
		30202 => to_signed(7980, LUT_AMPL_WIDTH),
		30203 => to_signed(7977, LUT_AMPL_WIDTH),
		30204 => to_signed(7974, LUT_AMPL_WIDTH),
		30205 => to_signed(7971, LUT_AMPL_WIDTH),
		30206 => to_signed(7968, LUT_AMPL_WIDTH),
		30207 => to_signed(7965, LUT_AMPL_WIDTH),
		30208 => to_signed(7962, LUT_AMPL_WIDTH),
		30209 => to_signed(7959, LUT_AMPL_WIDTH),
		30210 => to_signed(7956, LUT_AMPL_WIDTH),
		30211 => to_signed(7953, LUT_AMPL_WIDTH),
		30212 => to_signed(7950, LUT_AMPL_WIDTH),
		30213 => to_signed(7946, LUT_AMPL_WIDTH),
		30214 => to_signed(7943, LUT_AMPL_WIDTH),
		30215 => to_signed(7940, LUT_AMPL_WIDTH),
		30216 => to_signed(7937, LUT_AMPL_WIDTH),
		30217 => to_signed(7934, LUT_AMPL_WIDTH),
		30218 => to_signed(7931, LUT_AMPL_WIDTH),
		30219 => to_signed(7928, LUT_AMPL_WIDTH),
		30220 => to_signed(7925, LUT_AMPL_WIDTH),
		30221 => to_signed(7922, LUT_AMPL_WIDTH),
		30222 => to_signed(7919, LUT_AMPL_WIDTH),
		30223 => to_signed(7916, LUT_AMPL_WIDTH),
		30224 => to_signed(7913, LUT_AMPL_WIDTH),
		30225 => to_signed(7910, LUT_AMPL_WIDTH),
		30226 => to_signed(7907, LUT_AMPL_WIDTH),
		30227 => to_signed(7904, LUT_AMPL_WIDTH),
		30228 => to_signed(7901, LUT_AMPL_WIDTH),
		30229 => to_signed(7898, LUT_AMPL_WIDTH),
		30230 => to_signed(7895, LUT_AMPL_WIDTH),
		30231 => to_signed(7892, LUT_AMPL_WIDTH),
		30232 => to_signed(7889, LUT_AMPL_WIDTH),
		30233 => to_signed(7886, LUT_AMPL_WIDTH),
		30234 => to_signed(7882, LUT_AMPL_WIDTH),
		30235 => to_signed(7879, LUT_AMPL_WIDTH),
		30236 => to_signed(7876, LUT_AMPL_WIDTH),
		30237 => to_signed(7873, LUT_AMPL_WIDTH),
		30238 => to_signed(7870, LUT_AMPL_WIDTH),
		30239 => to_signed(7867, LUT_AMPL_WIDTH),
		30240 => to_signed(7864, LUT_AMPL_WIDTH),
		30241 => to_signed(7861, LUT_AMPL_WIDTH),
		30242 => to_signed(7858, LUT_AMPL_WIDTH),
		30243 => to_signed(7855, LUT_AMPL_WIDTH),
		30244 => to_signed(7852, LUT_AMPL_WIDTH),
		30245 => to_signed(7849, LUT_AMPL_WIDTH),
		30246 => to_signed(7846, LUT_AMPL_WIDTH),
		30247 => to_signed(7843, LUT_AMPL_WIDTH),
		30248 => to_signed(7840, LUT_AMPL_WIDTH),
		30249 => to_signed(7837, LUT_AMPL_WIDTH),
		30250 => to_signed(7834, LUT_AMPL_WIDTH),
		30251 => to_signed(7831, LUT_AMPL_WIDTH),
		30252 => to_signed(7828, LUT_AMPL_WIDTH),
		30253 => to_signed(7825, LUT_AMPL_WIDTH),
		30254 => to_signed(7821, LUT_AMPL_WIDTH),
		30255 => to_signed(7818, LUT_AMPL_WIDTH),
		30256 => to_signed(7815, LUT_AMPL_WIDTH),
		30257 => to_signed(7812, LUT_AMPL_WIDTH),
		30258 => to_signed(7809, LUT_AMPL_WIDTH),
		30259 => to_signed(7806, LUT_AMPL_WIDTH),
		30260 => to_signed(7803, LUT_AMPL_WIDTH),
		30261 => to_signed(7800, LUT_AMPL_WIDTH),
		30262 => to_signed(7797, LUT_AMPL_WIDTH),
		30263 => to_signed(7794, LUT_AMPL_WIDTH),
		30264 => to_signed(7791, LUT_AMPL_WIDTH),
		30265 => to_signed(7788, LUT_AMPL_WIDTH),
		30266 => to_signed(7785, LUT_AMPL_WIDTH),
		30267 => to_signed(7782, LUT_AMPL_WIDTH),
		30268 => to_signed(7779, LUT_AMPL_WIDTH),
		30269 => to_signed(7776, LUT_AMPL_WIDTH),
		30270 => to_signed(7773, LUT_AMPL_WIDTH),
		30271 => to_signed(7770, LUT_AMPL_WIDTH),
		30272 => to_signed(7767, LUT_AMPL_WIDTH),
		30273 => to_signed(7764, LUT_AMPL_WIDTH),
		30274 => to_signed(7760, LUT_AMPL_WIDTH),
		30275 => to_signed(7757, LUT_AMPL_WIDTH),
		30276 => to_signed(7754, LUT_AMPL_WIDTH),
		30277 => to_signed(7751, LUT_AMPL_WIDTH),
		30278 => to_signed(7748, LUT_AMPL_WIDTH),
		30279 => to_signed(7745, LUT_AMPL_WIDTH),
		30280 => to_signed(7742, LUT_AMPL_WIDTH),
		30281 => to_signed(7739, LUT_AMPL_WIDTH),
		30282 => to_signed(7736, LUT_AMPL_WIDTH),
		30283 => to_signed(7733, LUT_AMPL_WIDTH),
		30284 => to_signed(7730, LUT_AMPL_WIDTH),
		30285 => to_signed(7727, LUT_AMPL_WIDTH),
		30286 => to_signed(7724, LUT_AMPL_WIDTH),
		30287 => to_signed(7721, LUT_AMPL_WIDTH),
		30288 => to_signed(7718, LUT_AMPL_WIDTH),
		30289 => to_signed(7715, LUT_AMPL_WIDTH),
		30290 => to_signed(7712, LUT_AMPL_WIDTH),
		30291 => to_signed(7709, LUT_AMPL_WIDTH),
		30292 => to_signed(7705, LUT_AMPL_WIDTH),
		30293 => to_signed(7702, LUT_AMPL_WIDTH),
		30294 => to_signed(7699, LUT_AMPL_WIDTH),
		30295 => to_signed(7696, LUT_AMPL_WIDTH),
		30296 => to_signed(7693, LUT_AMPL_WIDTH),
		30297 => to_signed(7690, LUT_AMPL_WIDTH),
		30298 => to_signed(7687, LUT_AMPL_WIDTH),
		30299 => to_signed(7684, LUT_AMPL_WIDTH),
		30300 => to_signed(7681, LUT_AMPL_WIDTH),
		30301 => to_signed(7678, LUT_AMPL_WIDTH),
		30302 => to_signed(7675, LUT_AMPL_WIDTH),
		30303 => to_signed(7672, LUT_AMPL_WIDTH),
		30304 => to_signed(7669, LUT_AMPL_WIDTH),
		30305 => to_signed(7666, LUT_AMPL_WIDTH),
		30306 => to_signed(7663, LUT_AMPL_WIDTH),
		30307 => to_signed(7660, LUT_AMPL_WIDTH),
		30308 => to_signed(7657, LUT_AMPL_WIDTH),
		30309 => to_signed(7654, LUT_AMPL_WIDTH),
		30310 => to_signed(7651, LUT_AMPL_WIDTH),
		30311 => to_signed(7647, LUT_AMPL_WIDTH),
		30312 => to_signed(7644, LUT_AMPL_WIDTH),
		30313 => to_signed(7641, LUT_AMPL_WIDTH),
		30314 => to_signed(7638, LUT_AMPL_WIDTH),
		30315 => to_signed(7635, LUT_AMPL_WIDTH),
		30316 => to_signed(7632, LUT_AMPL_WIDTH),
		30317 => to_signed(7629, LUT_AMPL_WIDTH),
		30318 => to_signed(7626, LUT_AMPL_WIDTH),
		30319 => to_signed(7623, LUT_AMPL_WIDTH),
		30320 => to_signed(7620, LUT_AMPL_WIDTH),
		30321 => to_signed(7617, LUT_AMPL_WIDTH),
		30322 => to_signed(7614, LUT_AMPL_WIDTH),
		30323 => to_signed(7611, LUT_AMPL_WIDTH),
		30324 => to_signed(7608, LUT_AMPL_WIDTH),
		30325 => to_signed(7605, LUT_AMPL_WIDTH),
		30326 => to_signed(7602, LUT_AMPL_WIDTH),
		30327 => to_signed(7599, LUT_AMPL_WIDTH),
		30328 => to_signed(7596, LUT_AMPL_WIDTH),
		30329 => to_signed(7592, LUT_AMPL_WIDTH),
		30330 => to_signed(7589, LUT_AMPL_WIDTH),
		30331 => to_signed(7586, LUT_AMPL_WIDTH),
		30332 => to_signed(7583, LUT_AMPL_WIDTH),
		30333 => to_signed(7580, LUT_AMPL_WIDTH),
		30334 => to_signed(7577, LUT_AMPL_WIDTH),
		30335 => to_signed(7574, LUT_AMPL_WIDTH),
		30336 => to_signed(7571, LUT_AMPL_WIDTH),
		30337 => to_signed(7568, LUT_AMPL_WIDTH),
		30338 => to_signed(7565, LUT_AMPL_WIDTH),
		30339 => to_signed(7562, LUT_AMPL_WIDTH),
		30340 => to_signed(7559, LUT_AMPL_WIDTH),
		30341 => to_signed(7556, LUT_AMPL_WIDTH),
		30342 => to_signed(7553, LUT_AMPL_WIDTH),
		30343 => to_signed(7550, LUT_AMPL_WIDTH),
		30344 => to_signed(7547, LUT_AMPL_WIDTH),
		30345 => to_signed(7544, LUT_AMPL_WIDTH),
		30346 => to_signed(7541, LUT_AMPL_WIDTH),
		30347 => to_signed(7537, LUT_AMPL_WIDTH),
		30348 => to_signed(7534, LUT_AMPL_WIDTH),
		30349 => to_signed(7531, LUT_AMPL_WIDTH),
		30350 => to_signed(7528, LUT_AMPL_WIDTH),
		30351 => to_signed(7525, LUT_AMPL_WIDTH),
		30352 => to_signed(7522, LUT_AMPL_WIDTH),
		30353 => to_signed(7519, LUT_AMPL_WIDTH),
		30354 => to_signed(7516, LUT_AMPL_WIDTH),
		30355 => to_signed(7513, LUT_AMPL_WIDTH),
		30356 => to_signed(7510, LUT_AMPL_WIDTH),
		30357 => to_signed(7507, LUT_AMPL_WIDTH),
		30358 => to_signed(7504, LUT_AMPL_WIDTH),
		30359 => to_signed(7501, LUT_AMPL_WIDTH),
		30360 => to_signed(7498, LUT_AMPL_WIDTH),
		30361 => to_signed(7495, LUT_AMPL_WIDTH),
		30362 => to_signed(7492, LUT_AMPL_WIDTH),
		30363 => to_signed(7489, LUT_AMPL_WIDTH),
		30364 => to_signed(7485, LUT_AMPL_WIDTH),
		30365 => to_signed(7482, LUT_AMPL_WIDTH),
		30366 => to_signed(7479, LUT_AMPL_WIDTH),
		30367 => to_signed(7476, LUT_AMPL_WIDTH),
		30368 => to_signed(7473, LUT_AMPL_WIDTH),
		30369 => to_signed(7470, LUT_AMPL_WIDTH),
		30370 => to_signed(7467, LUT_AMPL_WIDTH),
		30371 => to_signed(7464, LUT_AMPL_WIDTH),
		30372 => to_signed(7461, LUT_AMPL_WIDTH),
		30373 => to_signed(7458, LUT_AMPL_WIDTH),
		30374 => to_signed(7455, LUT_AMPL_WIDTH),
		30375 => to_signed(7452, LUT_AMPL_WIDTH),
		30376 => to_signed(7449, LUT_AMPL_WIDTH),
		30377 => to_signed(7446, LUT_AMPL_WIDTH),
		30378 => to_signed(7443, LUT_AMPL_WIDTH),
		30379 => to_signed(7440, LUT_AMPL_WIDTH),
		30380 => to_signed(7437, LUT_AMPL_WIDTH),
		30381 => to_signed(7433, LUT_AMPL_WIDTH),
		30382 => to_signed(7430, LUT_AMPL_WIDTH),
		30383 => to_signed(7427, LUT_AMPL_WIDTH),
		30384 => to_signed(7424, LUT_AMPL_WIDTH),
		30385 => to_signed(7421, LUT_AMPL_WIDTH),
		30386 => to_signed(7418, LUT_AMPL_WIDTH),
		30387 => to_signed(7415, LUT_AMPL_WIDTH),
		30388 => to_signed(7412, LUT_AMPL_WIDTH),
		30389 => to_signed(7409, LUT_AMPL_WIDTH),
		30390 => to_signed(7406, LUT_AMPL_WIDTH),
		30391 => to_signed(7403, LUT_AMPL_WIDTH),
		30392 => to_signed(7400, LUT_AMPL_WIDTH),
		30393 => to_signed(7397, LUT_AMPL_WIDTH),
		30394 => to_signed(7394, LUT_AMPL_WIDTH),
		30395 => to_signed(7391, LUT_AMPL_WIDTH),
		30396 => to_signed(7388, LUT_AMPL_WIDTH),
		30397 => to_signed(7385, LUT_AMPL_WIDTH),
		30398 => to_signed(7381, LUT_AMPL_WIDTH),
		30399 => to_signed(7378, LUT_AMPL_WIDTH),
		30400 => to_signed(7375, LUT_AMPL_WIDTH),
		30401 => to_signed(7372, LUT_AMPL_WIDTH),
		30402 => to_signed(7369, LUT_AMPL_WIDTH),
		30403 => to_signed(7366, LUT_AMPL_WIDTH),
		30404 => to_signed(7363, LUT_AMPL_WIDTH),
		30405 => to_signed(7360, LUT_AMPL_WIDTH),
		30406 => to_signed(7357, LUT_AMPL_WIDTH),
		30407 => to_signed(7354, LUT_AMPL_WIDTH),
		30408 => to_signed(7351, LUT_AMPL_WIDTH),
		30409 => to_signed(7348, LUT_AMPL_WIDTH),
		30410 => to_signed(7345, LUT_AMPL_WIDTH),
		30411 => to_signed(7342, LUT_AMPL_WIDTH),
		30412 => to_signed(7339, LUT_AMPL_WIDTH),
		30413 => to_signed(7336, LUT_AMPL_WIDTH),
		30414 => to_signed(7332, LUT_AMPL_WIDTH),
		30415 => to_signed(7329, LUT_AMPL_WIDTH),
		30416 => to_signed(7326, LUT_AMPL_WIDTH),
		30417 => to_signed(7323, LUT_AMPL_WIDTH),
		30418 => to_signed(7320, LUT_AMPL_WIDTH),
		30419 => to_signed(7317, LUT_AMPL_WIDTH),
		30420 => to_signed(7314, LUT_AMPL_WIDTH),
		30421 => to_signed(7311, LUT_AMPL_WIDTH),
		30422 => to_signed(7308, LUT_AMPL_WIDTH),
		30423 => to_signed(7305, LUT_AMPL_WIDTH),
		30424 => to_signed(7302, LUT_AMPL_WIDTH),
		30425 => to_signed(7299, LUT_AMPL_WIDTH),
		30426 => to_signed(7296, LUT_AMPL_WIDTH),
		30427 => to_signed(7293, LUT_AMPL_WIDTH),
		30428 => to_signed(7290, LUT_AMPL_WIDTH),
		30429 => to_signed(7287, LUT_AMPL_WIDTH),
		30430 => to_signed(7283, LUT_AMPL_WIDTH),
		30431 => to_signed(7280, LUT_AMPL_WIDTH),
		30432 => to_signed(7277, LUT_AMPL_WIDTH),
		30433 => to_signed(7274, LUT_AMPL_WIDTH),
		30434 => to_signed(7271, LUT_AMPL_WIDTH),
		30435 => to_signed(7268, LUT_AMPL_WIDTH),
		30436 => to_signed(7265, LUT_AMPL_WIDTH),
		30437 => to_signed(7262, LUT_AMPL_WIDTH),
		30438 => to_signed(7259, LUT_AMPL_WIDTH),
		30439 => to_signed(7256, LUT_AMPL_WIDTH),
		30440 => to_signed(7253, LUT_AMPL_WIDTH),
		30441 => to_signed(7250, LUT_AMPL_WIDTH),
		30442 => to_signed(7247, LUT_AMPL_WIDTH),
		30443 => to_signed(7244, LUT_AMPL_WIDTH),
		30444 => to_signed(7241, LUT_AMPL_WIDTH),
		30445 => to_signed(7238, LUT_AMPL_WIDTH),
		30446 => to_signed(7234, LUT_AMPL_WIDTH),
		30447 => to_signed(7231, LUT_AMPL_WIDTH),
		30448 => to_signed(7228, LUT_AMPL_WIDTH),
		30449 => to_signed(7225, LUT_AMPL_WIDTH),
		30450 => to_signed(7222, LUT_AMPL_WIDTH),
		30451 => to_signed(7219, LUT_AMPL_WIDTH),
		30452 => to_signed(7216, LUT_AMPL_WIDTH),
		30453 => to_signed(7213, LUT_AMPL_WIDTH),
		30454 => to_signed(7210, LUT_AMPL_WIDTH),
		30455 => to_signed(7207, LUT_AMPL_WIDTH),
		30456 => to_signed(7204, LUT_AMPL_WIDTH),
		30457 => to_signed(7201, LUT_AMPL_WIDTH),
		30458 => to_signed(7198, LUT_AMPL_WIDTH),
		30459 => to_signed(7195, LUT_AMPL_WIDTH),
		30460 => to_signed(7192, LUT_AMPL_WIDTH),
		30461 => to_signed(7188, LUT_AMPL_WIDTH),
		30462 => to_signed(7185, LUT_AMPL_WIDTH),
		30463 => to_signed(7182, LUT_AMPL_WIDTH),
		30464 => to_signed(7179, LUT_AMPL_WIDTH),
		30465 => to_signed(7176, LUT_AMPL_WIDTH),
		30466 => to_signed(7173, LUT_AMPL_WIDTH),
		30467 => to_signed(7170, LUT_AMPL_WIDTH),
		30468 => to_signed(7167, LUT_AMPL_WIDTH),
		30469 => to_signed(7164, LUT_AMPL_WIDTH),
		30470 => to_signed(7161, LUT_AMPL_WIDTH),
		30471 => to_signed(7158, LUT_AMPL_WIDTH),
		30472 => to_signed(7155, LUT_AMPL_WIDTH),
		30473 => to_signed(7152, LUT_AMPL_WIDTH),
		30474 => to_signed(7149, LUT_AMPL_WIDTH),
		30475 => to_signed(7146, LUT_AMPL_WIDTH),
		30476 => to_signed(7143, LUT_AMPL_WIDTH),
		30477 => to_signed(7139, LUT_AMPL_WIDTH),
		30478 => to_signed(7136, LUT_AMPL_WIDTH),
		30479 => to_signed(7133, LUT_AMPL_WIDTH),
		30480 => to_signed(7130, LUT_AMPL_WIDTH),
		30481 => to_signed(7127, LUT_AMPL_WIDTH),
		30482 => to_signed(7124, LUT_AMPL_WIDTH),
		30483 => to_signed(7121, LUT_AMPL_WIDTH),
		30484 => to_signed(7118, LUT_AMPL_WIDTH),
		30485 => to_signed(7115, LUT_AMPL_WIDTH),
		30486 => to_signed(7112, LUT_AMPL_WIDTH),
		30487 => to_signed(7109, LUT_AMPL_WIDTH),
		30488 => to_signed(7106, LUT_AMPL_WIDTH),
		30489 => to_signed(7103, LUT_AMPL_WIDTH),
		30490 => to_signed(7100, LUT_AMPL_WIDTH),
		30491 => to_signed(7097, LUT_AMPL_WIDTH),
		30492 => to_signed(7093, LUT_AMPL_WIDTH),
		30493 => to_signed(7090, LUT_AMPL_WIDTH),
		30494 => to_signed(7087, LUT_AMPL_WIDTH),
		30495 => to_signed(7084, LUT_AMPL_WIDTH),
		30496 => to_signed(7081, LUT_AMPL_WIDTH),
		30497 => to_signed(7078, LUT_AMPL_WIDTH),
		30498 => to_signed(7075, LUT_AMPL_WIDTH),
		30499 => to_signed(7072, LUT_AMPL_WIDTH),
		30500 => to_signed(7069, LUT_AMPL_WIDTH),
		30501 => to_signed(7066, LUT_AMPL_WIDTH),
		30502 => to_signed(7063, LUT_AMPL_WIDTH),
		30503 => to_signed(7060, LUT_AMPL_WIDTH),
		30504 => to_signed(7057, LUT_AMPL_WIDTH),
		30505 => to_signed(7054, LUT_AMPL_WIDTH),
		30506 => to_signed(7050, LUT_AMPL_WIDTH),
		30507 => to_signed(7047, LUT_AMPL_WIDTH),
		30508 => to_signed(7044, LUT_AMPL_WIDTH),
		30509 => to_signed(7041, LUT_AMPL_WIDTH),
		30510 => to_signed(7038, LUT_AMPL_WIDTH),
		30511 => to_signed(7035, LUT_AMPL_WIDTH),
		30512 => to_signed(7032, LUT_AMPL_WIDTH),
		30513 => to_signed(7029, LUT_AMPL_WIDTH),
		30514 => to_signed(7026, LUT_AMPL_WIDTH),
		30515 => to_signed(7023, LUT_AMPL_WIDTH),
		30516 => to_signed(7020, LUT_AMPL_WIDTH),
		30517 => to_signed(7017, LUT_AMPL_WIDTH),
		30518 => to_signed(7014, LUT_AMPL_WIDTH),
		30519 => to_signed(7011, LUT_AMPL_WIDTH),
		30520 => to_signed(7008, LUT_AMPL_WIDTH),
		30521 => to_signed(7004, LUT_AMPL_WIDTH),
		30522 => to_signed(7001, LUT_AMPL_WIDTH),
		30523 => to_signed(6998, LUT_AMPL_WIDTH),
		30524 => to_signed(6995, LUT_AMPL_WIDTH),
		30525 => to_signed(6992, LUT_AMPL_WIDTH),
		30526 => to_signed(6989, LUT_AMPL_WIDTH),
		30527 => to_signed(6986, LUT_AMPL_WIDTH),
		30528 => to_signed(6983, LUT_AMPL_WIDTH),
		30529 => to_signed(6980, LUT_AMPL_WIDTH),
		30530 => to_signed(6977, LUT_AMPL_WIDTH),
		30531 => to_signed(6974, LUT_AMPL_WIDTH),
		30532 => to_signed(6971, LUT_AMPL_WIDTH),
		30533 => to_signed(6968, LUT_AMPL_WIDTH),
		30534 => to_signed(6965, LUT_AMPL_WIDTH),
		30535 => to_signed(6961, LUT_AMPL_WIDTH),
		30536 => to_signed(6958, LUT_AMPL_WIDTH),
		30537 => to_signed(6955, LUT_AMPL_WIDTH),
		30538 => to_signed(6952, LUT_AMPL_WIDTH),
		30539 => to_signed(6949, LUT_AMPL_WIDTH),
		30540 => to_signed(6946, LUT_AMPL_WIDTH),
		30541 => to_signed(6943, LUT_AMPL_WIDTH),
		30542 => to_signed(6940, LUT_AMPL_WIDTH),
		30543 => to_signed(6937, LUT_AMPL_WIDTH),
		30544 => to_signed(6934, LUT_AMPL_WIDTH),
		30545 => to_signed(6931, LUT_AMPL_WIDTH),
		30546 => to_signed(6928, LUT_AMPL_WIDTH),
		30547 => to_signed(6925, LUT_AMPL_WIDTH),
		30548 => to_signed(6922, LUT_AMPL_WIDTH),
		30549 => to_signed(6919, LUT_AMPL_WIDTH),
		30550 => to_signed(6915, LUT_AMPL_WIDTH),
		30551 => to_signed(6912, LUT_AMPL_WIDTH),
		30552 => to_signed(6909, LUT_AMPL_WIDTH),
		30553 => to_signed(6906, LUT_AMPL_WIDTH),
		30554 => to_signed(6903, LUT_AMPL_WIDTH),
		30555 => to_signed(6900, LUT_AMPL_WIDTH),
		30556 => to_signed(6897, LUT_AMPL_WIDTH),
		30557 => to_signed(6894, LUT_AMPL_WIDTH),
		30558 => to_signed(6891, LUT_AMPL_WIDTH),
		30559 => to_signed(6888, LUT_AMPL_WIDTH),
		30560 => to_signed(6885, LUT_AMPL_WIDTH),
		30561 => to_signed(6882, LUT_AMPL_WIDTH),
		30562 => to_signed(6879, LUT_AMPL_WIDTH),
		30563 => to_signed(6876, LUT_AMPL_WIDTH),
		30564 => to_signed(6872, LUT_AMPL_WIDTH),
		30565 => to_signed(6869, LUT_AMPL_WIDTH),
		30566 => to_signed(6866, LUT_AMPL_WIDTH),
		30567 => to_signed(6863, LUT_AMPL_WIDTH),
		30568 => to_signed(6860, LUT_AMPL_WIDTH),
		30569 => to_signed(6857, LUT_AMPL_WIDTH),
		30570 => to_signed(6854, LUT_AMPL_WIDTH),
		30571 => to_signed(6851, LUT_AMPL_WIDTH),
		30572 => to_signed(6848, LUT_AMPL_WIDTH),
		30573 => to_signed(6845, LUT_AMPL_WIDTH),
		30574 => to_signed(6842, LUT_AMPL_WIDTH),
		30575 => to_signed(6839, LUT_AMPL_WIDTH),
		30576 => to_signed(6836, LUT_AMPL_WIDTH),
		30577 => to_signed(6833, LUT_AMPL_WIDTH),
		30578 => to_signed(6829, LUT_AMPL_WIDTH),
		30579 => to_signed(6826, LUT_AMPL_WIDTH),
		30580 => to_signed(6823, LUT_AMPL_WIDTH),
		30581 => to_signed(6820, LUT_AMPL_WIDTH),
		30582 => to_signed(6817, LUT_AMPL_WIDTH),
		30583 => to_signed(6814, LUT_AMPL_WIDTH),
		30584 => to_signed(6811, LUT_AMPL_WIDTH),
		30585 => to_signed(6808, LUT_AMPL_WIDTH),
		30586 => to_signed(6805, LUT_AMPL_WIDTH),
		30587 => to_signed(6802, LUT_AMPL_WIDTH),
		30588 => to_signed(6799, LUT_AMPL_WIDTH),
		30589 => to_signed(6796, LUT_AMPL_WIDTH),
		30590 => to_signed(6793, LUT_AMPL_WIDTH),
		30591 => to_signed(6789, LUT_AMPL_WIDTH),
		30592 => to_signed(6786, LUT_AMPL_WIDTH),
		30593 => to_signed(6783, LUT_AMPL_WIDTH),
		30594 => to_signed(6780, LUT_AMPL_WIDTH),
		30595 => to_signed(6777, LUT_AMPL_WIDTH),
		30596 => to_signed(6774, LUT_AMPL_WIDTH),
		30597 => to_signed(6771, LUT_AMPL_WIDTH),
		30598 => to_signed(6768, LUT_AMPL_WIDTH),
		30599 => to_signed(6765, LUT_AMPL_WIDTH),
		30600 => to_signed(6762, LUT_AMPL_WIDTH),
		30601 => to_signed(6759, LUT_AMPL_WIDTH),
		30602 => to_signed(6756, LUT_AMPL_WIDTH),
		30603 => to_signed(6753, LUT_AMPL_WIDTH),
		30604 => to_signed(6750, LUT_AMPL_WIDTH),
		30605 => to_signed(6746, LUT_AMPL_WIDTH),
		30606 => to_signed(6743, LUT_AMPL_WIDTH),
		30607 => to_signed(6740, LUT_AMPL_WIDTH),
		30608 => to_signed(6737, LUT_AMPL_WIDTH),
		30609 => to_signed(6734, LUT_AMPL_WIDTH),
		30610 => to_signed(6731, LUT_AMPL_WIDTH),
		30611 => to_signed(6728, LUT_AMPL_WIDTH),
		30612 => to_signed(6725, LUT_AMPL_WIDTH),
		30613 => to_signed(6722, LUT_AMPL_WIDTH),
		30614 => to_signed(6719, LUT_AMPL_WIDTH),
		30615 => to_signed(6716, LUT_AMPL_WIDTH),
		30616 => to_signed(6713, LUT_AMPL_WIDTH),
		30617 => to_signed(6710, LUT_AMPL_WIDTH),
		30618 => to_signed(6706, LUT_AMPL_WIDTH),
		30619 => to_signed(6703, LUT_AMPL_WIDTH),
		30620 => to_signed(6700, LUT_AMPL_WIDTH),
		30621 => to_signed(6697, LUT_AMPL_WIDTH),
		30622 => to_signed(6694, LUT_AMPL_WIDTH),
		30623 => to_signed(6691, LUT_AMPL_WIDTH),
		30624 => to_signed(6688, LUT_AMPL_WIDTH),
		30625 => to_signed(6685, LUT_AMPL_WIDTH),
		30626 => to_signed(6682, LUT_AMPL_WIDTH),
		30627 => to_signed(6679, LUT_AMPL_WIDTH),
		30628 => to_signed(6676, LUT_AMPL_WIDTH),
		30629 => to_signed(6673, LUT_AMPL_WIDTH),
		30630 => to_signed(6670, LUT_AMPL_WIDTH),
		30631 => to_signed(6667, LUT_AMPL_WIDTH),
		30632 => to_signed(6663, LUT_AMPL_WIDTH),
		30633 => to_signed(6660, LUT_AMPL_WIDTH),
		30634 => to_signed(6657, LUT_AMPL_WIDTH),
		30635 => to_signed(6654, LUT_AMPL_WIDTH),
		30636 => to_signed(6651, LUT_AMPL_WIDTH),
		30637 => to_signed(6648, LUT_AMPL_WIDTH),
		30638 => to_signed(6645, LUT_AMPL_WIDTH),
		30639 => to_signed(6642, LUT_AMPL_WIDTH),
		30640 => to_signed(6639, LUT_AMPL_WIDTH),
		30641 => to_signed(6636, LUT_AMPL_WIDTH),
		30642 => to_signed(6633, LUT_AMPL_WIDTH),
		30643 => to_signed(6630, LUT_AMPL_WIDTH),
		30644 => to_signed(6627, LUT_AMPL_WIDTH),
		30645 => to_signed(6623, LUT_AMPL_WIDTH),
		30646 => to_signed(6620, LUT_AMPL_WIDTH),
		30647 => to_signed(6617, LUT_AMPL_WIDTH),
		30648 => to_signed(6614, LUT_AMPL_WIDTH),
		30649 => to_signed(6611, LUT_AMPL_WIDTH),
		30650 => to_signed(6608, LUT_AMPL_WIDTH),
		30651 => to_signed(6605, LUT_AMPL_WIDTH),
		30652 => to_signed(6602, LUT_AMPL_WIDTH),
		30653 => to_signed(6599, LUT_AMPL_WIDTH),
		30654 => to_signed(6596, LUT_AMPL_WIDTH),
		30655 => to_signed(6593, LUT_AMPL_WIDTH),
		30656 => to_signed(6590, LUT_AMPL_WIDTH),
		30657 => to_signed(6587, LUT_AMPL_WIDTH),
		30658 => to_signed(6583, LUT_AMPL_WIDTH),
		30659 => to_signed(6580, LUT_AMPL_WIDTH),
		30660 => to_signed(6577, LUT_AMPL_WIDTH),
		30661 => to_signed(6574, LUT_AMPL_WIDTH),
		30662 => to_signed(6571, LUT_AMPL_WIDTH),
		30663 => to_signed(6568, LUT_AMPL_WIDTH),
		30664 => to_signed(6565, LUT_AMPL_WIDTH),
		30665 => to_signed(6562, LUT_AMPL_WIDTH),
		30666 => to_signed(6559, LUT_AMPL_WIDTH),
		30667 => to_signed(6556, LUT_AMPL_WIDTH),
		30668 => to_signed(6553, LUT_AMPL_WIDTH),
		30669 => to_signed(6550, LUT_AMPL_WIDTH),
		30670 => to_signed(6547, LUT_AMPL_WIDTH),
		30671 => to_signed(6543, LUT_AMPL_WIDTH),
		30672 => to_signed(6540, LUT_AMPL_WIDTH),
		30673 => to_signed(6537, LUT_AMPL_WIDTH),
		30674 => to_signed(6534, LUT_AMPL_WIDTH),
		30675 => to_signed(6531, LUT_AMPL_WIDTH),
		30676 => to_signed(6528, LUT_AMPL_WIDTH),
		30677 => to_signed(6525, LUT_AMPL_WIDTH),
		30678 => to_signed(6522, LUT_AMPL_WIDTH),
		30679 => to_signed(6519, LUT_AMPL_WIDTH),
		30680 => to_signed(6516, LUT_AMPL_WIDTH),
		30681 => to_signed(6513, LUT_AMPL_WIDTH),
		30682 => to_signed(6510, LUT_AMPL_WIDTH),
		30683 => to_signed(6506, LUT_AMPL_WIDTH),
		30684 => to_signed(6503, LUT_AMPL_WIDTH),
		30685 => to_signed(6500, LUT_AMPL_WIDTH),
		30686 => to_signed(6497, LUT_AMPL_WIDTH),
		30687 => to_signed(6494, LUT_AMPL_WIDTH),
		30688 => to_signed(6491, LUT_AMPL_WIDTH),
		30689 => to_signed(6488, LUT_AMPL_WIDTH),
		30690 => to_signed(6485, LUT_AMPL_WIDTH),
		30691 => to_signed(6482, LUT_AMPL_WIDTH),
		30692 => to_signed(6479, LUT_AMPL_WIDTH),
		30693 => to_signed(6476, LUT_AMPL_WIDTH),
		30694 => to_signed(6473, LUT_AMPL_WIDTH),
		30695 => to_signed(6470, LUT_AMPL_WIDTH),
		30696 => to_signed(6466, LUT_AMPL_WIDTH),
		30697 => to_signed(6463, LUT_AMPL_WIDTH),
		30698 => to_signed(6460, LUT_AMPL_WIDTH),
		30699 => to_signed(6457, LUT_AMPL_WIDTH),
		30700 => to_signed(6454, LUT_AMPL_WIDTH),
		30701 => to_signed(6451, LUT_AMPL_WIDTH),
		30702 => to_signed(6448, LUT_AMPL_WIDTH),
		30703 => to_signed(6445, LUT_AMPL_WIDTH),
		30704 => to_signed(6442, LUT_AMPL_WIDTH),
		30705 => to_signed(6439, LUT_AMPL_WIDTH),
		30706 => to_signed(6436, LUT_AMPL_WIDTH),
		30707 => to_signed(6433, LUT_AMPL_WIDTH),
		30708 => to_signed(6429, LUT_AMPL_WIDTH),
		30709 => to_signed(6426, LUT_AMPL_WIDTH),
		30710 => to_signed(6423, LUT_AMPL_WIDTH),
		30711 => to_signed(6420, LUT_AMPL_WIDTH),
		30712 => to_signed(6417, LUT_AMPL_WIDTH),
		30713 => to_signed(6414, LUT_AMPL_WIDTH),
		30714 => to_signed(6411, LUT_AMPL_WIDTH),
		30715 => to_signed(6408, LUT_AMPL_WIDTH),
		30716 => to_signed(6405, LUT_AMPL_WIDTH),
		30717 => to_signed(6402, LUT_AMPL_WIDTH),
		30718 => to_signed(6399, LUT_AMPL_WIDTH),
		30719 => to_signed(6396, LUT_AMPL_WIDTH),
		30720 => to_signed(6393, LUT_AMPL_WIDTH),
		30721 => to_signed(6389, LUT_AMPL_WIDTH),
		30722 => to_signed(6386, LUT_AMPL_WIDTH),
		30723 => to_signed(6383, LUT_AMPL_WIDTH),
		30724 => to_signed(6380, LUT_AMPL_WIDTH),
		30725 => to_signed(6377, LUT_AMPL_WIDTH),
		30726 => to_signed(6374, LUT_AMPL_WIDTH),
		30727 => to_signed(6371, LUT_AMPL_WIDTH),
		30728 => to_signed(6368, LUT_AMPL_WIDTH),
		30729 => to_signed(6365, LUT_AMPL_WIDTH),
		30730 => to_signed(6362, LUT_AMPL_WIDTH),
		30731 => to_signed(6359, LUT_AMPL_WIDTH),
		30732 => to_signed(6356, LUT_AMPL_WIDTH),
		30733 => to_signed(6352, LUT_AMPL_WIDTH),
		30734 => to_signed(6349, LUT_AMPL_WIDTH),
		30735 => to_signed(6346, LUT_AMPL_WIDTH),
		30736 => to_signed(6343, LUT_AMPL_WIDTH),
		30737 => to_signed(6340, LUT_AMPL_WIDTH),
		30738 => to_signed(6337, LUT_AMPL_WIDTH),
		30739 => to_signed(6334, LUT_AMPL_WIDTH),
		30740 => to_signed(6331, LUT_AMPL_WIDTH),
		30741 => to_signed(6328, LUT_AMPL_WIDTH),
		30742 => to_signed(6325, LUT_AMPL_WIDTH),
		30743 => to_signed(6322, LUT_AMPL_WIDTH),
		30744 => to_signed(6319, LUT_AMPL_WIDTH),
		30745 => to_signed(6315, LUT_AMPL_WIDTH),
		30746 => to_signed(6312, LUT_AMPL_WIDTH),
		30747 => to_signed(6309, LUT_AMPL_WIDTH),
		30748 => to_signed(6306, LUT_AMPL_WIDTH),
		30749 => to_signed(6303, LUT_AMPL_WIDTH),
		30750 => to_signed(6300, LUT_AMPL_WIDTH),
		30751 => to_signed(6297, LUT_AMPL_WIDTH),
		30752 => to_signed(6294, LUT_AMPL_WIDTH),
		30753 => to_signed(6291, LUT_AMPL_WIDTH),
		30754 => to_signed(6288, LUT_AMPL_WIDTH),
		30755 => to_signed(6285, LUT_AMPL_WIDTH),
		30756 => to_signed(6282, LUT_AMPL_WIDTH),
		30757 => to_signed(6278, LUT_AMPL_WIDTH),
		30758 => to_signed(6275, LUT_AMPL_WIDTH),
		30759 => to_signed(6272, LUT_AMPL_WIDTH),
		30760 => to_signed(6269, LUT_AMPL_WIDTH),
		30761 => to_signed(6266, LUT_AMPL_WIDTH),
		30762 => to_signed(6263, LUT_AMPL_WIDTH),
		30763 => to_signed(6260, LUT_AMPL_WIDTH),
		30764 => to_signed(6257, LUT_AMPL_WIDTH),
		30765 => to_signed(6254, LUT_AMPL_WIDTH),
		30766 => to_signed(6251, LUT_AMPL_WIDTH),
		30767 => to_signed(6248, LUT_AMPL_WIDTH),
		30768 => to_signed(6245, LUT_AMPL_WIDTH),
		30769 => to_signed(6241, LUT_AMPL_WIDTH),
		30770 => to_signed(6238, LUT_AMPL_WIDTH),
		30771 => to_signed(6235, LUT_AMPL_WIDTH),
		30772 => to_signed(6232, LUT_AMPL_WIDTH),
		30773 => to_signed(6229, LUT_AMPL_WIDTH),
		30774 => to_signed(6226, LUT_AMPL_WIDTH),
		30775 => to_signed(6223, LUT_AMPL_WIDTH),
		30776 => to_signed(6220, LUT_AMPL_WIDTH),
		30777 => to_signed(6217, LUT_AMPL_WIDTH),
		30778 => to_signed(6214, LUT_AMPL_WIDTH),
		30779 => to_signed(6211, LUT_AMPL_WIDTH),
		30780 => to_signed(6208, LUT_AMPL_WIDTH),
		30781 => to_signed(6204, LUT_AMPL_WIDTH),
		30782 => to_signed(6201, LUT_AMPL_WIDTH),
		30783 => to_signed(6198, LUT_AMPL_WIDTH),
		30784 => to_signed(6195, LUT_AMPL_WIDTH),
		30785 => to_signed(6192, LUT_AMPL_WIDTH),
		30786 => to_signed(6189, LUT_AMPL_WIDTH),
		30787 => to_signed(6186, LUT_AMPL_WIDTH),
		30788 => to_signed(6183, LUT_AMPL_WIDTH),
		30789 => to_signed(6180, LUT_AMPL_WIDTH),
		30790 => to_signed(6177, LUT_AMPL_WIDTH),
		30791 => to_signed(6174, LUT_AMPL_WIDTH),
		30792 => to_signed(6171, LUT_AMPL_WIDTH),
		30793 => to_signed(6167, LUT_AMPL_WIDTH),
		30794 => to_signed(6164, LUT_AMPL_WIDTH),
		30795 => to_signed(6161, LUT_AMPL_WIDTH),
		30796 => to_signed(6158, LUT_AMPL_WIDTH),
		30797 => to_signed(6155, LUT_AMPL_WIDTH),
		30798 => to_signed(6152, LUT_AMPL_WIDTH),
		30799 => to_signed(6149, LUT_AMPL_WIDTH),
		30800 => to_signed(6146, LUT_AMPL_WIDTH),
		30801 => to_signed(6143, LUT_AMPL_WIDTH),
		30802 => to_signed(6140, LUT_AMPL_WIDTH),
		30803 => to_signed(6137, LUT_AMPL_WIDTH),
		30804 => to_signed(6134, LUT_AMPL_WIDTH),
		30805 => to_signed(6130, LUT_AMPL_WIDTH),
		30806 => to_signed(6127, LUT_AMPL_WIDTH),
		30807 => to_signed(6124, LUT_AMPL_WIDTH),
		30808 => to_signed(6121, LUT_AMPL_WIDTH),
		30809 => to_signed(6118, LUT_AMPL_WIDTH),
		30810 => to_signed(6115, LUT_AMPL_WIDTH),
		30811 => to_signed(6112, LUT_AMPL_WIDTH),
		30812 => to_signed(6109, LUT_AMPL_WIDTH),
		30813 => to_signed(6106, LUT_AMPL_WIDTH),
		30814 => to_signed(6103, LUT_AMPL_WIDTH),
		30815 => to_signed(6100, LUT_AMPL_WIDTH),
		30816 => to_signed(6096, LUT_AMPL_WIDTH),
		30817 => to_signed(6093, LUT_AMPL_WIDTH),
		30818 => to_signed(6090, LUT_AMPL_WIDTH),
		30819 => to_signed(6087, LUT_AMPL_WIDTH),
		30820 => to_signed(6084, LUT_AMPL_WIDTH),
		30821 => to_signed(6081, LUT_AMPL_WIDTH),
		30822 => to_signed(6078, LUT_AMPL_WIDTH),
		30823 => to_signed(6075, LUT_AMPL_WIDTH),
		30824 => to_signed(6072, LUT_AMPL_WIDTH),
		30825 => to_signed(6069, LUT_AMPL_WIDTH),
		30826 => to_signed(6066, LUT_AMPL_WIDTH),
		30827 => to_signed(6063, LUT_AMPL_WIDTH),
		30828 => to_signed(6059, LUT_AMPL_WIDTH),
		30829 => to_signed(6056, LUT_AMPL_WIDTH),
		30830 => to_signed(6053, LUT_AMPL_WIDTH),
		30831 => to_signed(6050, LUT_AMPL_WIDTH),
		30832 => to_signed(6047, LUT_AMPL_WIDTH),
		30833 => to_signed(6044, LUT_AMPL_WIDTH),
		30834 => to_signed(6041, LUT_AMPL_WIDTH),
		30835 => to_signed(6038, LUT_AMPL_WIDTH),
		30836 => to_signed(6035, LUT_AMPL_WIDTH),
		30837 => to_signed(6032, LUT_AMPL_WIDTH),
		30838 => to_signed(6029, LUT_AMPL_WIDTH),
		30839 => to_signed(6025, LUT_AMPL_WIDTH),
		30840 => to_signed(6022, LUT_AMPL_WIDTH),
		30841 => to_signed(6019, LUT_AMPL_WIDTH),
		30842 => to_signed(6016, LUT_AMPL_WIDTH),
		30843 => to_signed(6013, LUT_AMPL_WIDTH),
		30844 => to_signed(6010, LUT_AMPL_WIDTH),
		30845 => to_signed(6007, LUT_AMPL_WIDTH),
		30846 => to_signed(6004, LUT_AMPL_WIDTH),
		30847 => to_signed(6001, LUT_AMPL_WIDTH),
		30848 => to_signed(5998, LUT_AMPL_WIDTH),
		30849 => to_signed(5995, LUT_AMPL_WIDTH),
		30850 => to_signed(5991, LUT_AMPL_WIDTH),
		30851 => to_signed(5988, LUT_AMPL_WIDTH),
		30852 => to_signed(5985, LUT_AMPL_WIDTH),
		30853 => to_signed(5982, LUT_AMPL_WIDTH),
		30854 => to_signed(5979, LUT_AMPL_WIDTH),
		30855 => to_signed(5976, LUT_AMPL_WIDTH),
		30856 => to_signed(5973, LUT_AMPL_WIDTH),
		30857 => to_signed(5970, LUT_AMPL_WIDTH),
		30858 => to_signed(5967, LUT_AMPL_WIDTH),
		30859 => to_signed(5964, LUT_AMPL_WIDTH),
		30860 => to_signed(5961, LUT_AMPL_WIDTH),
		30861 => to_signed(5958, LUT_AMPL_WIDTH),
		30862 => to_signed(5954, LUT_AMPL_WIDTH),
		30863 => to_signed(5951, LUT_AMPL_WIDTH),
		30864 => to_signed(5948, LUT_AMPL_WIDTH),
		30865 => to_signed(5945, LUT_AMPL_WIDTH),
		30866 => to_signed(5942, LUT_AMPL_WIDTH),
		30867 => to_signed(5939, LUT_AMPL_WIDTH),
		30868 => to_signed(5936, LUT_AMPL_WIDTH),
		30869 => to_signed(5933, LUT_AMPL_WIDTH),
		30870 => to_signed(5930, LUT_AMPL_WIDTH),
		30871 => to_signed(5927, LUT_AMPL_WIDTH),
		30872 => to_signed(5924, LUT_AMPL_WIDTH),
		30873 => to_signed(5920, LUT_AMPL_WIDTH),
		30874 => to_signed(5917, LUT_AMPL_WIDTH),
		30875 => to_signed(5914, LUT_AMPL_WIDTH),
		30876 => to_signed(5911, LUT_AMPL_WIDTH),
		30877 => to_signed(5908, LUT_AMPL_WIDTH),
		30878 => to_signed(5905, LUT_AMPL_WIDTH),
		30879 => to_signed(5902, LUT_AMPL_WIDTH),
		30880 => to_signed(5899, LUT_AMPL_WIDTH),
		30881 => to_signed(5896, LUT_AMPL_WIDTH),
		30882 => to_signed(5893, LUT_AMPL_WIDTH),
		30883 => to_signed(5890, LUT_AMPL_WIDTH),
		30884 => to_signed(5886, LUT_AMPL_WIDTH),
		30885 => to_signed(5883, LUT_AMPL_WIDTH),
		30886 => to_signed(5880, LUT_AMPL_WIDTH),
		30887 => to_signed(5877, LUT_AMPL_WIDTH),
		30888 => to_signed(5874, LUT_AMPL_WIDTH),
		30889 => to_signed(5871, LUT_AMPL_WIDTH),
		30890 => to_signed(5868, LUT_AMPL_WIDTH),
		30891 => to_signed(5865, LUT_AMPL_WIDTH),
		30892 => to_signed(5862, LUT_AMPL_WIDTH),
		30893 => to_signed(5859, LUT_AMPL_WIDTH),
		30894 => to_signed(5856, LUT_AMPL_WIDTH),
		30895 => to_signed(5852, LUT_AMPL_WIDTH),
		30896 => to_signed(5849, LUT_AMPL_WIDTH),
		30897 => to_signed(5846, LUT_AMPL_WIDTH),
		30898 => to_signed(5843, LUT_AMPL_WIDTH),
		30899 => to_signed(5840, LUT_AMPL_WIDTH),
		30900 => to_signed(5837, LUT_AMPL_WIDTH),
		30901 => to_signed(5834, LUT_AMPL_WIDTH),
		30902 => to_signed(5831, LUT_AMPL_WIDTH),
		30903 => to_signed(5828, LUT_AMPL_WIDTH),
		30904 => to_signed(5825, LUT_AMPL_WIDTH),
		30905 => to_signed(5822, LUT_AMPL_WIDTH),
		30906 => to_signed(5818, LUT_AMPL_WIDTH),
		30907 => to_signed(5815, LUT_AMPL_WIDTH),
		30908 => to_signed(5812, LUT_AMPL_WIDTH),
		30909 => to_signed(5809, LUT_AMPL_WIDTH),
		30910 => to_signed(5806, LUT_AMPL_WIDTH),
		30911 => to_signed(5803, LUT_AMPL_WIDTH),
		30912 => to_signed(5800, LUT_AMPL_WIDTH),
		30913 => to_signed(5797, LUT_AMPL_WIDTH),
		30914 => to_signed(5794, LUT_AMPL_WIDTH),
		30915 => to_signed(5791, LUT_AMPL_WIDTH),
		30916 => to_signed(5788, LUT_AMPL_WIDTH),
		30917 => to_signed(5784, LUT_AMPL_WIDTH),
		30918 => to_signed(5781, LUT_AMPL_WIDTH),
		30919 => to_signed(5778, LUT_AMPL_WIDTH),
		30920 => to_signed(5775, LUT_AMPL_WIDTH),
		30921 => to_signed(5772, LUT_AMPL_WIDTH),
		30922 => to_signed(5769, LUT_AMPL_WIDTH),
		30923 => to_signed(5766, LUT_AMPL_WIDTH),
		30924 => to_signed(5763, LUT_AMPL_WIDTH),
		30925 => to_signed(5760, LUT_AMPL_WIDTH),
		30926 => to_signed(5757, LUT_AMPL_WIDTH),
		30927 => to_signed(5754, LUT_AMPL_WIDTH),
		30928 => to_signed(5750, LUT_AMPL_WIDTH),
		30929 => to_signed(5747, LUT_AMPL_WIDTH),
		30930 => to_signed(5744, LUT_AMPL_WIDTH),
		30931 => to_signed(5741, LUT_AMPL_WIDTH),
		30932 => to_signed(5738, LUT_AMPL_WIDTH),
		30933 => to_signed(5735, LUT_AMPL_WIDTH),
		30934 => to_signed(5732, LUT_AMPL_WIDTH),
		30935 => to_signed(5729, LUT_AMPL_WIDTH),
		30936 => to_signed(5726, LUT_AMPL_WIDTH),
		30937 => to_signed(5723, LUT_AMPL_WIDTH),
		30938 => to_signed(5719, LUT_AMPL_WIDTH),
		30939 => to_signed(5716, LUT_AMPL_WIDTH),
		30940 => to_signed(5713, LUT_AMPL_WIDTH),
		30941 => to_signed(5710, LUT_AMPL_WIDTH),
		30942 => to_signed(5707, LUT_AMPL_WIDTH),
		30943 => to_signed(5704, LUT_AMPL_WIDTH),
		30944 => to_signed(5701, LUT_AMPL_WIDTH),
		30945 => to_signed(5698, LUT_AMPL_WIDTH),
		30946 => to_signed(5695, LUT_AMPL_WIDTH),
		30947 => to_signed(5692, LUT_AMPL_WIDTH),
		30948 => to_signed(5689, LUT_AMPL_WIDTH),
		30949 => to_signed(5685, LUT_AMPL_WIDTH),
		30950 => to_signed(5682, LUT_AMPL_WIDTH),
		30951 => to_signed(5679, LUT_AMPL_WIDTH),
		30952 => to_signed(5676, LUT_AMPL_WIDTH),
		30953 => to_signed(5673, LUT_AMPL_WIDTH),
		30954 => to_signed(5670, LUT_AMPL_WIDTH),
		30955 => to_signed(5667, LUT_AMPL_WIDTH),
		30956 => to_signed(5664, LUT_AMPL_WIDTH),
		30957 => to_signed(5661, LUT_AMPL_WIDTH),
		30958 => to_signed(5658, LUT_AMPL_WIDTH),
		30959 => to_signed(5655, LUT_AMPL_WIDTH),
		30960 => to_signed(5651, LUT_AMPL_WIDTH),
		30961 => to_signed(5648, LUT_AMPL_WIDTH),
		30962 => to_signed(5645, LUT_AMPL_WIDTH),
		30963 => to_signed(5642, LUT_AMPL_WIDTH),
		30964 => to_signed(5639, LUT_AMPL_WIDTH),
		30965 => to_signed(5636, LUT_AMPL_WIDTH),
		30966 => to_signed(5633, LUT_AMPL_WIDTH),
		30967 => to_signed(5630, LUT_AMPL_WIDTH),
		30968 => to_signed(5627, LUT_AMPL_WIDTH),
		30969 => to_signed(5624, LUT_AMPL_WIDTH),
		30970 => to_signed(5620, LUT_AMPL_WIDTH),
		30971 => to_signed(5617, LUT_AMPL_WIDTH),
		30972 => to_signed(5614, LUT_AMPL_WIDTH),
		30973 => to_signed(5611, LUT_AMPL_WIDTH),
		30974 => to_signed(5608, LUT_AMPL_WIDTH),
		30975 => to_signed(5605, LUT_AMPL_WIDTH),
		30976 => to_signed(5602, LUT_AMPL_WIDTH),
		30977 => to_signed(5599, LUT_AMPL_WIDTH),
		30978 => to_signed(5596, LUT_AMPL_WIDTH),
		30979 => to_signed(5593, LUT_AMPL_WIDTH),
		30980 => to_signed(5590, LUT_AMPL_WIDTH),
		30981 => to_signed(5586, LUT_AMPL_WIDTH),
		30982 => to_signed(5583, LUT_AMPL_WIDTH),
		30983 => to_signed(5580, LUT_AMPL_WIDTH),
		30984 => to_signed(5577, LUT_AMPL_WIDTH),
		30985 => to_signed(5574, LUT_AMPL_WIDTH),
		30986 => to_signed(5571, LUT_AMPL_WIDTH),
		30987 => to_signed(5568, LUT_AMPL_WIDTH),
		30988 => to_signed(5565, LUT_AMPL_WIDTH),
		30989 => to_signed(5562, LUT_AMPL_WIDTH),
		30990 => to_signed(5559, LUT_AMPL_WIDTH),
		30991 => to_signed(5555, LUT_AMPL_WIDTH),
		30992 => to_signed(5552, LUT_AMPL_WIDTH),
		30993 => to_signed(5549, LUT_AMPL_WIDTH),
		30994 => to_signed(5546, LUT_AMPL_WIDTH),
		30995 => to_signed(5543, LUT_AMPL_WIDTH),
		30996 => to_signed(5540, LUT_AMPL_WIDTH),
		30997 => to_signed(5537, LUT_AMPL_WIDTH),
		30998 => to_signed(5534, LUT_AMPL_WIDTH),
		30999 => to_signed(5531, LUT_AMPL_WIDTH),
		31000 => to_signed(5528, LUT_AMPL_WIDTH),
		31001 => to_signed(5525, LUT_AMPL_WIDTH),
		31002 => to_signed(5521, LUT_AMPL_WIDTH),
		31003 => to_signed(5518, LUT_AMPL_WIDTH),
		31004 => to_signed(5515, LUT_AMPL_WIDTH),
		31005 => to_signed(5512, LUT_AMPL_WIDTH),
		31006 => to_signed(5509, LUT_AMPL_WIDTH),
		31007 => to_signed(5506, LUT_AMPL_WIDTH),
		31008 => to_signed(5503, LUT_AMPL_WIDTH),
		31009 => to_signed(5500, LUT_AMPL_WIDTH),
		31010 => to_signed(5497, LUT_AMPL_WIDTH),
		31011 => to_signed(5494, LUT_AMPL_WIDTH),
		31012 => to_signed(5490, LUT_AMPL_WIDTH),
		31013 => to_signed(5487, LUT_AMPL_WIDTH),
		31014 => to_signed(5484, LUT_AMPL_WIDTH),
		31015 => to_signed(5481, LUT_AMPL_WIDTH),
		31016 => to_signed(5478, LUT_AMPL_WIDTH),
		31017 => to_signed(5475, LUT_AMPL_WIDTH),
		31018 => to_signed(5472, LUT_AMPL_WIDTH),
		31019 => to_signed(5469, LUT_AMPL_WIDTH),
		31020 => to_signed(5466, LUT_AMPL_WIDTH),
		31021 => to_signed(5463, LUT_AMPL_WIDTH),
		31022 => to_signed(5459, LUT_AMPL_WIDTH),
		31023 => to_signed(5456, LUT_AMPL_WIDTH),
		31024 => to_signed(5453, LUT_AMPL_WIDTH),
		31025 => to_signed(5450, LUT_AMPL_WIDTH),
		31026 => to_signed(5447, LUT_AMPL_WIDTH),
		31027 => to_signed(5444, LUT_AMPL_WIDTH),
		31028 => to_signed(5441, LUT_AMPL_WIDTH),
		31029 => to_signed(5438, LUT_AMPL_WIDTH),
		31030 => to_signed(5435, LUT_AMPL_WIDTH),
		31031 => to_signed(5432, LUT_AMPL_WIDTH),
		31032 => to_signed(5428, LUT_AMPL_WIDTH),
		31033 => to_signed(5425, LUT_AMPL_WIDTH),
		31034 => to_signed(5422, LUT_AMPL_WIDTH),
		31035 => to_signed(5419, LUT_AMPL_WIDTH),
		31036 => to_signed(5416, LUT_AMPL_WIDTH),
		31037 => to_signed(5413, LUT_AMPL_WIDTH),
		31038 => to_signed(5410, LUT_AMPL_WIDTH),
		31039 => to_signed(5407, LUT_AMPL_WIDTH),
		31040 => to_signed(5404, LUT_AMPL_WIDTH),
		31041 => to_signed(5401, LUT_AMPL_WIDTH),
		31042 => to_signed(5398, LUT_AMPL_WIDTH),
		31043 => to_signed(5394, LUT_AMPL_WIDTH),
		31044 => to_signed(5391, LUT_AMPL_WIDTH),
		31045 => to_signed(5388, LUT_AMPL_WIDTH),
		31046 => to_signed(5385, LUT_AMPL_WIDTH),
		31047 => to_signed(5382, LUT_AMPL_WIDTH),
		31048 => to_signed(5379, LUT_AMPL_WIDTH),
		31049 => to_signed(5376, LUT_AMPL_WIDTH),
		31050 => to_signed(5373, LUT_AMPL_WIDTH),
		31051 => to_signed(5370, LUT_AMPL_WIDTH),
		31052 => to_signed(5367, LUT_AMPL_WIDTH),
		31053 => to_signed(5363, LUT_AMPL_WIDTH),
		31054 => to_signed(5360, LUT_AMPL_WIDTH),
		31055 => to_signed(5357, LUT_AMPL_WIDTH),
		31056 => to_signed(5354, LUT_AMPL_WIDTH),
		31057 => to_signed(5351, LUT_AMPL_WIDTH),
		31058 => to_signed(5348, LUT_AMPL_WIDTH),
		31059 => to_signed(5345, LUT_AMPL_WIDTH),
		31060 => to_signed(5342, LUT_AMPL_WIDTH),
		31061 => to_signed(5339, LUT_AMPL_WIDTH),
		31062 => to_signed(5336, LUT_AMPL_WIDTH),
		31063 => to_signed(5332, LUT_AMPL_WIDTH),
		31064 => to_signed(5329, LUT_AMPL_WIDTH),
		31065 => to_signed(5326, LUT_AMPL_WIDTH),
		31066 => to_signed(5323, LUT_AMPL_WIDTH),
		31067 => to_signed(5320, LUT_AMPL_WIDTH),
		31068 => to_signed(5317, LUT_AMPL_WIDTH),
		31069 => to_signed(5314, LUT_AMPL_WIDTH),
		31070 => to_signed(5311, LUT_AMPL_WIDTH),
		31071 => to_signed(5308, LUT_AMPL_WIDTH),
		31072 => to_signed(5305, LUT_AMPL_WIDTH),
		31073 => to_signed(5301, LUT_AMPL_WIDTH),
		31074 => to_signed(5298, LUT_AMPL_WIDTH),
		31075 => to_signed(5295, LUT_AMPL_WIDTH),
		31076 => to_signed(5292, LUT_AMPL_WIDTH),
		31077 => to_signed(5289, LUT_AMPL_WIDTH),
		31078 => to_signed(5286, LUT_AMPL_WIDTH),
		31079 => to_signed(5283, LUT_AMPL_WIDTH),
		31080 => to_signed(5280, LUT_AMPL_WIDTH),
		31081 => to_signed(5277, LUT_AMPL_WIDTH),
		31082 => to_signed(5274, LUT_AMPL_WIDTH),
		31083 => to_signed(5270, LUT_AMPL_WIDTH),
		31084 => to_signed(5267, LUT_AMPL_WIDTH),
		31085 => to_signed(5264, LUT_AMPL_WIDTH),
		31086 => to_signed(5261, LUT_AMPL_WIDTH),
		31087 => to_signed(5258, LUT_AMPL_WIDTH),
		31088 => to_signed(5255, LUT_AMPL_WIDTH),
		31089 => to_signed(5252, LUT_AMPL_WIDTH),
		31090 => to_signed(5249, LUT_AMPL_WIDTH),
		31091 => to_signed(5246, LUT_AMPL_WIDTH),
		31092 => to_signed(5243, LUT_AMPL_WIDTH),
		31093 => to_signed(5239, LUT_AMPL_WIDTH),
		31094 => to_signed(5236, LUT_AMPL_WIDTH),
		31095 => to_signed(5233, LUT_AMPL_WIDTH),
		31096 => to_signed(5230, LUT_AMPL_WIDTH),
		31097 => to_signed(5227, LUT_AMPL_WIDTH),
		31098 => to_signed(5224, LUT_AMPL_WIDTH),
		31099 => to_signed(5221, LUT_AMPL_WIDTH),
		31100 => to_signed(5218, LUT_AMPL_WIDTH),
		31101 => to_signed(5215, LUT_AMPL_WIDTH),
		31102 => to_signed(5212, LUT_AMPL_WIDTH),
		31103 => to_signed(5208, LUT_AMPL_WIDTH),
		31104 => to_signed(5205, LUT_AMPL_WIDTH),
		31105 => to_signed(5202, LUT_AMPL_WIDTH),
		31106 => to_signed(5199, LUT_AMPL_WIDTH),
		31107 => to_signed(5196, LUT_AMPL_WIDTH),
		31108 => to_signed(5193, LUT_AMPL_WIDTH),
		31109 => to_signed(5190, LUT_AMPL_WIDTH),
		31110 => to_signed(5187, LUT_AMPL_WIDTH),
		31111 => to_signed(5184, LUT_AMPL_WIDTH),
		31112 => to_signed(5180, LUT_AMPL_WIDTH),
		31113 => to_signed(5177, LUT_AMPL_WIDTH),
		31114 => to_signed(5174, LUT_AMPL_WIDTH),
		31115 => to_signed(5171, LUT_AMPL_WIDTH),
		31116 => to_signed(5168, LUT_AMPL_WIDTH),
		31117 => to_signed(5165, LUT_AMPL_WIDTH),
		31118 => to_signed(5162, LUT_AMPL_WIDTH),
		31119 => to_signed(5159, LUT_AMPL_WIDTH),
		31120 => to_signed(5156, LUT_AMPL_WIDTH),
		31121 => to_signed(5153, LUT_AMPL_WIDTH),
		31122 => to_signed(5149, LUT_AMPL_WIDTH),
		31123 => to_signed(5146, LUT_AMPL_WIDTH),
		31124 => to_signed(5143, LUT_AMPL_WIDTH),
		31125 => to_signed(5140, LUT_AMPL_WIDTH),
		31126 => to_signed(5137, LUT_AMPL_WIDTH),
		31127 => to_signed(5134, LUT_AMPL_WIDTH),
		31128 => to_signed(5131, LUT_AMPL_WIDTH),
		31129 => to_signed(5128, LUT_AMPL_WIDTH),
		31130 => to_signed(5125, LUT_AMPL_WIDTH),
		31131 => to_signed(5122, LUT_AMPL_WIDTH),
		31132 => to_signed(5118, LUT_AMPL_WIDTH),
		31133 => to_signed(5115, LUT_AMPL_WIDTH),
		31134 => to_signed(5112, LUT_AMPL_WIDTH),
		31135 => to_signed(5109, LUT_AMPL_WIDTH),
		31136 => to_signed(5106, LUT_AMPL_WIDTH),
		31137 => to_signed(5103, LUT_AMPL_WIDTH),
		31138 => to_signed(5100, LUT_AMPL_WIDTH),
		31139 => to_signed(5097, LUT_AMPL_WIDTH),
		31140 => to_signed(5094, LUT_AMPL_WIDTH),
		31141 => to_signed(5091, LUT_AMPL_WIDTH),
		31142 => to_signed(5087, LUT_AMPL_WIDTH),
		31143 => to_signed(5084, LUT_AMPL_WIDTH),
		31144 => to_signed(5081, LUT_AMPL_WIDTH),
		31145 => to_signed(5078, LUT_AMPL_WIDTH),
		31146 => to_signed(5075, LUT_AMPL_WIDTH),
		31147 => to_signed(5072, LUT_AMPL_WIDTH),
		31148 => to_signed(5069, LUT_AMPL_WIDTH),
		31149 => to_signed(5066, LUT_AMPL_WIDTH),
		31150 => to_signed(5063, LUT_AMPL_WIDTH),
		31151 => to_signed(5059, LUT_AMPL_WIDTH),
		31152 => to_signed(5056, LUT_AMPL_WIDTH),
		31153 => to_signed(5053, LUT_AMPL_WIDTH),
		31154 => to_signed(5050, LUT_AMPL_WIDTH),
		31155 => to_signed(5047, LUT_AMPL_WIDTH),
		31156 => to_signed(5044, LUT_AMPL_WIDTH),
		31157 => to_signed(5041, LUT_AMPL_WIDTH),
		31158 => to_signed(5038, LUT_AMPL_WIDTH),
		31159 => to_signed(5035, LUT_AMPL_WIDTH),
		31160 => to_signed(5032, LUT_AMPL_WIDTH),
		31161 => to_signed(5028, LUT_AMPL_WIDTH),
		31162 => to_signed(5025, LUT_AMPL_WIDTH),
		31163 => to_signed(5022, LUT_AMPL_WIDTH),
		31164 => to_signed(5019, LUT_AMPL_WIDTH),
		31165 => to_signed(5016, LUT_AMPL_WIDTH),
		31166 => to_signed(5013, LUT_AMPL_WIDTH),
		31167 => to_signed(5010, LUT_AMPL_WIDTH),
		31168 => to_signed(5007, LUT_AMPL_WIDTH),
		31169 => to_signed(5004, LUT_AMPL_WIDTH),
		31170 => to_signed(5000, LUT_AMPL_WIDTH),
		31171 => to_signed(4997, LUT_AMPL_WIDTH),
		31172 => to_signed(4994, LUT_AMPL_WIDTH),
		31173 => to_signed(4991, LUT_AMPL_WIDTH),
		31174 => to_signed(4988, LUT_AMPL_WIDTH),
		31175 => to_signed(4985, LUT_AMPL_WIDTH),
		31176 => to_signed(4982, LUT_AMPL_WIDTH),
		31177 => to_signed(4979, LUT_AMPL_WIDTH),
		31178 => to_signed(4976, LUT_AMPL_WIDTH),
		31179 => to_signed(4973, LUT_AMPL_WIDTH),
		31180 => to_signed(4969, LUT_AMPL_WIDTH),
		31181 => to_signed(4966, LUT_AMPL_WIDTH),
		31182 => to_signed(4963, LUT_AMPL_WIDTH),
		31183 => to_signed(4960, LUT_AMPL_WIDTH),
		31184 => to_signed(4957, LUT_AMPL_WIDTH),
		31185 => to_signed(4954, LUT_AMPL_WIDTH),
		31186 => to_signed(4951, LUT_AMPL_WIDTH),
		31187 => to_signed(4948, LUT_AMPL_WIDTH),
		31188 => to_signed(4945, LUT_AMPL_WIDTH),
		31189 => to_signed(4941, LUT_AMPL_WIDTH),
		31190 => to_signed(4938, LUT_AMPL_WIDTH),
		31191 => to_signed(4935, LUT_AMPL_WIDTH),
		31192 => to_signed(4932, LUT_AMPL_WIDTH),
		31193 => to_signed(4929, LUT_AMPL_WIDTH),
		31194 => to_signed(4926, LUT_AMPL_WIDTH),
		31195 => to_signed(4923, LUT_AMPL_WIDTH),
		31196 => to_signed(4920, LUT_AMPL_WIDTH),
		31197 => to_signed(4917, LUT_AMPL_WIDTH),
		31198 => to_signed(4914, LUT_AMPL_WIDTH),
		31199 => to_signed(4910, LUT_AMPL_WIDTH),
		31200 => to_signed(4907, LUT_AMPL_WIDTH),
		31201 => to_signed(4904, LUT_AMPL_WIDTH),
		31202 => to_signed(4901, LUT_AMPL_WIDTH),
		31203 => to_signed(4898, LUT_AMPL_WIDTH),
		31204 => to_signed(4895, LUT_AMPL_WIDTH),
		31205 => to_signed(4892, LUT_AMPL_WIDTH),
		31206 => to_signed(4889, LUT_AMPL_WIDTH),
		31207 => to_signed(4886, LUT_AMPL_WIDTH),
		31208 => to_signed(4882, LUT_AMPL_WIDTH),
		31209 => to_signed(4879, LUT_AMPL_WIDTH),
		31210 => to_signed(4876, LUT_AMPL_WIDTH),
		31211 => to_signed(4873, LUT_AMPL_WIDTH),
		31212 => to_signed(4870, LUT_AMPL_WIDTH),
		31213 => to_signed(4867, LUT_AMPL_WIDTH),
		31214 => to_signed(4864, LUT_AMPL_WIDTH),
		31215 => to_signed(4861, LUT_AMPL_WIDTH),
		31216 => to_signed(4858, LUT_AMPL_WIDTH),
		31217 => to_signed(4855, LUT_AMPL_WIDTH),
		31218 => to_signed(4851, LUT_AMPL_WIDTH),
		31219 => to_signed(4848, LUT_AMPL_WIDTH),
		31220 => to_signed(4845, LUT_AMPL_WIDTH),
		31221 => to_signed(4842, LUT_AMPL_WIDTH),
		31222 => to_signed(4839, LUT_AMPL_WIDTH),
		31223 => to_signed(4836, LUT_AMPL_WIDTH),
		31224 => to_signed(4833, LUT_AMPL_WIDTH),
		31225 => to_signed(4830, LUT_AMPL_WIDTH),
		31226 => to_signed(4827, LUT_AMPL_WIDTH),
		31227 => to_signed(4823, LUT_AMPL_WIDTH),
		31228 => to_signed(4820, LUT_AMPL_WIDTH),
		31229 => to_signed(4817, LUT_AMPL_WIDTH),
		31230 => to_signed(4814, LUT_AMPL_WIDTH),
		31231 => to_signed(4811, LUT_AMPL_WIDTH),
		31232 => to_signed(4808, LUT_AMPL_WIDTH),
		31233 => to_signed(4805, LUT_AMPL_WIDTH),
		31234 => to_signed(4802, LUT_AMPL_WIDTH),
		31235 => to_signed(4799, LUT_AMPL_WIDTH),
		31236 => to_signed(4795, LUT_AMPL_WIDTH),
		31237 => to_signed(4792, LUT_AMPL_WIDTH),
		31238 => to_signed(4789, LUT_AMPL_WIDTH),
		31239 => to_signed(4786, LUT_AMPL_WIDTH),
		31240 => to_signed(4783, LUT_AMPL_WIDTH),
		31241 => to_signed(4780, LUT_AMPL_WIDTH),
		31242 => to_signed(4777, LUT_AMPL_WIDTH),
		31243 => to_signed(4774, LUT_AMPL_WIDTH),
		31244 => to_signed(4771, LUT_AMPL_WIDTH),
		31245 => to_signed(4768, LUT_AMPL_WIDTH),
		31246 => to_signed(4764, LUT_AMPL_WIDTH),
		31247 => to_signed(4761, LUT_AMPL_WIDTH),
		31248 => to_signed(4758, LUT_AMPL_WIDTH),
		31249 => to_signed(4755, LUT_AMPL_WIDTH),
		31250 => to_signed(4752, LUT_AMPL_WIDTH),
		31251 => to_signed(4749, LUT_AMPL_WIDTH),
		31252 => to_signed(4746, LUT_AMPL_WIDTH),
		31253 => to_signed(4743, LUT_AMPL_WIDTH),
		31254 => to_signed(4740, LUT_AMPL_WIDTH),
		31255 => to_signed(4736, LUT_AMPL_WIDTH),
		31256 => to_signed(4733, LUT_AMPL_WIDTH),
		31257 => to_signed(4730, LUT_AMPL_WIDTH),
		31258 => to_signed(4727, LUT_AMPL_WIDTH),
		31259 => to_signed(4724, LUT_AMPL_WIDTH),
		31260 => to_signed(4721, LUT_AMPL_WIDTH),
		31261 => to_signed(4718, LUT_AMPL_WIDTH),
		31262 => to_signed(4715, LUT_AMPL_WIDTH),
		31263 => to_signed(4712, LUT_AMPL_WIDTH),
		31264 => to_signed(4708, LUT_AMPL_WIDTH),
		31265 => to_signed(4705, LUT_AMPL_WIDTH),
		31266 => to_signed(4702, LUT_AMPL_WIDTH),
		31267 => to_signed(4699, LUT_AMPL_WIDTH),
		31268 => to_signed(4696, LUT_AMPL_WIDTH),
		31269 => to_signed(4693, LUT_AMPL_WIDTH),
		31270 => to_signed(4690, LUT_AMPL_WIDTH),
		31271 => to_signed(4687, LUT_AMPL_WIDTH),
		31272 => to_signed(4684, LUT_AMPL_WIDTH),
		31273 => to_signed(4680, LUT_AMPL_WIDTH),
		31274 => to_signed(4677, LUT_AMPL_WIDTH),
		31275 => to_signed(4674, LUT_AMPL_WIDTH),
		31276 => to_signed(4671, LUT_AMPL_WIDTH),
		31277 => to_signed(4668, LUT_AMPL_WIDTH),
		31278 => to_signed(4665, LUT_AMPL_WIDTH),
		31279 => to_signed(4662, LUT_AMPL_WIDTH),
		31280 => to_signed(4659, LUT_AMPL_WIDTH),
		31281 => to_signed(4656, LUT_AMPL_WIDTH),
		31282 => to_signed(4652, LUT_AMPL_WIDTH),
		31283 => to_signed(4649, LUT_AMPL_WIDTH),
		31284 => to_signed(4646, LUT_AMPL_WIDTH),
		31285 => to_signed(4643, LUT_AMPL_WIDTH),
		31286 => to_signed(4640, LUT_AMPL_WIDTH),
		31287 => to_signed(4637, LUT_AMPL_WIDTH),
		31288 => to_signed(4634, LUT_AMPL_WIDTH),
		31289 => to_signed(4631, LUT_AMPL_WIDTH),
		31290 => to_signed(4628, LUT_AMPL_WIDTH),
		31291 => to_signed(4624, LUT_AMPL_WIDTH),
		31292 => to_signed(4621, LUT_AMPL_WIDTH),
		31293 => to_signed(4618, LUT_AMPL_WIDTH),
		31294 => to_signed(4615, LUT_AMPL_WIDTH),
		31295 => to_signed(4612, LUT_AMPL_WIDTH),
		31296 => to_signed(4609, LUT_AMPL_WIDTH),
		31297 => to_signed(4606, LUT_AMPL_WIDTH),
		31298 => to_signed(4603, LUT_AMPL_WIDTH),
		31299 => to_signed(4600, LUT_AMPL_WIDTH),
		31300 => to_signed(4597, LUT_AMPL_WIDTH),
		31301 => to_signed(4593, LUT_AMPL_WIDTH),
		31302 => to_signed(4590, LUT_AMPL_WIDTH),
		31303 => to_signed(4587, LUT_AMPL_WIDTH),
		31304 => to_signed(4584, LUT_AMPL_WIDTH),
		31305 => to_signed(4581, LUT_AMPL_WIDTH),
		31306 => to_signed(4578, LUT_AMPL_WIDTH),
		31307 => to_signed(4575, LUT_AMPL_WIDTH),
		31308 => to_signed(4572, LUT_AMPL_WIDTH),
		31309 => to_signed(4569, LUT_AMPL_WIDTH),
		31310 => to_signed(4565, LUT_AMPL_WIDTH),
		31311 => to_signed(4562, LUT_AMPL_WIDTH),
		31312 => to_signed(4559, LUT_AMPL_WIDTH),
		31313 => to_signed(4556, LUT_AMPL_WIDTH),
		31314 => to_signed(4553, LUT_AMPL_WIDTH),
		31315 => to_signed(4550, LUT_AMPL_WIDTH),
		31316 => to_signed(4547, LUT_AMPL_WIDTH),
		31317 => to_signed(4544, LUT_AMPL_WIDTH),
		31318 => to_signed(4541, LUT_AMPL_WIDTH),
		31319 => to_signed(4537, LUT_AMPL_WIDTH),
		31320 => to_signed(4534, LUT_AMPL_WIDTH),
		31321 => to_signed(4531, LUT_AMPL_WIDTH),
		31322 => to_signed(4528, LUT_AMPL_WIDTH),
		31323 => to_signed(4525, LUT_AMPL_WIDTH),
		31324 => to_signed(4522, LUT_AMPL_WIDTH),
		31325 => to_signed(4519, LUT_AMPL_WIDTH),
		31326 => to_signed(4516, LUT_AMPL_WIDTH),
		31327 => to_signed(4513, LUT_AMPL_WIDTH),
		31328 => to_signed(4509, LUT_AMPL_WIDTH),
		31329 => to_signed(4506, LUT_AMPL_WIDTH),
		31330 => to_signed(4503, LUT_AMPL_WIDTH),
		31331 => to_signed(4500, LUT_AMPL_WIDTH),
		31332 => to_signed(4497, LUT_AMPL_WIDTH),
		31333 => to_signed(4494, LUT_AMPL_WIDTH),
		31334 => to_signed(4491, LUT_AMPL_WIDTH),
		31335 => to_signed(4488, LUT_AMPL_WIDTH),
		31336 => to_signed(4485, LUT_AMPL_WIDTH),
		31337 => to_signed(4481, LUT_AMPL_WIDTH),
		31338 => to_signed(4478, LUT_AMPL_WIDTH),
		31339 => to_signed(4475, LUT_AMPL_WIDTH),
		31340 => to_signed(4472, LUT_AMPL_WIDTH),
		31341 => to_signed(4469, LUT_AMPL_WIDTH),
		31342 => to_signed(4466, LUT_AMPL_WIDTH),
		31343 => to_signed(4463, LUT_AMPL_WIDTH),
		31344 => to_signed(4460, LUT_AMPL_WIDTH),
		31345 => to_signed(4456, LUT_AMPL_WIDTH),
		31346 => to_signed(4453, LUT_AMPL_WIDTH),
		31347 => to_signed(4450, LUT_AMPL_WIDTH),
		31348 => to_signed(4447, LUT_AMPL_WIDTH),
		31349 => to_signed(4444, LUT_AMPL_WIDTH),
		31350 => to_signed(4441, LUT_AMPL_WIDTH),
		31351 => to_signed(4438, LUT_AMPL_WIDTH),
		31352 => to_signed(4435, LUT_AMPL_WIDTH),
		31353 => to_signed(4432, LUT_AMPL_WIDTH),
		31354 => to_signed(4428, LUT_AMPL_WIDTH),
		31355 => to_signed(4425, LUT_AMPL_WIDTH),
		31356 => to_signed(4422, LUT_AMPL_WIDTH),
		31357 => to_signed(4419, LUT_AMPL_WIDTH),
		31358 => to_signed(4416, LUT_AMPL_WIDTH),
		31359 => to_signed(4413, LUT_AMPL_WIDTH),
		31360 => to_signed(4410, LUT_AMPL_WIDTH),
		31361 => to_signed(4407, LUT_AMPL_WIDTH),
		31362 => to_signed(4404, LUT_AMPL_WIDTH),
		31363 => to_signed(4400, LUT_AMPL_WIDTH),
		31364 => to_signed(4397, LUT_AMPL_WIDTH),
		31365 => to_signed(4394, LUT_AMPL_WIDTH),
		31366 => to_signed(4391, LUT_AMPL_WIDTH),
		31367 => to_signed(4388, LUT_AMPL_WIDTH),
		31368 => to_signed(4385, LUT_AMPL_WIDTH),
		31369 => to_signed(4382, LUT_AMPL_WIDTH),
		31370 => to_signed(4379, LUT_AMPL_WIDTH),
		31371 => to_signed(4376, LUT_AMPL_WIDTH),
		31372 => to_signed(4372, LUT_AMPL_WIDTH),
		31373 => to_signed(4369, LUT_AMPL_WIDTH),
		31374 => to_signed(4366, LUT_AMPL_WIDTH),
		31375 => to_signed(4363, LUT_AMPL_WIDTH),
		31376 => to_signed(4360, LUT_AMPL_WIDTH),
		31377 => to_signed(4357, LUT_AMPL_WIDTH),
		31378 => to_signed(4354, LUT_AMPL_WIDTH),
		31379 => to_signed(4351, LUT_AMPL_WIDTH),
		31380 => to_signed(4348, LUT_AMPL_WIDTH),
		31381 => to_signed(4344, LUT_AMPL_WIDTH),
		31382 => to_signed(4341, LUT_AMPL_WIDTH),
		31383 => to_signed(4338, LUT_AMPL_WIDTH),
		31384 => to_signed(4335, LUT_AMPL_WIDTH),
		31385 => to_signed(4332, LUT_AMPL_WIDTH),
		31386 => to_signed(4329, LUT_AMPL_WIDTH),
		31387 => to_signed(4326, LUT_AMPL_WIDTH),
		31388 => to_signed(4323, LUT_AMPL_WIDTH),
		31389 => to_signed(4320, LUT_AMPL_WIDTH),
		31390 => to_signed(4316, LUT_AMPL_WIDTH),
		31391 => to_signed(4313, LUT_AMPL_WIDTH),
		31392 => to_signed(4310, LUT_AMPL_WIDTH),
		31393 => to_signed(4307, LUT_AMPL_WIDTH),
		31394 => to_signed(4304, LUT_AMPL_WIDTH),
		31395 => to_signed(4301, LUT_AMPL_WIDTH),
		31396 => to_signed(4298, LUT_AMPL_WIDTH),
		31397 => to_signed(4295, LUT_AMPL_WIDTH),
		31398 => to_signed(4291, LUT_AMPL_WIDTH),
		31399 => to_signed(4288, LUT_AMPL_WIDTH),
		31400 => to_signed(4285, LUT_AMPL_WIDTH),
		31401 => to_signed(4282, LUT_AMPL_WIDTH),
		31402 => to_signed(4279, LUT_AMPL_WIDTH),
		31403 => to_signed(4276, LUT_AMPL_WIDTH),
		31404 => to_signed(4273, LUT_AMPL_WIDTH),
		31405 => to_signed(4270, LUT_AMPL_WIDTH),
		31406 => to_signed(4267, LUT_AMPL_WIDTH),
		31407 => to_signed(4263, LUT_AMPL_WIDTH),
		31408 => to_signed(4260, LUT_AMPL_WIDTH),
		31409 => to_signed(4257, LUT_AMPL_WIDTH),
		31410 => to_signed(4254, LUT_AMPL_WIDTH),
		31411 => to_signed(4251, LUT_AMPL_WIDTH),
		31412 => to_signed(4248, LUT_AMPL_WIDTH),
		31413 => to_signed(4245, LUT_AMPL_WIDTH),
		31414 => to_signed(4242, LUT_AMPL_WIDTH),
		31415 => to_signed(4239, LUT_AMPL_WIDTH),
		31416 => to_signed(4235, LUT_AMPL_WIDTH),
		31417 => to_signed(4232, LUT_AMPL_WIDTH),
		31418 => to_signed(4229, LUT_AMPL_WIDTH),
		31419 => to_signed(4226, LUT_AMPL_WIDTH),
		31420 => to_signed(4223, LUT_AMPL_WIDTH),
		31421 => to_signed(4220, LUT_AMPL_WIDTH),
		31422 => to_signed(4217, LUT_AMPL_WIDTH),
		31423 => to_signed(4214, LUT_AMPL_WIDTH),
		31424 => to_signed(4210, LUT_AMPL_WIDTH),
		31425 => to_signed(4207, LUT_AMPL_WIDTH),
		31426 => to_signed(4204, LUT_AMPL_WIDTH),
		31427 => to_signed(4201, LUT_AMPL_WIDTH),
		31428 => to_signed(4198, LUT_AMPL_WIDTH),
		31429 => to_signed(4195, LUT_AMPL_WIDTH),
		31430 => to_signed(4192, LUT_AMPL_WIDTH),
		31431 => to_signed(4189, LUT_AMPL_WIDTH),
		31432 => to_signed(4186, LUT_AMPL_WIDTH),
		31433 => to_signed(4182, LUT_AMPL_WIDTH),
		31434 => to_signed(4179, LUT_AMPL_WIDTH),
		31435 => to_signed(4176, LUT_AMPL_WIDTH),
		31436 => to_signed(4173, LUT_AMPL_WIDTH),
		31437 => to_signed(4170, LUT_AMPL_WIDTH),
		31438 => to_signed(4167, LUT_AMPL_WIDTH),
		31439 => to_signed(4164, LUT_AMPL_WIDTH),
		31440 => to_signed(4161, LUT_AMPL_WIDTH),
		31441 => to_signed(4158, LUT_AMPL_WIDTH),
		31442 => to_signed(4154, LUT_AMPL_WIDTH),
		31443 => to_signed(4151, LUT_AMPL_WIDTH),
		31444 => to_signed(4148, LUT_AMPL_WIDTH),
		31445 => to_signed(4145, LUT_AMPL_WIDTH),
		31446 => to_signed(4142, LUT_AMPL_WIDTH),
		31447 => to_signed(4139, LUT_AMPL_WIDTH),
		31448 => to_signed(4136, LUT_AMPL_WIDTH),
		31449 => to_signed(4133, LUT_AMPL_WIDTH),
		31450 => to_signed(4129, LUT_AMPL_WIDTH),
		31451 => to_signed(4126, LUT_AMPL_WIDTH),
		31452 => to_signed(4123, LUT_AMPL_WIDTH),
		31453 => to_signed(4120, LUT_AMPL_WIDTH),
		31454 => to_signed(4117, LUT_AMPL_WIDTH),
		31455 => to_signed(4114, LUT_AMPL_WIDTH),
		31456 => to_signed(4111, LUT_AMPL_WIDTH),
		31457 => to_signed(4108, LUT_AMPL_WIDTH),
		31458 => to_signed(4105, LUT_AMPL_WIDTH),
		31459 => to_signed(4101, LUT_AMPL_WIDTH),
		31460 => to_signed(4098, LUT_AMPL_WIDTH),
		31461 => to_signed(4095, LUT_AMPL_WIDTH),
		31462 => to_signed(4092, LUT_AMPL_WIDTH),
		31463 => to_signed(4089, LUT_AMPL_WIDTH),
		31464 => to_signed(4086, LUT_AMPL_WIDTH),
		31465 => to_signed(4083, LUT_AMPL_WIDTH),
		31466 => to_signed(4080, LUT_AMPL_WIDTH),
		31467 => to_signed(4076, LUT_AMPL_WIDTH),
		31468 => to_signed(4073, LUT_AMPL_WIDTH),
		31469 => to_signed(4070, LUT_AMPL_WIDTH),
		31470 => to_signed(4067, LUT_AMPL_WIDTH),
		31471 => to_signed(4064, LUT_AMPL_WIDTH),
		31472 => to_signed(4061, LUT_AMPL_WIDTH),
		31473 => to_signed(4058, LUT_AMPL_WIDTH),
		31474 => to_signed(4055, LUT_AMPL_WIDTH),
		31475 => to_signed(4052, LUT_AMPL_WIDTH),
		31476 => to_signed(4048, LUT_AMPL_WIDTH),
		31477 => to_signed(4045, LUT_AMPL_WIDTH),
		31478 => to_signed(4042, LUT_AMPL_WIDTH),
		31479 => to_signed(4039, LUT_AMPL_WIDTH),
		31480 => to_signed(4036, LUT_AMPL_WIDTH),
		31481 => to_signed(4033, LUT_AMPL_WIDTH),
		31482 => to_signed(4030, LUT_AMPL_WIDTH),
		31483 => to_signed(4027, LUT_AMPL_WIDTH),
		31484 => to_signed(4024, LUT_AMPL_WIDTH),
		31485 => to_signed(4020, LUT_AMPL_WIDTH),
		31486 => to_signed(4017, LUT_AMPL_WIDTH),
		31487 => to_signed(4014, LUT_AMPL_WIDTH),
		31488 => to_signed(4011, LUT_AMPL_WIDTH),
		31489 => to_signed(4008, LUT_AMPL_WIDTH),
		31490 => to_signed(4005, LUT_AMPL_WIDTH),
		31491 => to_signed(4002, LUT_AMPL_WIDTH),
		31492 => to_signed(3999, LUT_AMPL_WIDTH),
		31493 => to_signed(3995, LUT_AMPL_WIDTH),
		31494 => to_signed(3992, LUT_AMPL_WIDTH),
		31495 => to_signed(3989, LUT_AMPL_WIDTH),
		31496 => to_signed(3986, LUT_AMPL_WIDTH),
		31497 => to_signed(3983, LUT_AMPL_WIDTH),
		31498 => to_signed(3980, LUT_AMPL_WIDTH),
		31499 => to_signed(3977, LUT_AMPL_WIDTH),
		31500 => to_signed(3974, LUT_AMPL_WIDTH),
		31501 => to_signed(3970, LUT_AMPL_WIDTH),
		31502 => to_signed(3967, LUT_AMPL_WIDTH),
		31503 => to_signed(3964, LUT_AMPL_WIDTH),
		31504 => to_signed(3961, LUT_AMPL_WIDTH),
		31505 => to_signed(3958, LUT_AMPL_WIDTH),
		31506 => to_signed(3955, LUT_AMPL_WIDTH),
		31507 => to_signed(3952, LUT_AMPL_WIDTH),
		31508 => to_signed(3949, LUT_AMPL_WIDTH),
		31509 => to_signed(3946, LUT_AMPL_WIDTH),
		31510 => to_signed(3942, LUT_AMPL_WIDTH),
		31511 => to_signed(3939, LUT_AMPL_WIDTH),
		31512 => to_signed(3936, LUT_AMPL_WIDTH),
		31513 => to_signed(3933, LUT_AMPL_WIDTH),
		31514 => to_signed(3930, LUT_AMPL_WIDTH),
		31515 => to_signed(3927, LUT_AMPL_WIDTH),
		31516 => to_signed(3924, LUT_AMPL_WIDTH),
		31517 => to_signed(3921, LUT_AMPL_WIDTH),
		31518 => to_signed(3917, LUT_AMPL_WIDTH),
		31519 => to_signed(3914, LUT_AMPL_WIDTH),
		31520 => to_signed(3911, LUT_AMPL_WIDTH),
		31521 => to_signed(3908, LUT_AMPL_WIDTH),
		31522 => to_signed(3905, LUT_AMPL_WIDTH),
		31523 => to_signed(3902, LUT_AMPL_WIDTH),
		31524 => to_signed(3899, LUT_AMPL_WIDTH),
		31525 => to_signed(3896, LUT_AMPL_WIDTH),
		31526 => to_signed(3893, LUT_AMPL_WIDTH),
		31527 => to_signed(3889, LUT_AMPL_WIDTH),
		31528 => to_signed(3886, LUT_AMPL_WIDTH),
		31529 => to_signed(3883, LUT_AMPL_WIDTH),
		31530 => to_signed(3880, LUT_AMPL_WIDTH),
		31531 => to_signed(3877, LUT_AMPL_WIDTH),
		31532 => to_signed(3874, LUT_AMPL_WIDTH),
		31533 => to_signed(3871, LUT_AMPL_WIDTH),
		31534 => to_signed(3868, LUT_AMPL_WIDTH),
		31535 => to_signed(3864, LUT_AMPL_WIDTH),
		31536 => to_signed(3861, LUT_AMPL_WIDTH),
		31537 => to_signed(3858, LUT_AMPL_WIDTH),
		31538 => to_signed(3855, LUT_AMPL_WIDTH),
		31539 => to_signed(3852, LUT_AMPL_WIDTH),
		31540 => to_signed(3849, LUT_AMPL_WIDTH),
		31541 => to_signed(3846, LUT_AMPL_WIDTH),
		31542 => to_signed(3843, LUT_AMPL_WIDTH),
		31543 => to_signed(3839, LUT_AMPL_WIDTH),
		31544 => to_signed(3836, LUT_AMPL_WIDTH),
		31545 => to_signed(3833, LUT_AMPL_WIDTH),
		31546 => to_signed(3830, LUT_AMPL_WIDTH),
		31547 => to_signed(3827, LUT_AMPL_WIDTH),
		31548 => to_signed(3824, LUT_AMPL_WIDTH),
		31549 => to_signed(3821, LUT_AMPL_WIDTH),
		31550 => to_signed(3818, LUT_AMPL_WIDTH),
		31551 => to_signed(3815, LUT_AMPL_WIDTH),
		31552 => to_signed(3811, LUT_AMPL_WIDTH),
		31553 => to_signed(3808, LUT_AMPL_WIDTH),
		31554 => to_signed(3805, LUT_AMPL_WIDTH),
		31555 => to_signed(3802, LUT_AMPL_WIDTH),
		31556 => to_signed(3799, LUT_AMPL_WIDTH),
		31557 => to_signed(3796, LUT_AMPL_WIDTH),
		31558 => to_signed(3793, LUT_AMPL_WIDTH),
		31559 => to_signed(3790, LUT_AMPL_WIDTH),
		31560 => to_signed(3786, LUT_AMPL_WIDTH),
		31561 => to_signed(3783, LUT_AMPL_WIDTH),
		31562 => to_signed(3780, LUT_AMPL_WIDTH),
		31563 => to_signed(3777, LUT_AMPL_WIDTH),
		31564 => to_signed(3774, LUT_AMPL_WIDTH),
		31565 => to_signed(3771, LUT_AMPL_WIDTH),
		31566 => to_signed(3768, LUT_AMPL_WIDTH),
		31567 => to_signed(3765, LUT_AMPL_WIDTH),
		31568 => to_signed(3761, LUT_AMPL_WIDTH),
		31569 => to_signed(3758, LUT_AMPL_WIDTH),
		31570 => to_signed(3755, LUT_AMPL_WIDTH),
		31571 => to_signed(3752, LUT_AMPL_WIDTH),
		31572 => to_signed(3749, LUT_AMPL_WIDTH),
		31573 => to_signed(3746, LUT_AMPL_WIDTH),
		31574 => to_signed(3743, LUT_AMPL_WIDTH),
		31575 => to_signed(3740, LUT_AMPL_WIDTH),
		31576 => to_signed(3737, LUT_AMPL_WIDTH),
		31577 => to_signed(3733, LUT_AMPL_WIDTH),
		31578 => to_signed(3730, LUT_AMPL_WIDTH),
		31579 => to_signed(3727, LUT_AMPL_WIDTH),
		31580 => to_signed(3724, LUT_AMPL_WIDTH),
		31581 => to_signed(3721, LUT_AMPL_WIDTH),
		31582 => to_signed(3718, LUT_AMPL_WIDTH),
		31583 => to_signed(3715, LUT_AMPL_WIDTH),
		31584 => to_signed(3712, LUT_AMPL_WIDTH),
		31585 => to_signed(3708, LUT_AMPL_WIDTH),
		31586 => to_signed(3705, LUT_AMPL_WIDTH),
		31587 => to_signed(3702, LUT_AMPL_WIDTH),
		31588 => to_signed(3699, LUT_AMPL_WIDTH),
		31589 => to_signed(3696, LUT_AMPL_WIDTH),
		31590 => to_signed(3693, LUT_AMPL_WIDTH),
		31591 => to_signed(3690, LUT_AMPL_WIDTH),
		31592 => to_signed(3687, LUT_AMPL_WIDTH),
		31593 => to_signed(3683, LUT_AMPL_WIDTH),
		31594 => to_signed(3680, LUT_AMPL_WIDTH),
		31595 => to_signed(3677, LUT_AMPL_WIDTH),
		31596 => to_signed(3674, LUT_AMPL_WIDTH),
		31597 => to_signed(3671, LUT_AMPL_WIDTH),
		31598 => to_signed(3668, LUT_AMPL_WIDTH),
		31599 => to_signed(3665, LUT_AMPL_WIDTH),
		31600 => to_signed(3662, LUT_AMPL_WIDTH),
		31601 => to_signed(3658, LUT_AMPL_WIDTH),
		31602 => to_signed(3655, LUT_AMPL_WIDTH),
		31603 => to_signed(3652, LUT_AMPL_WIDTH),
		31604 => to_signed(3649, LUT_AMPL_WIDTH),
		31605 => to_signed(3646, LUT_AMPL_WIDTH),
		31606 => to_signed(3643, LUT_AMPL_WIDTH),
		31607 => to_signed(3640, LUT_AMPL_WIDTH),
		31608 => to_signed(3637, LUT_AMPL_WIDTH),
		31609 => to_signed(3634, LUT_AMPL_WIDTH),
		31610 => to_signed(3630, LUT_AMPL_WIDTH),
		31611 => to_signed(3627, LUT_AMPL_WIDTH),
		31612 => to_signed(3624, LUT_AMPL_WIDTH),
		31613 => to_signed(3621, LUT_AMPL_WIDTH),
		31614 => to_signed(3618, LUT_AMPL_WIDTH),
		31615 => to_signed(3615, LUT_AMPL_WIDTH),
		31616 => to_signed(3612, LUT_AMPL_WIDTH),
		31617 => to_signed(3609, LUT_AMPL_WIDTH),
		31618 => to_signed(3605, LUT_AMPL_WIDTH),
		31619 => to_signed(3602, LUT_AMPL_WIDTH),
		31620 => to_signed(3599, LUT_AMPL_WIDTH),
		31621 => to_signed(3596, LUT_AMPL_WIDTH),
		31622 => to_signed(3593, LUT_AMPL_WIDTH),
		31623 => to_signed(3590, LUT_AMPL_WIDTH),
		31624 => to_signed(3587, LUT_AMPL_WIDTH),
		31625 => to_signed(3584, LUT_AMPL_WIDTH),
		31626 => to_signed(3580, LUT_AMPL_WIDTH),
		31627 => to_signed(3577, LUT_AMPL_WIDTH),
		31628 => to_signed(3574, LUT_AMPL_WIDTH),
		31629 => to_signed(3571, LUT_AMPL_WIDTH),
		31630 => to_signed(3568, LUT_AMPL_WIDTH),
		31631 => to_signed(3565, LUT_AMPL_WIDTH),
		31632 => to_signed(3562, LUT_AMPL_WIDTH),
		31633 => to_signed(3559, LUT_AMPL_WIDTH),
		31634 => to_signed(3555, LUT_AMPL_WIDTH),
		31635 => to_signed(3552, LUT_AMPL_WIDTH),
		31636 => to_signed(3549, LUT_AMPL_WIDTH),
		31637 => to_signed(3546, LUT_AMPL_WIDTH),
		31638 => to_signed(3543, LUT_AMPL_WIDTH),
		31639 => to_signed(3540, LUT_AMPL_WIDTH),
		31640 => to_signed(3537, LUT_AMPL_WIDTH),
		31641 => to_signed(3534, LUT_AMPL_WIDTH),
		31642 => to_signed(3530, LUT_AMPL_WIDTH),
		31643 => to_signed(3527, LUT_AMPL_WIDTH),
		31644 => to_signed(3524, LUT_AMPL_WIDTH),
		31645 => to_signed(3521, LUT_AMPL_WIDTH),
		31646 => to_signed(3518, LUT_AMPL_WIDTH),
		31647 => to_signed(3515, LUT_AMPL_WIDTH),
		31648 => to_signed(3512, LUT_AMPL_WIDTH),
		31649 => to_signed(3509, LUT_AMPL_WIDTH),
		31650 => to_signed(3505, LUT_AMPL_WIDTH),
		31651 => to_signed(3502, LUT_AMPL_WIDTH),
		31652 => to_signed(3499, LUT_AMPL_WIDTH),
		31653 => to_signed(3496, LUT_AMPL_WIDTH),
		31654 => to_signed(3493, LUT_AMPL_WIDTH),
		31655 => to_signed(3490, LUT_AMPL_WIDTH),
		31656 => to_signed(3487, LUT_AMPL_WIDTH),
		31657 => to_signed(3484, LUT_AMPL_WIDTH),
		31658 => to_signed(3480, LUT_AMPL_WIDTH),
		31659 => to_signed(3477, LUT_AMPL_WIDTH),
		31660 => to_signed(3474, LUT_AMPL_WIDTH),
		31661 => to_signed(3471, LUT_AMPL_WIDTH),
		31662 => to_signed(3468, LUT_AMPL_WIDTH),
		31663 => to_signed(3465, LUT_AMPL_WIDTH),
		31664 => to_signed(3462, LUT_AMPL_WIDTH),
		31665 => to_signed(3459, LUT_AMPL_WIDTH),
		31666 => to_signed(3455, LUT_AMPL_WIDTH),
		31667 => to_signed(3452, LUT_AMPL_WIDTH),
		31668 => to_signed(3449, LUT_AMPL_WIDTH),
		31669 => to_signed(3446, LUT_AMPL_WIDTH),
		31670 => to_signed(3443, LUT_AMPL_WIDTH),
		31671 => to_signed(3440, LUT_AMPL_WIDTH),
		31672 => to_signed(3437, LUT_AMPL_WIDTH),
		31673 => to_signed(3434, LUT_AMPL_WIDTH),
		31674 => to_signed(3430, LUT_AMPL_WIDTH),
		31675 => to_signed(3427, LUT_AMPL_WIDTH),
		31676 => to_signed(3424, LUT_AMPL_WIDTH),
		31677 => to_signed(3421, LUT_AMPL_WIDTH),
		31678 => to_signed(3418, LUT_AMPL_WIDTH),
		31679 => to_signed(3415, LUT_AMPL_WIDTH),
		31680 => to_signed(3412, LUT_AMPL_WIDTH),
		31681 => to_signed(3409, LUT_AMPL_WIDTH),
		31682 => to_signed(3406, LUT_AMPL_WIDTH),
		31683 => to_signed(3402, LUT_AMPL_WIDTH),
		31684 => to_signed(3399, LUT_AMPL_WIDTH),
		31685 => to_signed(3396, LUT_AMPL_WIDTH),
		31686 => to_signed(3393, LUT_AMPL_WIDTH),
		31687 => to_signed(3390, LUT_AMPL_WIDTH),
		31688 => to_signed(3387, LUT_AMPL_WIDTH),
		31689 => to_signed(3384, LUT_AMPL_WIDTH),
		31690 => to_signed(3381, LUT_AMPL_WIDTH),
		31691 => to_signed(3377, LUT_AMPL_WIDTH),
		31692 => to_signed(3374, LUT_AMPL_WIDTH),
		31693 => to_signed(3371, LUT_AMPL_WIDTH),
		31694 => to_signed(3368, LUT_AMPL_WIDTH),
		31695 => to_signed(3365, LUT_AMPL_WIDTH),
		31696 => to_signed(3362, LUT_AMPL_WIDTH),
		31697 => to_signed(3359, LUT_AMPL_WIDTH),
		31698 => to_signed(3356, LUT_AMPL_WIDTH),
		31699 => to_signed(3352, LUT_AMPL_WIDTH),
		31700 => to_signed(3349, LUT_AMPL_WIDTH),
		31701 => to_signed(3346, LUT_AMPL_WIDTH),
		31702 => to_signed(3343, LUT_AMPL_WIDTH),
		31703 => to_signed(3340, LUT_AMPL_WIDTH),
		31704 => to_signed(3337, LUT_AMPL_WIDTH),
		31705 => to_signed(3334, LUT_AMPL_WIDTH),
		31706 => to_signed(3331, LUT_AMPL_WIDTH),
		31707 => to_signed(3327, LUT_AMPL_WIDTH),
		31708 => to_signed(3324, LUT_AMPL_WIDTH),
		31709 => to_signed(3321, LUT_AMPL_WIDTH),
		31710 => to_signed(3318, LUT_AMPL_WIDTH),
		31711 => to_signed(3315, LUT_AMPL_WIDTH),
		31712 => to_signed(3312, LUT_AMPL_WIDTH),
		31713 => to_signed(3309, LUT_AMPL_WIDTH),
		31714 => to_signed(3306, LUT_AMPL_WIDTH),
		31715 => to_signed(3302, LUT_AMPL_WIDTH),
		31716 => to_signed(3299, LUT_AMPL_WIDTH),
		31717 => to_signed(3296, LUT_AMPL_WIDTH),
		31718 => to_signed(3293, LUT_AMPL_WIDTH),
		31719 => to_signed(3290, LUT_AMPL_WIDTH),
		31720 => to_signed(3287, LUT_AMPL_WIDTH),
		31721 => to_signed(3284, LUT_AMPL_WIDTH),
		31722 => to_signed(3281, LUT_AMPL_WIDTH),
		31723 => to_signed(3277, LUT_AMPL_WIDTH),
		31724 => to_signed(3274, LUT_AMPL_WIDTH),
		31725 => to_signed(3271, LUT_AMPL_WIDTH),
		31726 => to_signed(3268, LUT_AMPL_WIDTH),
		31727 => to_signed(3265, LUT_AMPL_WIDTH),
		31728 => to_signed(3262, LUT_AMPL_WIDTH),
		31729 => to_signed(3259, LUT_AMPL_WIDTH),
		31730 => to_signed(3255, LUT_AMPL_WIDTH),
		31731 => to_signed(3252, LUT_AMPL_WIDTH),
		31732 => to_signed(3249, LUT_AMPL_WIDTH),
		31733 => to_signed(3246, LUT_AMPL_WIDTH),
		31734 => to_signed(3243, LUT_AMPL_WIDTH),
		31735 => to_signed(3240, LUT_AMPL_WIDTH),
		31736 => to_signed(3237, LUT_AMPL_WIDTH),
		31737 => to_signed(3234, LUT_AMPL_WIDTH),
		31738 => to_signed(3230, LUT_AMPL_WIDTH),
		31739 => to_signed(3227, LUT_AMPL_WIDTH),
		31740 => to_signed(3224, LUT_AMPL_WIDTH),
		31741 => to_signed(3221, LUT_AMPL_WIDTH),
		31742 => to_signed(3218, LUT_AMPL_WIDTH),
		31743 => to_signed(3215, LUT_AMPL_WIDTH),
		31744 => to_signed(3212, LUT_AMPL_WIDTH),
		31745 => to_signed(3209, LUT_AMPL_WIDTH),
		31746 => to_signed(3205, LUT_AMPL_WIDTH),
		31747 => to_signed(3202, LUT_AMPL_WIDTH),
		31748 => to_signed(3199, LUT_AMPL_WIDTH),
		31749 => to_signed(3196, LUT_AMPL_WIDTH),
		31750 => to_signed(3193, LUT_AMPL_WIDTH),
		31751 => to_signed(3190, LUT_AMPL_WIDTH),
		31752 => to_signed(3187, LUT_AMPL_WIDTH),
		31753 => to_signed(3184, LUT_AMPL_WIDTH),
		31754 => to_signed(3180, LUT_AMPL_WIDTH),
		31755 => to_signed(3177, LUT_AMPL_WIDTH),
		31756 => to_signed(3174, LUT_AMPL_WIDTH),
		31757 => to_signed(3171, LUT_AMPL_WIDTH),
		31758 => to_signed(3168, LUT_AMPL_WIDTH),
		31759 => to_signed(3165, LUT_AMPL_WIDTH),
		31760 => to_signed(3162, LUT_AMPL_WIDTH),
		31761 => to_signed(3159, LUT_AMPL_WIDTH),
		31762 => to_signed(3155, LUT_AMPL_WIDTH),
		31763 => to_signed(3152, LUT_AMPL_WIDTH),
		31764 => to_signed(3149, LUT_AMPL_WIDTH),
		31765 => to_signed(3146, LUT_AMPL_WIDTH),
		31766 => to_signed(3143, LUT_AMPL_WIDTH),
		31767 => to_signed(3140, LUT_AMPL_WIDTH),
		31768 => to_signed(3137, LUT_AMPL_WIDTH),
		31769 => to_signed(3134, LUT_AMPL_WIDTH),
		31770 => to_signed(3130, LUT_AMPL_WIDTH),
		31771 => to_signed(3127, LUT_AMPL_WIDTH),
		31772 => to_signed(3124, LUT_AMPL_WIDTH),
		31773 => to_signed(3121, LUT_AMPL_WIDTH),
		31774 => to_signed(3118, LUT_AMPL_WIDTH),
		31775 => to_signed(3115, LUT_AMPL_WIDTH),
		31776 => to_signed(3112, LUT_AMPL_WIDTH),
		31777 => to_signed(3109, LUT_AMPL_WIDTH),
		31778 => to_signed(3105, LUT_AMPL_WIDTH),
		31779 => to_signed(3102, LUT_AMPL_WIDTH),
		31780 => to_signed(3099, LUT_AMPL_WIDTH),
		31781 => to_signed(3096, LUT_AMPL_WIDTH),
		31782 => to_signed(3093, LUT_AMPL_WIDTH),
		31783 => to_signed(3090, LUT_AMPL_WIDTH),
		31784 => to_signed(3087, LUT_AMPL_WIDTH),
		31785 => to_signed(3084, LUT_AMPL_WIDTH),
		31786 => to_signed(3080, LUT_AMPL_WIDTH),
		31787 => to_signed(3077, LUT_AMPL_WIDTH),
		31788 => to_signed(3074, LUT_AMPL_WIDTH),
		31789 => to_signed(3071, LUT_AMPL_WIDTH),
		31790 => to_signed(3068, LUT_AMPL_WIDTH),
		31791 => to_signed(3065, LUT_AMPL_WIDTH),
		31792 => to_signed(3062, LUT_AMPL_WIDTH),
		31793 => to_signed(3059, LUT_AMPL_WIDTH),
		31794 => to_signed(3055, LUT_AMPL_WIDTH),
		31795 => to_signed(3052, LUT_AMPL_WIDTH),
		31796 => to_signed(3049, LUT_AMPL_WIDTH),
		31797 => to_signed(3046, LUT_AMPL_WIDTH),
		31798 => to_signed(3043, LUT_AMPL_WIDTH),
		31799 => to_signed(3040, LUT_AMPL_WIDTH),
		31800 => to_signed(3037, LUT_AMPL_WIDTH),
		31801 => to_signed(3033, LUT_AMPL_WIDTH),
		31802 => to_signed(3030, LUT_AMPL_WIDTH),
		31803 => to_signed(3027, LUT_AMPL_WIDTH),
		31804 => to_signed(3024, LUT_AMPL_WIDTH),
		31805 => to_signed(3021, LUT_AMPL_WIDTH),
		31806 => to_signed(3018, LUT_AMPL_WIDTH),
		31807 => to_signed(3015, LUT_AMPL_WIDTH),
		31808 => to_signed(3012, LUT_AMPL_WIDTH),
		31809 => to_signed(3008, LUT_AMPL_WIDTH),
		31810 => to_signed(3005, LUT_AMPL_WIDTH),
		31811 => to_signed(3002, LUT_AMPL_WIDTH),
		31812 => to_signed(2999, LUT_AMPL_WIDTH),
		31813 => to_signed(2996, LUT_AMPL_WIDTH),
		31814 => to_signed(2993, LUT_AMPL_WIDTH),
		31815 => to_signed(2990, LUT_AMPL_WIDTH),
		31816 => to_signed(2987, LUT_AMPL_WIDTH),
		31817 => to_signed(2983, LUT_AMPL_WIDTH),
		31818 => to_signed(2980, LUT_AMPL_WIDTH),
		31819 => to_signed(2977, LUT_AMPL_WIDTH),
		31820 => to_signed(2974, LUT_AMPL_WIDTH),
		31821 => to_signed(2971, LUT_AMPL_WIDTH),
		31822 => to_signed(2968, LUT_AMPL_WIDTH),
		31823 => to_signed(2965, LUT_AMPL_WIDTH),
		31824 => to_signed(2962, LUT_AMPL_WIDTH),
		31825 => to_signed(2958, LUT_AMPL_WIDTH),
		31826 => to_signed(2955, LUT_AMPL_WIDTH),
		31827 => to_signed(2952, LUT_AMPL_WIDTH),
		31828 => to_signed(2949, LUT_AMPL_WIDTH),
		31829 => to_signed(2946, LUT_AMPL_WIDTH),
		31830 => to_signed(2943, LUT_AMPL_WIDTH),
		31831 => to_signed(2940, LUT_AMPL_WIDTH),
		31832 => to_signed(2936, LUT_AMPL_WIDTH),
		31833 => to_signed(2933, LUT_AMPL_WIDTH),
		31834 => to_signed(2930, LUT_AMPL_WIDTH),
		31835 => to_signed(2927, LUT_AMPL_WIDTH),
		31836 => to_signed(2924, LUT_AMPL_WIDTH),
		31837 => to_signed(2921, LUT_AMPL_WIDTH),
		31838 => to_signed(2918, LUT_AMPL_WIDTH),
		31839 => to_signed(2915, LUT_AMPL_WIDTH),
		31840 => to_signed(2911, LUT_AMPL_WIDTH),
		31841 => to_signed(2908, LUT_AMPL_WIDTH),
		31842 => to_signed(2905, LUT_AMPL_WIDTH),
		31843 => to_signed(2902, LUT_AMPL_WIDTH),
		31844 => to_signed(2899, LUT_AMPL_WIDTH),
		31845 => to_signed(2896, LUT_AMPL_WIDTH),
		31846 => to_signed(2893, LUT_AMPL_WIDTH),
		31847 => to_signed(2890, LUT_AMPL_WIDTH),
		31848 => to_signed(2886, LUT_AMPL_WIDTH),
		31849 => to_signed(2883, LUT_AMPL_WIDTH),
		31850 => to_signed(2880, LUT_AMPL_WIDTH),
		31851 => to_signed(2877, LUT_AMPL_WIDTH),
		31852 => to_signed(2874, LUT_AMPL_WIDTH),
		31853 => to_signed(2871, LUT_AMPL_WIDTH),
		31854 => to_signed(2868, LUT_AMPL_WIDTH),
		31855 => to_signed(2865, LUT_AMPL_WIDTH),
		31856 => to_signed(2861, LUT_AMPL_WIDTH),
		31857 => to_signed(2858, LUT_AMPL_WIDTH),
		31858 => to_signed(2855, LUT_AMPL_WIDTH),
		31859 => to_signed(2852, LUT_AMPL_WIDTH),
		31860 => to_signed(2849, LUT_AMPL_WIDTH),
		31861 => to_signed(2846, LUT_AMPL_WIDTH),
		31862 => to_signed(2843, LUT_AMPL_WIDTH),
		31863 => to_signed(2839, LUT_AMPL_WIDTH),
		31864 => to_signed(2836, LUT_AMPL_WIDTH),
		31865 => to_signed(2833, LUT_AMPL_WIDTH),
		31866 => to_signed(2830, LUT_AMPL_WIDTH),
		31867 => to_signed(2827, LUT_AMPL_WIDTH),
		31868 => to_signed(2824, LUT_AMPL_WIDTH),
		31869 => to_signed(2821, LUT_AMPL_WIDTH),
		31870 => to_signed(2818, LUT_AMPL_WIDTH),
		31871 => to_signed(2814, LUT_AMPL_WIDTH),
		31872 => to_signed(2811, LUT_AMPL_WIDTH),
		31873 => to_signed(2808, LUT_AMPL_WIDTH),
		31874 => to_signed(2805, LUT_AMPL_WIDTH),
		31875 => to_signed(2802, LUT_AMPL_WIDTH),
		31876 => to_signed(2799, LUT_AMPL_WIDTH),
		31877 => to_signed(2796, LUT_AMPL_WIDTH),
		31878 => to_signed(2793, LUT_AMPL_WIDTH),
		31879 => to_signed(2789, LUT_AMPL_WIDTH),
		31880 => to_signed(2786, LUT_AMPL_WIDTH),
		31881 => to_signed(2783, LUT_AMPL_WIDTH),
		31882 => to_signed(2780, LUT_AMPL_WIDTH),
		31883 => to_signed(2777, LUT_AMPL_WIDTH),
		31884 => to_signed(2774, LUT_AMPL_WIDTH),
		31885 => to_signed(2771, LUT_AMPL_WIDTH),
		31886 => to_signed(2767, LUT_AMPL_WIDTH),
		31887 => to_signed(2764, LUT_AMPL_WIDTH),
		31888 => to_signed(2761, LUT_AMPL_WIDTH),
		31889 => to_signed(2758, LUT_AMPL_WIDTH),
		31890 => to_signed(2755, LUT_AMPL_WIDTH),
		31891 => to_signed(2752, LUT_AMPL_WIDTH),
		31892 => to_signed(2749, LUT_AMPL_WIDTH),
		31893 => to_signed(2746, LUT_AMPL_WIDTH),
		31894 => to_signed(2742, LUT_AMPL_WIDTH),
		31895 => to_signed(2739, LUT_AMPL_WIDTH),
		31896 => to_signed(2736, LUT_AMPL_WIDTH),
		31897 => to_signed(2733, LUT_AMPL_WIDTH),
		31898 => to_signed(2730, LUT_AMPL_WIDTH),
		31899 => to_signed(2727, LUT_AMPL_WIDTH),
		31900 => to_signed(2724, LUT_AMPL_WIDTH),
		31901 => to_signed(2721, LUT_AMPL_WIDTH),
		31902 => to_signed(2717, LUT_AMPL_WIDTH),
		31903 => to_signed(2714, LUT_AMPL_WIDTH),
		31904 => to_signed(2711, LUT_AMPL_WIDTH),
		31905 => to_signed(2708, LUT_AMPL_WIDTH),
		31906 => to_signed(2705, LUT_AMPL_WIDTH),
		31907 => to_signed(2702, LUT_AMPL_WIDTH),
		31908 => to_signed(2699, LUT_AMPL_WIDTH),
		31909 => to_signed(2695, LUT_AMPL_WIDTH),
		31910 => to_signed(2692, LUT_AMPL_WIDTH),
		31911 => to_signed(2689, LUT_AMPL_WIDTH),
		31912 => to_signed(2686, LUT_AMPL_WIDTH),
		31913 => to_signed(2683, LUT_AMPL_WIDTH),
		31914 => to_signed(2680, LUT_AMPL_WIDTH),
		31915 => to_signed(2677, LUT_AMPL_WIDTH),
		31916 => to_signed(2674, LUT_AMPL_WIDTH),
		31917 => to_signed(2670, LUT_AMPL_WIDTH),
		31918 => to_signed(2667, LUT_AMPL_WIDTH),
		31919 => to_signed(2664, LUT_AMPL_WIDTH),
		31920 => to_signed(2661, LUT_AMPL_WIDTH),
		31921 => to_signed(2658, LUT_AMPL_WIDTH),
		31922 => to_signed(2655, LUT_AMPL_WIDTH),
		31923 => to_signed(2652, LUT_AMPL_WIDTH),
		31924 => to_signed(2649, LUT_AMPL_WIDTH),
		31925 => to_signed(2645, LUT_AMPL_WIDTH),
		31926 => to_signed(2642, LUT_AMPL_WIDTH),
		31927 => to_signed(2639, LUT_AMPL_WIDTH),
		31928 => to_signed(2636, LUT_AMPL_WIDTH),
		31929 => to_signed(2633, LUT_AMPL_WIDTH),
		31930 => to_signed(2630, LUT_AMPL_WIDTH),
		31931 => to_signed(2627, LUT_AMPL_WIDTH),
		31932 => to_signed(2623, LUT_AMPL_WIDTH),
		31933 => to_signed(2620, LUT_AMPL_WIDTH),
		31934 => to_signed(2617, LUT_AMPL_WIDTH),
		31935 => to_signed(2614, LUT_AMPL_WIDTH),
		31936 => to_signed(2611, LUT_AMPL_WIDTH),
		31937 => to_signed(2608, LUT_AMPL_WIDTH),
		31938 => to_signed(2605, LUT_AMPL_WIDTH),
		31939 => to_signed(2602, LUT_AMPL_WIDTH),
		31940 => to_signed(2598, LUT_AMPL_WIDTH),
		31941 => to_signed(2595, LUT_AMPL_WIDTH),
		31942 => to_signed(2592, LUT_AMPL_WIDTH),
		31943 => to_signed(2589, LUT_AMPL_WIDTH),
		31944 => to_signed(2586, LUT_AMPL_WIDTH),
		31945 => to_signed(2583, LUT_AMPL_WIDTH),
		31946 => to_signed(2580, LUT_AMPL_WIDTH),
		31947 => to_signed(2577, LUT_AMPL_WIDTH),
		31948 => to_signed(2573, LUT_AMPL_WIDTH),
		31949 => to_signed(2570, LUT_AMPL_WIDTH),
		31950 => to_signed(2567, LUT_AMPL_WIDTH),
		31951 => to_signed(2564, LUT_AMPL_WIDTH),
		31952 => to_signed(2561, LUT_AMPL_WIDTH),
		31953 => to_signed(2558, LUT_AMPL_WIDTH),
		31954 => to_signed(2555, LUT_AMPL_WIDTH),
		31955 => to_signed(2551, LUT_AMPL_WIDTH),
		31956 => to_signed(2548, LUT_AMPL_WIDTH),
		31957 => to_signed(2545, LUT_AMPL_WIDTH),
		31958 => to_signed(2542, LUT_AMPL_WIDTH),
		31959 => to_signed(2539, LUT_AMPL_WIDTH),
		31960 => to_signed(2536, LUT_AMPL_WIDTH),
		31961 => to_signed(2533, LUT_AMPL_WIDTH),
		31962 => to_signed(2530, LUT_AMPL_WIDTH),
		31963 => to_signed(2526, LUT_AMPL_WIDTH),
		31964 => to_signed(2523, LUT_AMPL_WIDTH),
		31965 => to_signed(2520, LUT_AMPL_WIDTH),
		31966 => to_signed(2517, LUT_AMPL_WIDTH),
		31967 => to_signed(2514, LUT_AMPL_WIDTH),
		31968 => to_signed(2511, LUT_AMPL_WIDTH),
		31969 => to_signed(2508, LUT_AMPL_WIDTH),
		31970 => to_signed(2504, LUT_AMPL_WIDTH),
		31971 => to_signed(2501, LUT_AMPL_WIDTH),
		31972 => to_signed(2498, LUT_AMPL_WIDTH),
		31973 => to_signed(2495, LUT_AMPL_WIDTH),
		31974 => to_signed(2492, LUT_AMPL_WIDTH),
		31975 => to_signed(2489, LUT_AMPL_WIDTH),
		31976 => to_signed(2486, LUT_AMPL_WIDTH),
		31977 => to_signed(2483, LUT_AMPL_WIDTH),
		31978 => to_signed(2479, LUT_AMPL_WIDTH),
		31979 => to_signed(2476, LUT_AMPL_WIDTH),
		31980 => to_signed(2473, LUT_AMPL_WIDTH),
		31981 => to_signed(2470, LUT_AMPL_WIDTH),
		31982 => to_signed(2467, LUT_AMPL_WIDTH),
		31983 => to_signed(2464, LUT_AMPL_WIDTH),
		31984 => to_signed(2461, LUT_AMPL_WIDTH),
		31985 => to_signed(2457, LUT_AMPL_WIDTH),
		31986 => to_signed(2454, LUT_AMPL_WIDTH),
		31987 => to_signed(2451, LUT_AMPL_WIDTH),
		31988 => to_signed(2448, LUT_AMPL_WIDTH),
		31989 => to_signed(2445, LUT_AMPL_WIDTH),
		31990 => to_signed(2442, LUT_AMPL_WIDTH),
		31991 => to_signed(2439, LUT_AMPL_WIDTH),
		31992 => to_signed(2436, LUT_AMPL_WIDTH),
		31993 => to_signed(2432, LUT_AMPL_WIDTH),
		31994 => to_signed(2429, LUT_AMPL_WIDTH),
		31995 => to_signed(2426, LUT_AMPL_WIDTH),
		31996 => to_signed(2423, LUT_AMPL_WIDTH),
		31997 => to_signed(2420, LUT_AMPL_WIDTH),
		31998 => to_signed(2417, LUT_AMPL_WIDTH),
		31999 => to_signed(2414, LUT_AMPL_WIDTH),
		32000 => to_signed(2410, LUT_AMPL_WIDTH),
		32001 => to_signed(2407, LUT_AMPL_WIDTH),
		32002 => to_signed(2404, LUT_AMPL_WIDTH),
		32003 => to_signed(2401, LUT_AMPL_WIDTH),
		32004 => to_signed(2398, LUT_AMPL_WIDTH),
		32005 => to_signed(2395, LUT_AMPL_WIDTH),
		32006 => to_signed(2392, LUT_AMPL_WIDTH),
		32007 => to_signed(2389, LUT_AMPL_WIDTH),
		32008 => to_signed(2385, LUT_AMPL_WIDTH),
		32009 => to_signed(2382, LUT_AMPL_WIDTH),
		32010 => to_signed(2379, LUT_AMPL_WIDTH),
		32011 => to_signed(2376, LUT_AMPL_WIDTH),
		32012 => to_signed(2373, LUT_AMPL_WIDTH),
		32013 => to_signed(2370, LUT_AMPL_WIDTH),
		32014 => to_signed(2367, LUT_AMPL_WIDTH),
		32015 => to_signed(2363, LUT_AMPL_WIDTH),
		32016 => to_signed(2360, LUT_AMPL_WIDTH),
		32017 => to_signed(2357, LUT_AMPL_WIDTH),
		32018 => to_signed(2354, LUT_AMPL_WIDTH),
		32019 => to_signed(2351, LUT_AMPL_WIDTH),
		32020 => to_signed(2348, LUT_AMPL_WIDTH),
		32021 => to_signed(2345, LUT_AMPL_WIDTH),
		32022 => to_signed(2342, LUT_AMPL_WIDTH),
		32023 => to_signed(2338, LUT_AMPL_WIDTH),
		32024 => to_signed(2335, LUT_AMPL_WIDTH),
		32025 => to_signed(2332, LUT_AMPL_WIDTH),
		32026 => to_signed(2329, LUT_AMPL_WIDTH),
		32027 => to_signed(2326, LUT_AMPL_WIDTH),
		32028 => to_signed(2323, LUT_AMPL_WIDTH),
		32029 => to_signed(2320, LUT_AMPL_WIDTH),
		32030 => to_signed(2316, LUT_AMPL_WIDTH),
		32031 => to_signed(2313, LUT_AMPL_WIDTH),
		32032 => to_signed(2310, LUT_AMPL_WIDTH),
		32033 => to_signed(2307, LUT_AMPL_WIDTH),
		32034 => to_signed(2304, LUT_AMPL_WIDTH),
		32035 => to_signed(2301, LUT_AMPL_WIDTH),
		32036 => to_signed(2298, LUT_AMPL_WIDTH),
		32037 => to_signed(2295, LUT_AMPL_WIDTH),
		32038 => to_signed(2291, LUT_AMPL_WIDTH),
		32039 => to_signed(2288, LUT_AMPL_WIDTH),
		32040 => to_signed(2285, LUT_AMPL_WIDTH),
		32041 => to_signed(2282, LUT_AMPL_WIDTH),
		32042 => to_signed(2279, LUT_AMPL_WIDTH),
		32043 => to_signed(2276, LUT_AMPL_WIDTH),
		32044 => to_signed(2273, LUT_AMPL_WIDTH),
		32045 => to_signed(2269, LUT_AMPL_WIDTH),
		32046 => to_signed(2266, LUT_AMPL_WIDTH),
		32047 => to_signed(2263, LUT_AMPL_WIDTH),
		32048 => to_signed(2260, LUT_AMPL_WIDTH),
		32049 => to_signed(2257, LUT_AMPL_WIDTH),
		32050 => to_signed(2254, LUT_AMPL_WIDTH),
		32051 => to_signed(2251, LUT_AMPL_WIDTH),
		32052 => to_signed(2248, LUT_AMPL_WIDTH),
		32053 => to_signed(2244, LUT_AMPL_WIDTH),
		32054 => to_signed(2241, LUT_AMPL_WIDTH),
		32055 => to_signed(2238, LUT_AMPL_WIDTH),
		32056 => to_signed(2235, LUT_AMPL_WIDTH),
		32057 => to_signed(2232, LUT_AMPL_WIDTH),
		32058 => to_signed(2229, LUT_AMPL_WIDTH),
		32059 => to_signed(2226, LUT_AMPL_WIDTH),
		32060 => to_signed(2222, LUT_AMPL_WIDTH),
		32061 => to_signed(2219, LUT_AMPL_WIDTH),
		32062 => to_signed(2216, LUT_AMPL_WIDTH),
		32063 => to_signed(2213, LUT_AMPL_WIDTH),
		32064 => to_signed(2210, LUT_AMPL_WIDTH),
		32065 => to_signed(2207, LUT_AMPL_WIDTH),
		32066 => to_signed(2204, LUT_AMPL_WIDTH),
		32067 => to_signed(2201, LUT_AMPL_WIDTH),
		32068 => to_signed(2197, LUT_AMPL_WIDTH),
		32069 => to_signed(2194, LUT_AMPL_WIDTH),
		32070 => to_signed(2191, LUT_AMPL_WIDTH),
		32071 => to_signed(2188, LUT_AMPL_WIDTH),
		32072 => to_signed(2185, LUT_AMPL_WIDTH),
		32073 => to_signed(2182, LUT_AMPL_WIDTH),
		32074 => to_signed(2179, LUT_AMPL_WIDTH),
		32075 => to_signed(2175, LUT_AMPL_WIDTH),
		32076 => to_signed(2172, LUT_AMPL_WIDTH),
		32077 => to_signed(2169, LUT_AMPL_WIDTH),
		32078 => to_signed(2166, LUT_AMPL_WIDTH),
		32079 => to_signed(2163, LUT_AMPL_WIDTH),
		32080 => to_signed(2160, LUT_AMPL_WIDTH),
		32081 => to_signed(2157, LUT_AMPL_WIDTH),
		32082 => to_signed(2154, LUT_AMPL_WIDTH),
		32083 => to_signed(2150, LUT_AMPL_WIDTH),
		32084 => to_signed(2147, LUT_AMPL_WIDTH),
		32085 => to_signed(2144, LUT_AMPL_WIDTH),
		32086 => to_signed(2141, LUT_AMPL_WIDTH),
		32087 => to_signed(2138, LUT_AMPL_WIDTH),
		32088 => to_signed(2135, LUT_AMPL_WIDTH),
		32089 => to_signed(2132, LUT_AMPL_WIDTH),
		32090 => to_signed(2128, LUT_AMPL_WIDTH),
		32091 => to_signed(2125, LUT_AMPL_WIDTH),
		32092 => to_signed(2122, LUT_AMPL_WIDTH),
		32093 => to_signed(2119, LUT_AMPL_WIDTH),
		32094 => to_signed(2116, LUT_AMPL_WIDTH),
		32095 => to_signed(2113, LUT_AMPL_WIDTH),
		32096 => to_signed(2110, LUT_AMPL_WIDTH),
		32097 => to_signed(2106, LUT_AMPL_WIDTH),
		32098 => to_signed(2103, LUT_AMPL_WIDTH),
		32099 => to_signed(2100, LUT_AMPL_WIDTH),
		32100 => to_signed(2097, LUT_AMPL_WIDTH),
		32101 => to_signed(2094, LUT_AMPL_WIDTH),
		32102 => to_signed(2091, LUT_AMPL_WIDTH),
		32103 => to_signed(2088, LUT_AMPL_WIDTH),
		32104 => to_signed(2085, LUT_AMPL_WIDTH),
		32105 => to_signed(2081, LUT_AMPL_WIDTH),
		32106 => to_signed(2078, LUT_AMPL_WIDTH),
		32107 => to_signed(2075, LUT_AMPL_WIDTH),
		32108 => to_signed(2072, LUT_AMPL_WIDTH),
		32109 => to_signed(2069, LUT_AMPL_WIDTH),
		32110 => to_signed(2066, LUT_AMPL_WIDTH),
		32111 => to_signed(2063, LUT_AMPL_WIDTH),
		32112 => to_signed(2059, LUT_AMPL_WIDTH),
		32113 => to_signed(2056, LUT_AMPL_WIDTH),
		32114 => to_signed(2053, LUT_AMPL_WIDTH),
		32115 => to_signed(2050, LUT_AMPL_WIDTH),
		32116 => to_signed(2047, LUT_AMPL_WIDTH),
		32117 => to_signed(2044, LUT_AMPL_WIDTH),
		32118 => to_signed(2041, LUT_AMPL_WIDTH),
		32119 => to_signed(2038, LUT_AMPL_WIDTH),
		32120 => to_signed(2034, LUT_AMPL_WIDTH),
		32121 => to_signed(2031, LUT_AMPL_WIDTH),
		32122 => to_signed(2028, LUT_AMPL_WIDTH),
		32123 => to_signed(2025, LUT_AMPL_WIDTH),
		32124 => to_signed(2022, LUT_AMPL_WIDTH),
		32125 => to_signed(2019, LUT_AMPL_WIDTH),
		32126 => to_signed(2016, LUT_AMPL_WIDTH),
		32127 => to_signed(2012, LUT_AMPL_WIDTH),
		32128 => to_signed(2009, LUT_AMPL_WIDTH),
		32129 => to_signed(2006, LUT_AMPL_WIDTH),
		32130 => to_signed(2003, LUT_AMPL_WIDTH),
		32131 => to_signed(2000, LUT_AMPL_WIDTH),
		32132 => to_signed(1997, LUT_AMPL_WIDTH),
		32133 => to_signed(1994, LUT_AMPL_WIDTH),
		32134 => to_signed(1990, LUT_AMPL_WIDTH),
		32135 => to_signed(1987, LUT_AMPL_WIDTH),
		32136 => to_signed(1984, LUT_AMPL_WIDTH),
		32137 => to_signed(1981, LUT_AMPL_WIDTH),
		32138 => to_signed(1978, LUT_AMPL_WIDTH),
		32139 => to_signed(1975, LUT_AMPL_WIDTH),
		32140 => to_signed(1972, LUT_AMPL_WIDTH),
		32141 => to_signed(1969, LUT_AMPL_WIDTH),
		32142 => to_signed(1965, LUT_AMPL_WIDTH),
		32143 => to_signed(1962, LUT_AMPL_WIDTH),
		32144 => to_signed(1959, LUT_AMPL_WIDTH),
		32145 => to_signed(1956, LUT_AMPL_WIDTH),
		32146 => to_signed(1953, LUT_AMPL_WIDTH),
		32147 => to_signed(1950, LUT_AMPL_WIDTH),
		32148 => to_signed(1947, LUT_AMPL_WIDTH),
		32149 => to_signed(1943, LUT_AMPL_WIDTH),
		32150 => to_signed(1940, LUT_AMPL_WIDTH),
		32151 => to_signed(1937, LUT_AMPL_WIDTH),
		32152 => to_signed(1934, LUT_AMPL_WIDTH),
		32153 => to_signed(1931, LUT_AMPL_WIDTH),
		32154 => to_signed(1928, LUT_AMPL_WIDTH),
		32155 => to_signed(1925, LUT_AMPL_WIDTH),
		32156 => to_signed(1921, LUT_AMPL_WIDTH),
		32157 => to_signed(1918, LUT_AMPL_WIDTH),
		32158 => to_signed(1915, LUT_AMPL_WIDTH),
		32159 => to_signed(1912, LUT_AMPL_WIDTH),
		32160 => to_signed(1909, LUT_AMPL_WIDTH),
		32161 => to_signed(1906, LUT_AMPL_WIDTH),
		32162 => to_signed(1903, LUT_AMPL_WIDTH),
		32163 => to_signed(1900, LUT_AMPL_WIDTH),
		32164 => to_signed(1896, LUT_AMPL_WIDTH),
		32165 => to_signed(1893, LUT_AMPL_WIDTH),
		32166 => to_signed(1890, LUT_AMPL_WIDTH),
		32167 => to_signed(1887, LUT_AMPL_WIDTH),
		32168 => to_signed(1884, LUT_AMPL_WIDTH),
		32169 => to_signed(1881, LUT_AMPL_WIDTH),
		32170 => to_signed(1878, LUT_AMPL_WIDTH),
		32171 => to_signed(1874, LUT_AMPL_WIDTH),
		32172 => to_signed(1871, LUT_AMPL_WIDTH),
		32173 => to_signed(1868, LUT_AMPL_WIDTH),
		32174 => to_signed(1865, LUT_AMPL_WIDTH),
		32175 => to_signed(1862, LUT_AMPL_WIDTH),
		32176 => to_signed(1859, LUT_AMPL_WIDTH),
		32177 => to_signed(1856, LUT_AMPL_WIDTH),
		32178 => to_signed(1852, LUT_AMPL_WIDTH),
		32179 => to_signed(1849, LUT_AMPL_WIDTH),
		32180 => to_signed(1846, LUT_AMPL_WIDTH),
		32181 => to_signed(1843, LUT_AMPL_WIDTH),
		32182 => to_signed(1840, LUT_AMPL_WIDTH),
		32183 => to_signed(1837, LUT_AMPL_WIDTH),
		32184 => to_signed(1834, LUT_AMPL_WIDTH),
		32185 => to_signed(1831, LUT_AMPL_WIDTH),
		32186 => to_signed(1827, LUT_AMPL_WIDTH),
		32187 => to_signed(1824, LUT_AMPL_WIDTH),
		32188 => to_signed(1821, LUT_AMPL_WIDTH),
		32189 => to_signed(1818, LUT_AMPL_WIDTH),
		32190 => to_signed(1815, LUT_AMPL_WIDTH),
		32191 => to_signed(1812, LUT_AMPL_WIDTH),
		32192 => to_signed(1809, LUT_AMPL_WIDTH),
		32193 => to_signed(1805, LUT_AMPL_WIDTH),
		32194 => to_signed(1802, LUT_AMPL_WIDTH),
		32195 => to_signed(1799, LUT_AMPL_WIDTH),
		32196 => to_signed(1796, LUT_AMPL_WIDTH),
		32197 => to_signed(1793, LUT_AMPL_WIDTH),
		32198 => to_signed(1790, LUT_AMPL_WIDTH),
		32199 => to_signed(1787, LUT_AMPL_WIDTH),
		32200 => to_signed(1783, LUT_AMPL_WIDTH),
		32201 => to_signed(1780, LUT_AMPL_WIDTH),
		32202 => to_signed(1777, LUT_AMPL_WIDTH),
		32203 => to_signed(1774, LUT_AMPL_WIDTH),
		32204 => to_signed(1771, LUT_AMPL_WIDTH),
		32205 => to_signed(1768, LUT_AMPL_WIDTH),
		32206 => to_signed(1765, LUT_AMPL_WIDTH),
		32207 => to_signed(1762, LUT_AMPL_WIDTH),
		32208 => to_signed(1758, LUT_AMPL_WIDTH),
		32209 => to_signed(1755, LUT_AMPL_WIDTH),
		32210 => to_signed(1752, LUT_AMPL_WIDTH),
		32211 => to_signed(1749, LUT_AMPL_WIDTH),
		32212 => to_signed(1746, LUT_AMPL_WIDTH),
		32213 => to_signed(1743, LUT_AMPL_WIDTH),
		32214 => to_signed(1740, LUT_AMPL_WIDTH),
		32215 => to_signed(1736, LUT_AMPL_WIDTH),
		32216 => to_signed(1733, LUT_AMPL_WIDTH),
		32217 => to_signed(1730, LUT_AMPL_WIDTH),
		32218 => to_signed(1727, LUT_AMPL_WIDTH),
		32219 => to_signed(1724, LUT_AMPL_WIDTH),
		32220 => to_signed(1721, LUT_AMPL_WIDTH),
		32221 => to_signed(1718, LUT_AMPL_WIDTH),
		32222 => to_signed(1714, LUT_AMPL_WIDTH),
		32223 => to_signed(1711, LUT_AMPL_WIDTH),
		32224 => to_signed(1708, LUT_AMPL_WIDTH),
		32225 => to_signed(1705, LUT_AMPL_WIDTH),
		32226 => to_signed(1702, LUT_AMPL_WIDTH),
		32227 => to_signed(1699, LUT_AMPL_WIDTH),
		32228 => to_signed(1696, LUT_AMPL_WIDTH),
		32229 => to_signed(1693, LUT_AMPL_WIDTH),
		32230 => to_signed(1689, LUT_AMPL_WIDTH),
		32231 => to_signed(1686, LUT_AMPL_WIDTH),
		32232 => to_signed(1683, LUT_AMPL_WIDTH),
		32233 => to_signed(1680, LUT_AMPL_WIDTH),
		32234 => to_signed(1677, LUT_AMPL_WIDTH),
		32235 => to_signed(1674, LUT_AMPL_WIDTH),
		32236 => to_signed(1671, LUT_AMPL_WIDTH),
		32237 => to_signed(1667, LUT_AMPL_WIDTH),
		32238 => to_signed(1664, LUT_AMPL_WIDTH),
		32239 => to_signed(1661, LUT_AMPL_WIDTH),
		32240 => to_signed(1658, LUT_AMPL_WIDTH),
		32241 => to_signed(1655, LUT_AMPL_WIDTH),
		32242 => to_signed(1652, LUT_AMPL_WIDTH),
		32243 => to_signed(1649, LUT_AMPL_WIDTH),
		32244 => to_signed(1645, LUT_AMPL_WIDTH),
		32245 => to_signed(1642, LUT_AMPL_WIDTH),
		32246 => to_signed(1639, LUT_AMPL_WIDTH),
		32247 => to_signed(1636, LUT_AMPL_WIDTH),
		32248 => to_signed(1633, LUT_AMPL_WIDTH),
		32249 => to_signed(1630, LUT_AMPL_WIDTH),
		32250 => to_signed(1627, LUT_AMPL_WIDTH),
		32251 => to_signed(1623, LUT_AMPL_WIDTH),
		32252 => to_signed(1620, LUT_AMPL_WIDTH),
		32253 => to_signed(1617, LUT_AMPL_WIDTH),
		32254 => to_signed(1614, LUT_AMPL_WIDTH),
		32255 => to_signed(1611, LUT_AMPL_WIDTH),
		32256 => to_signed(1608, LUT_AMPL_WIDTH),
		32257 => to_signed(1605, LUT_AMPL_WIDTH),
		32258 => to_signed(1602, LUT_AMPL_WIDTH),
		32259 => to_signed(1598, LUT_AMPL_WIDTH),
		32260 => to_signed(1595, LUT_AMPL_WIDTH),
		32261 => to_signed(1592, LUT_AMPL_WIDTH),
		32262 => to_signed(1589, LUT_AMPL_WIDTH),
		32263 => to_signed(1586, LUT_AMPL_WIDTH),
		32264 => to_signed(1583, LUT_AMPL_WIDTH),
		32265 => to_signed(1580, LUT_AMPL_WIDTH),
		32266 => to_signed(1576, LUT_AMPL_WIDTH),
		32267 => to_signed(1573, LUT_AMPL_WIDTH),
		32268 => to_signed(1570, LUT_AMPL_WIDTH),
		32269 => to_signed(1567, LUT_AMPL_WIDTH),
		32270 => to_signed(1564, LUT_AMPL_WIDTH),
		32271 => to_signed(1561, LUT_AMPL_WIDTH),
		32272 => to_signed(1558, LUT_AMPL_WIDTH),
		32273 => to_signed(1554, LUT_AMPL_WIDTH),
		32274 => to_signed(1551, LUT_AMPL_WIDTH),
		32275 => to_signed(1548, LUT_AMPL_WIDTH),
		32276 => to_signed(1545, LUT_AMPL_WIDTH),
		32277 => to_signed(1542, LUT_AMPL_WIDTH),
		32278 => to_signed(1539, LUT_AMPL_WIDTH),
		32279 => to_signed(1536, LUT_AMPL_WIDTH),
		32280 => to_signed(1532, LUT_AMPL_WIDTH),
		32281 => to_signed(1529, LUT_AMPL_WIDTH),
		32282 => to_signed(1526, LUT_AMPL_WIDTH),
		32283 => to_signed(1523, LUT_AMPL_WIDTH),
		32284 => to_signed(1520, LUT_AMPL_WIDTH),
		32285 => to_signed(1517, LUT_AMPL_WIDTH),
		32286 => to_signed(1514, LUT_AMPL_WIDTH),
		32287 => to_signed(1511, LUT_AMPL_WIDTH),
		32288 => to_signed(1507, LUT_AMPL_WIDTH),
		32289 => to_signed(1504, LUT_AMPL_WIDTH),
		32290 => to_signed(1501, LUT_AMPL_WIDTH),
		32291 => to_signed(1498, LUT_AMPL_WIDTH),
		32292 => to_signed(1495, LUT_AMPL_WIDTH),
		32293 => to_signed(1492, LUT_AMPL_WIDTH),
		32294 => to_signed(1489, LUT_AMPL_WIDTH),
		32295 => to_signed(1485, LUT_AMPL_WIDTH),
		32296 => to_signed(1482, LUT_AMPL_WIDTH),
		32297 => to_signed(1479, LUT_AMPL_WIDTH),
		32298 => to_signed(1476, LUT_AMPL_WIDTH),
		32299 => to_signed(1473, LUT_AMPL_WIDTH),
		32300 => to_signed(1470, LUT_AMPL_WIDTH),
		32301 => to_signed(1467, LUT_AMPL_WIDTH),
		32302 => to_signed(1463, LUT_AMPL_WIDTH),
		32303 => to_signed(1460, LUT_AMPL_WIDTH),
		32304 => to_signed(1457, LUT_AMPL_WIDTH),
		32305 => to_signed(1454, LUT_AMPL_WIDTH),
		32306 => to_signed(1451, LUT_AMPL_WIDTH),
		32307 => to_signed(1448, LUT_AMPL_WIDTH),
		32308 => to_signed(1445, LUT_AMPL_WIDTH),
		32309 => to_signed(1441, LUT_AMPL_WIDTH),
		32310 => to_signed(1438, LUT_AMPL_WIDTH),
		32311 => to_signed(1435, LUT_AMPL_WIDTH),
		32312 => to_signed(1432, LUT_AMPL_WIDTH),
		32313 => to_signed(1429, LUT_AMPL_WIDTH),
		32314 => to_signed(1426, LUT_AMPL_WIDTH),
		32315 => to_signed(1423, LUT_AMPL_WIDTH),
		32316 => to_signed(1420, LUT_AMPL_WIDTH),
		32317 => to_signed(1416, LUT_AMPL_WIDTH),
		32318 => to_signed(1413, LUT_AMPL_WIDTH),
		32319 => to_signed(1410, LUT_AMPL_WIDTH),
		32320 => to_signed(1407, LUT_AMPL_WIDTH),
		32321 => to_signed(1404, LUT_AMPL_WIDTH),
		32322 => to_signed(1401, LUT_AMPL_WIDTH),
		32323 => to_signed(1398, LUT_AMPL_WIDTH),
		32324 => to_signed(1394, LUT_AMPL_WIDTH),
		32325 => to_signed(1391, LUT_AMPL_WIDTH),
		32326 => to_signed(1388, LUT_AMPL_WIDTH),
		32327 => to_signed(1385, LUT_AMPL_WIDTH),
		32328 => to_signed(1382, LUT_AMPL_WIDTH),
		32329 => to_signed(1379, LUT_AMPL_WIDTH),
		32330 => to_signed(1376, LUT_AMPL_WIDTH),
		32331 => to_signed(1372, LUT_AMPL_WIDTH),
		32332 => to_signed(1369, LUT_AMPL_WIDTH),
		32333 => to_signed(1366, LUT_AMPL_WIDTH),
		32334 => to_signed(1363, LUT_AMPL_WIDTH),
		32335 => to_signed(1360, LUT_AMPL_WIDTH),
		32336 => to_signed(1357, LUT_AMPL_WIDTH),
		32337 => to_signed(1354, LUT_AMPL_WIDTH),
		32338 => to_signed(1350, LUT_AMPL_WIDTH),
		32339 => to_signed(1347, LUT_AMPL_WIDTH),
		32340 => to_signed(1344, LUT_AMPL_WIDTH),
		32341 => to_signed(1341, LUT_AMPL_WIDTH),
		32342 => to_signed(1338, LUT_AMPL_WIDTH),
		32343 => to_signed(1335, LUT_AMPL_WIDTH),
		32344 => to_signed(1332, LUT_AMPL_WIDTH),
		32345 => to_signed(1328, LUT_AMPL_WIDTH),
		32346 => to_signed(1325, LUT_AMPL_WIDTH),
		32347 => to_signed(1322, LUT_AMPL_WIDTH),
		32348 => to_signed(1319, LUT_AMPL_WIDTH),
		32349 => to_signed(1316, LUT_AMPL_WIDTH),
		32350 => to_signed(1313, LUT_AMPL_WIDTH),
		32351 => to_signed(1310, LUT_AMPL_WIDTH),
		32352 => to_signed(1307, LUT_AMPL_WIDTH),
		32353 => to_signed(1303, LUT_AMPL_WIDTH),
		32354 => to_signed(1300, LUT_AMPL_WIDTH),
		32355 => to_signed(1297, LUT_AMPL_WIDTH),
		32356 => to_signed(1294, LUT_AMPL_WIDTH),
		32357 => to_signed(1291, LUT_AMPL_WIDTH),
		32358 => to_signed(1288, LUT_AMPL_WIDTH),
		32359 => to_signed(1285, LUT_AMPL_WIDTH),
		32360 => to_signed(1281, LUT_AMPL_WIDTH),
		32361 => to_signed(1278, LUT_AMPL_WIDTH),
		32362 => to_signed(1275, LUT_AMPL_WIDTH),
		32363 => to_signed(1272, LUT_AMPL_WIDTH),
		32364 => to_signed(1269, LUT_AMPL_WIDTH),
		32365 => to_signed(1266, LUT_AMPL_WIDTH),
		32366 => to_signed(1263, LUT_AMPL_WIDTH),
		32367 => to_signed(1259, LUT_AMPL_WIDTH),
		32368 => to_signed(1256, LUT_AMPL_WIDTH),
		32369 => to_signed(1253, LUT_AMPL_WIDTH),
		32370 => to_signed(1250, LUT_AMPL_WIDTH),
		32371 => to_signed(1247, LUT_AMPL_WIDTH),
		32372 => to_signed(1244, LUT_AMPL_WIDTH),
		32373 => to_signed(1241, LUT_AMPL_WIDTH),
		32374 => to_signed(1237, LUT_AMPL_WIDTH),
		32375 => to_signed(1234, LUT_AMPL_WIDTH),
		32376 => to_signed(1231, LUT_AMPL_WIDTH),
		32377 => to_signed(1228, LUT_AMPL_WIDTH),
		32378 => to_signed(1225, LUT_AMPL_WIDTH),
		32379 => to_signed(1222, LUT_AMPL_WIDTH),
		32380 => to_signed(1219, LUT_AMPL_WIDTH),
		32381 => to_signed(1215, LUT_AMPL_WIDTH),
		32382 => to_signed(1212, LUT_AMPL_WIDTH),
		32383 => to_signed(1209, LUT_AMPL_WIDTH),
		32384 => to_signed(1206, LUT_AMPL_WIDTH),
		32385 => to_signed(1203, LUT_AMPL_WIDTH),
		32386 => to_signed(1200, LUT_AMPL_WIDTH),
		32387 => to_signed(1197, LUT_AMPL_WIDTH),
		32388 => to_signed(1194, LUT_AMPL_WIDTH),
		32389 => to_signed(1190, LUT_AMPL_WIDTH),
		32390 => to_signed(1187, LUT_AMPL_WIDTH),
		32391 => to_signed(1184, LUT_AMPL_WIDTH),
		32392 => to_signed(1181, LUT_AMPL_WIDTH),
		32393 => to_signed(1178, LUT_AMPL_WIDTH),
		32394 => to_signed(1175, LUT_AMPL_WIDTH),
		32395 => to_signed(1172, LUT_AMPL_WIDTH),
		32396 => to_signed(1168, LUT_AMPL_WIDTH),
		32397 => to_signed(1165, LUT_AMPL_WIDTH),
		32398 => to_signed(1162, LUT_AMPL_WIDTH),
		32399 => to_signed(1159, LUT_AMPL_WIDTH),
		32400 => to_signed(1156, LUT_AMPL_WIDTH),
		32401 => to_signed(1153, LUT_AMPL_WIDTH),
		32402 => to_signed(1150, LUT_AMPL_WIDTH),
		32403 => to_signed(1146, LUT_AMPL_WIDTH),
		32404 => to_signed(1143, LUT_AMPL_WIDTH),
		32405 => to_signed(1140, LUT_AMPL_WIDTH),
		32406 => to_signed(1137, LUT_AMPL_WIDTH),
		32407 => to_signed(1134, LUT_AMPL_WIDTH),
		32408 => to_signed(1131, LUT_AMPL_WIDTH),
		32409 => to_signed(1128, LUT_AMPL_WIDTH),
		32410 => to_signed(1124, LUT_AMPL_WIDTH),
		32411 => to_signed(1121, LUT_AMPL_WIDTH),
		32412 => to_signed(1118, LUT_AMPL_WIDTH),
		32413 => to_signed(1115, LUT_AMPL_WIDTH),
		32414 => to_signed(1112, LUT_AMPL_WIDTH),
		32415 => to_signed(1109, LUT_AMPL_WIDTH),
		32416 => to_signed(1106, LUT_AMPL_WIDTH),
		32417 => to_signed(1102, LUT_AMPL_WIDTH),
		32418 => to_signed(1099, LUT_AMPL_WIDTH),
		32419 => to_signed(1096, LUT_AMPL_WIDTH),
		32420 => to_signed(1093, LUT_AMPL_WIDTH),
		32421 => to_signed(1090, LUT_AMPL_WIDTH),
		32422 => to_signed(1087, LUT_AMPL_WIDTH),
		32423 => to_signed(1084, LUT_AMPL_WIDTH),
		32424 => to_signed(1080, LUT_AMPL_WIDTH),
		32425 => to_signed(1077, LUT_AMPL_WIDTH),
		32426 => to_signed(1074, LUT_AMPL_WIDTH),
		32427 => to_signed(1071, LUT_AMPL_WIDTH),
		32428 => to_signed(1068, LUT_AMPL_WIDTH),
		32429 => to_signed(1065, LUT_AMPL_WIDTH),
		32430 => to_signed(1062, LUT_AMPL_WIDTH),
		32431 => to_signed(1059, LUT_AMPL_WIDTH),
		32432 => to_signed(1055, LUT_AMPL_WIDTH),
		32433 => to_signed(1052, LUT_AMPL_WIDTH),
		32434 => to_signed(1049, LUT_AMPL_WIDTH),
		32435 => to_signed(1046, LUT_AMPL_WIDTH),
		32436 => to_signed(1043, LUT_AMPL_WIDTH),
		32437 => to_signed(1040, LUT_AMPL_WIDTH),
		32438 => to_signed(1037, LUT_AMPL_WIDTH),
		32439 => to_signed(1033, LUT_AMPL_WIDTH),
		32440 => to_signed(1030, LUT_AMPL_WIDTH),
		32441 => to_signed(1027, LUT_AMPL_WIDTH),
		32442 => to_signed(1024, LUT_AMPL_WIDTH),
		32443 => to_signed(1021, LUT_AMPL_WIDTH),
		32444 => to_signed(1018, LUT_AMPL_WIDTH),
		32445 => to_signed(1015, LUT_AMPL_WIDTH),
		32446 => to_signed(1011, LUT_AMPL_WIDTH),
		32447 => to_signed(1008, LUT_AMPL_WIDTH),
		32448 => to_signed(1005, LUT_AMPL_WIDTH),
		32449 => to_signed(1002, LUT_AMPL_WIDTH),
		32450 => to_signed(999, LUT_AMPL_WIDTH),
		32451 => to_signed(996, LUT_AMPL_WIDTH),
		32452 => to_signed(993, LUT_AMPL_WIDTH),
		32453 => to_signed(989, LUT_AMPL_WIDTH),
		32454 => to_signed(986, LUT_AMPL_WIDTH),
		32455 => to_signed(983, LUT_AMPL_WIDTH),
		32456 => to_signed(980, LUT_AMPL_WIDTH),
		32457 => to_signed(977, LUT_AMPL_WIDTH),
		32458 => to_signed(974, LUT_AMPL_WIDTH),
		32459 => to_signed(971, LUT_AMPL_WIDTH),
		32460 => to_signed(967, LUT_AMPL_WIDTH),
		32461 => to_signed(964, LUT_AMPL_WIDTH),
		32462 => to_signed(961, LUT_AMPL_WIDTH),
		32463 => to_signed(958, LUT_AMPL_WIDTH),
		32464 => to_signed(955, LUT_AMPL_WIDTH),
		32465 => to_signed(952, LUT_AMPL_WIDTH),
		32466 => to_signed(949, LUT_AMPL_WIDTH),
		32467 => to_signed(945, LUT_AMPL_WIDTH),
		32468 => to_signed(942, LUT_AMPL_WIDTH),
		32469 => to_signed(939, LUT_AMPL_WIDTH),
		32470 => to_signed(936, LUT_AMPL_WIDTH),
		32471 => to_signed(933, LUT_AMPL_WIDTH),
		32472 => to_signed(930, LUT_AMPL_WIDTH),
		32473 => to_signed(927, LUT_AMPL_WIDTH),
		32474 => to_signed(923, LUT_AMPL_WIDTH),
		32475 => to_signed(920, LUT_AMPL_WIDTH),
		32476 => to_signed(917, LUT_AMPL_WIDTH),
		32477 => to_signed(914, LUT_AMPL_WIDTH),
		32478 => to_signed(911, LUT_AMPL_WIDTH),
		32479 => to_signed(908, LUT_AMPL_WIDTH),
		32480 => to_signed(905, LUT_AMPL_WIDTH),
		32481 => to_signed(901, LUT_AMPL_WIDTH),
		32482 => to_signed(898, LUT_AMPL_WIDTH),
		32483 => to_signed(895, LUT_AMPL_WIDTH),
		32484 => to_signed(892, LUT_AMPL_WIDTH),
		32485 => to_signed(889, LUT_AMPL_WIDTH),
		32486 => to_signed(886, LUT_AMPL_WIDTH),
		32487 => to_signed(883, LUT_AMPL_WIDTH),
		32488 => to_signed(880, LUT_AMPL_WIDTH),
		32489 => to_signed(876, LUT_AMPL_WIDTH),
		32490 => to_signed(873, LUT_AMPL_WIDTH),
		32491 => to_signed(870, LUT_AMPL_WIDTH),
		32492 => to_signed(867, LUT_AMPL_WIDTH),
		32493 => to_signed(864, LUT_AMPL_WIDTH),
		32494 => to_signed(861, LUT_AMPL_WIDTH),
		32495 => to_signed(858, LUT_AMPL_WIDTH),
		32496 => to_signed(854, LUT_AMPL_WIDTH),
		32497 => to_signed(851, LUT_AMPL_WIDTH),
		32498 => to_signed(848, LUT_AMPL_WIDTH),
		32499 => to_signed(845, LUT_AMPL_WIDTH),
		32500 => to_signed(842, LUT_AMPL_WIDTH),
		32501 => to_signed(839, LUT_AMPL_WIDTH),
		32502 => to_signed(836, LUT_AMPL_WIDTH),
		32503 => to_signed(832, LUT_AMPL_WIDTH),
		32504 => to_signed(829, LUT_AMPL_WIDTH),
		32505 => to_signed(826, LUT_AMPL_WIDTH),
		32506 => to_signed(823, LUT_AMPL_WIDTH),
		32507 => to_signed(820, LUT_AMPL_WIDTH),
		32508 => to_signed(817, LUT_AMPL_WIDTH),
		32509 => to_signed(814, LUT_AMPL_WIDTH),
		32510 => to_signed(810, LUT_AMPL_WIDTH),
		32511 => to_signed(807, LUT_AMPL_WIDTH),
		32512 => to_signed(804, LUT_AMPL_WIDTH),
		32513 => to_signed(801, LUT_AMPL_WIDTH),
		32514 => to_signed(798, LUT_AMPL_WIDTH),
		32515 => to_signed(795, LUT_AMPL_WIDTH),
		32516 => to_signed(792, LUT_AMPL_WIDTH),
		32517 => to_signed(788, LUT_AMPL_WIDTH),
		32518 => to_signed(785, LUT_AMPL_WIDTH),
		32519 => to_signed(782, LUT_AMPL_WIDTH),
		32520 => to_signed(779, LUT_AMPL_WIDTH),
		32521 => to_signed(776, LUT_AMPL_WIDTH),
		32522 => to_signed(773, LUT_AMPL_WIDTH),
		32523 => to_signed(770, LUT_AMPL_WIDTH),
		32524 => to_signed(766, LUT_AMPL_WIDTH),
		32525 => to_signed(763, LUT_AMPL_WIDTH),
		32526 => to_signed(760, LUT_AMPL_WIDTH),
		32527 => to_signed(757, LUT_AMPL_WIDTH),
		32528 => to_signed(754, LUT_AMPL_WIDTH),
		32529 => to_signed(751, LUT_AMPL_WIDTH),
		32530 => to_signed(748, LUT_AMPL_WIDTH),
		32531 => to_signed(744, LUT_AMPL_WIDTH),
		32532 => to_signed(741, LUT_AMPL_WIDTH),
		32533 => to_signed(738, LUT_AMPL_WIDTH),
		32534 => to_signed(735, LUT_AMPL_WIDTH),
		32535 => to_signed(732, LUT_AMPL_WIDTH),
		32536 => to_signed(729, LUT_AMPL_WIDTH),
		32537 => to_signed(726, LUT_AMPL_WIDTH),
		32538 => to_signed(722, LUT_AMPL_WIDTH),
		32539 => to_signed(719, LUT_AMPL_WIDTH),
		32540 => to_signed(716, LUT_AMPL_WIDTH),
		32541 => to_signed(713, LUT_AMPL_WIDTH),
		32542 => to_signed(710, LUT_AMPL_WIDTH),
		32543 => to_signed(707, LUT_AMPL_WIDTH),
		32544 => to_signed(704, LUT_AMPL_WIDTH),
		32545 => to_signed(701, LUT_AMPL_WIDTH),
		32546 => to_signed(697, LUT_AMPL_WIDTH),
		32547 => to_signed(694, LUT_AMPL_WIDTH),
		32548 => to_signed(691, LUT_AMPL_WIDTH),
		32549 => to_signed(688, LUT_AMPL_WIDTH),
		32550 => to_signed(685, LUT_AMPL_WIDTH),
		32551 => to_signed(682, LUT_AMPL_WIDTH),
		32552 => to_signed(679, LUT_AMPL_WIDTH),
		32553 => to_signed(675, LUT_AMPL_WIDTH),
		32554 => to_signed(672, LUT_AMPL_WIDTH),
		32555 => to_signed(669, LUT_AMPL_WIDTH),
		32556 => to_signed(666, LUT_AMPL_WIDTH),
		32557 => to_signed(663, LUT_AMPL_WIDTH),
		32558 => to_signed(660, LUT_AMPL_WIDTH),
		32559 => to_signed(657, LUT_AMPL_WIDTH),
		32560 => to_signed(653, LUT_AMPL_WIDTH),
		32561 => to_signed(650, LUT_AMPL_WIDTH),
		32562 => to_signed(647, LUT_AMPL_WIDTH),
		32563 => to_signed(644, LUT_AMPL_WIDTH),
		32564 => to_signed(641, LUT_AMPL_WIDTH),
		32565 => to_signed(638, LUT_AMPL_WIDTH),
		32566 => to_signed(635, LUT_AMPL_WIDTH),
		32567 => to_signed(631, LUT_AMPL_WIDTH),
		32568 => to_signed(628, LUT_AMPL_WIDTH),
		32569 => to_signed(625, LUT_AMPL_WIDTH),
		32570 => to_signed(622, LUT_AMPL_WIDTH),
		32571 => to_signed(619, LUT_AMPL_WIDTH),
		32572 => to_signed(616, LUT_AMPL_WIDTH),
		32573 => to_signed(613, LUT_AMPL_WIDTH),
		32574 => to_signed(609, LUT_AMPL_WIDTH),
		32575 => to_signed(606, LUT_AMPL_WIDTH),
		32576 => to_signed(603, LUT_AMPL_WIDTH),
		32577 => to_signed(600, LUT_AMPL_WIDTH),
		32578 => to_signed(597, LUT_AMPL_WIDTH),
		32579 => to_signed(594, LUT_AMPL_WIDTH),
		32580 => to_signed(591, LUT_AMPL_WIDTH),
		32581 => to_signed(587, LUT_AMPL_WIDTH),
		32582 => to_signed(584, LUT_AMPL_WIDTH),
		32583 => to_signed(581, LUT_AMPL_WIDTH),
		32584 => to_signed(578, LUT_AMPL_WIDTH),
		32585 => to_signed(575, LUT_AMPL_WIDTH),
		32586 => to_signed(572, LUT_AMPL_WIDTH),
		32587 => to_signed(569, LUT_AMPL_WIDTH),
		32588 => to_signed(565, LUT_AMPL_WIDTH),
		32589 => to_signed(562, LUT_AMPL_WIDTH),
		32590 => to_signed(559, LUT_AMPL_WIDTH),
		32591 => to_signed(556, LUT_AMPL_WIDTH),
		32592 => to_signed(553, LUT_AMPL_WIDTH),
		32593 => to_signed(550, LUT_AMPL_WIDTH),
		32594 => to_signed(547, LUT_AMPL_WIDTH),
		32595 => to_signed(543, LUT_AMPL_WIDTH),
		32596 => to_signed(540, LUT_AMPL_WIDTH),
		32597 => to_signed(537, LUT_AMPL_WIDTH),
		32598 => to_signed(534, LUT_AMPL_WIDTH),
		32599 => to_signed(531, LUT_AMPL_WIDTH),
		32600 => to_signed(528, LUT_AMPL_WIDTH),
		32601 => to_signed(525, LUT_AMPL_WIDTH),
		32602 => to_signed(521, LUT_AMPL_WIDTH),
		32603 => to_signed(518, LUT_AMPL_WIDTH),
		32604 => to_signed(515, LUT_AMPL_WIDTH),
		32605 => to_signed(512, LUT_AMPL_WIDTH),
		32606 => to_signed(509, LUT_AMPL_WIDTH),
		32607 => to_signed(506, LUT_AMPL_WIDTH),
		32608 => to_signed(503, LUT_AMPL_WIDTH),
		32609 => to_signed(499, LUT_AMPL_WIDTH),
		32610 => to_signed(496, LUT_AMPL_WIDTH),
		32611 => to_signed(493, LUT_AMPL_WIDTH),
		32612 => to_signed(490, LUT_AMPL_WIDTH),
		32613 => to_signed(487, LUT_AMPL_WIDTH),
		32614 => to_signed(484, LUT_AMPL_WIDTH),
		32615 => to_signed(481, LUT_AMPL_WIDTH),
		32616 => to_signed(477, LUT_AMPL_WIDTH),
		32617 => to_signed(474, LUT_AMPL_WIDTH),
		32618 => to_signed(471, LUT_AMPL_WIDTH),
		32619 => to_signed(468, LUT_AMPL_WIDTH),
		32620 => to_signed(465, LUT_AMPL_WIDTH),
		32621 => to_signed(462, LUT_AMPL_WIDTH),
		32622 => to_signed(459, LUT_AMPL_WIDTH),
		32623 => to_signed(456, LUT_AMPL_WIDTH),
		32624 => to_signed(452, LUT_AMPL_WIDTH),
		32625 => to_signed(449, LUT_AMPL_WIDTH),
		32626 => to_signed(446, LUT_AMPL_WIDTH),
		32627 => to_signed(443, LUT_AMPL_WIDTH),
		32628 => to_signed(440, LUT_AMPL_WIDTH),
		32629 => to_signed(437, LUT_AMPL_WIDTH),
		32630 => to_signed(434, LUT_AMPL_WIDTH),
		32631 => to_signed(430, LUT_AMPL_WIDTH),
		32632 => to_signed(427, LUT_AMPL_WIDTH),
		32633 => to_signed(424, LUT_AMPL_WIDTH),
		32634 => to_signed(421, LUT_AMPL_WIDTH),
		32635 => to_signed(418, LUT_AMPL_WIDTH),
		32636 => to_signed(415, LUT_AMPL_WIDTH),
		32637 => to_signed(412, LUT_AMPL_WIDTH),
		32638 => to_signed(408, LUT_AMPL_WIDTH),
		32639 => to_signed(405, LUT_AMPL_WIDTH),
		32640 => to_signed(402, LUT_AMPL_WIDTH),
		32641 => to_signed(399, LUT_AMPL_WIDTH),
		32642 => to_signed(396, LUT_AMPL_WIDTH),
		32643 => to_signed(393, LUT_AMPL_WIDTH),
		32644 => to_signed(390, LUT_AMPL_WIDTH),
		32645 => to_signed(386, LUT_AMPL_WIDTH),
		32646 => to_signed(383, LUT_AMPL_WIDTH),
		32647 => to_signed(380, LUT_AMPL_WIDTH),
		32648 => to_signed(377, LUT_AMPL_WIDTH),
		32649 => to_signed(374, LUT_AMPL_WIDTH),
		32650 => to_signed(371, LUT_AMPL_WIDTH),
		32651 => to_signed(368, LUT_AMPL_WIDTH),
		32652 => to_signed(364, LUT_AMPL_WIDTH),
		32653 => to_signed(361, LUT_AMPL_WIDTH),
		32654 => to_signed(358, LUT_AMPL_WIDTH),
		32655 => to_signed(355, LUT_AMPL_WIDTH),
		32656 => to_signed(352, LUT_AMPL_WIDTH),
		32657 => to_signed(349, LUT_AMPL_WIDTH),
		32658 => to_signed(346, LUT_AMPL_WIDTH),
		32659 => to_signed(342, LUT_AMPL_WIDTH),
		32660 => to_signed(339, LUT_AMPL_WIDTH),
		32661 => to_signed(336, LUT_AMPL_WIDTH),
		32662 => to_signed(333, LUT_AMPL_WIDTH),
		32663 => to_signed(330, LUT_AMPL_WIDTH),
		32664 => to_signed(327, LUT_AMPL_WIDTH),
		32665 => to_signed(324, LUT_AMPL_WIDTH),
		32666 => to_signed(320, LUT_AMPL_WIDTH),
		32667 => to_signed(317, LUT_AMPL_WIDTH),
		32668 => to_signed(314, LUT_AMPL_WIDTH),
		32669 => to_signed(311, LUT_AMPL_WIDTH),
		32670 => to_signed(308, LUT_AMPL_WIDTH),
		32671 => to_signed(305, LUT_AMPL_WIDTH),
		32672 => to_signed(302, LUT_AMPL_WIDTH),
		32673 => to_signed(298, LUT_AMPL_WIDTH),
		32674 => to_signed(295, LUT_AMPL_WIDTH),
		32675 => to_signed(292, LUT_AMPL_WIDTH),
		32676 => to_signed(289, LUT_AMPL_WIDTH),
		32677 => to_signed(286, LUT_AMPL_WIDTH),
		32678 => to_signed(283, LUT_AMPL_WIDTH),
		32679 => to_signed(280, LUT_AMPL_WIDTH),
		32680 => to_signed(276, LUT_AMPL_WIDTH),
		32681 => to_signed(273, LUT_AMPL_WIDTH),
		32682 => to_signed(270, LUT_AMPL_WIDTH),
		32683 => to_signed(267, LUT_AMPL_WIDTH),
		32684 => to_signed(264, LUT_AMPL_WIDTH),
		32685 => to_signed(261, LUT_AMPL_WIDTH),
		32686 => to_signed(258, LUT_AMPL_WIDTH),
		32687 => to_signed(254, LUT_AMPL_WIDTH),
		32688 => to_signed(251, LUT_AMPL_WIDTH),
		32689 => to_signed(248, LUT_AMPL_WIDTH),
		32690 => to_signed(245, LUT_AMPL_WIDTH),
		32691 => to_signed(242, LUT_AMPL_WIDTH),
		32692 => to_signed(239, LUT_AMPL_WIDTH),
		32693 => to_signed(236, LUT_AMPL_WIDTH),
		32694 => to_signed(232, LUT_AMPL_WIDTH),
		32695 => to_signed(229, LUT_AMPL_WIDTH),
		32696 => to_signed(226, LUT_AMPL_WIDTH),
		32697 => to_signed(223, LUT_AMPL_WIDTH),
		32698 => to_signed(220, LUT_AMPL_WIDTH),
		32699 => to_signed(217, LUT_AMPL_WIDTH),
		32700 => to_signed(214, LUT_AMPL_WIDTH),
		32701 => to_signed(210, LUT_AMPL_WIDTH),
		32702 => to_signed(207, LUT_AMPL_WIDTH),
		32703 => to_signed(204, LUT_AMPL_WIDTH),
		32704 => to_signed(201, LUT_AMPL_WIDTH),
		32705 => to_signed(198, LUT_AMPL_WIDTH),
		32706 => to_signed(195, LUT_AMPL_WIDTH),
		32707 => to_signed(192, LUT_AMPL_WIDTH),
		32708 => to_signed(188, LUT_AMPL_WIDTH),
		32709 => to_signed(185, LUT_AMPL_WIDTH),
		32710 => to_signed(182, LUT_AMPL_WIDTH),
		32711 => to_signed(179, LUT_AMPL_WIDTH),
		32712 => to_signed(176, LUT_AMPL_WIDTH),
		32713 => to_signed(173, LUT_AMPL_WIDTH),
		32714 => to_signed(170, LUT_AMPL_WIDTH),
		32715 => to_signed(166, LUT_AMPL_WIDTH),
		32716 => to_signed(163, LUT_AMPL_WIDTH),
		32717 => to_signed(160, LUT_AMPL_WIDTH),
		32718 => to_signed(157, LUT_AMPL_WIDTH),
		32719 => to_signed(154, LUT_AMPL_WIDTH),
		32720 => to_signed(151, LUT_AMPL_WIDTH),
		32721 => to_signed(148, LUT_AMPL_WIDTH),
		32722 => to_signed(145, LUT_AMPL_WIDTH),
		32723 => to_signed(141, LUT_AMPL_WIDTH),
		32724 => to_signed(138, LUT_AMPL_WIDTH),
		32725 => to_signed(135, LUT_AMPL_WIDTH),
		32726 => to_signed(132, LUT_AMPL_WIDTH),
		32727 => to_signed(129, LUT_AMPL_WIDTH),
		32728 => to_signed(126, LUT_AMPL_WIDTH),
		32729 => to_signed(123, LUT_AMPL_WIDTH),
		32730 => to_signed(119, LUT_AMPL_WIDTH),
		32731 => to_signed(116, LUT_AMPL_WIDTH),
		32732 => to_signed(113, LUT_AMPL_WIDTH),
		32733 => to_signed(110, LUT_AMPL_WIDTH),
		32734 => to_signed(107, LUT_AMPL_WIDTH),
		32735 => to_signed(104, LUT_AMPL_WIDTH),
		32736 => to_signed(101, LUT_AMPL_WIDTH),
		32737 => to_signed(97, LUT_AMPL_WIDTH),
		32738 => to_signed(94, LUT_AMPL_WIDTH),
		32739 => to_signed(91, LUT_AMPL_WIDTH),
		32740 => to_signed(88, LUT_AMPL_WIDTH),
		32741 => to_signed(85, LUT_AMPL_WIDTH),
		32742 => to_signed(82, LUT_AMPL_WIDTH),
		32743 => to_signed(79, LUT_AMPL_WIDTH),
		32744 => to_signed(75, LUT_AMPL_WIDTH),
		32745 => to_signed(72, LUT_AMPL_WIDTH),
		32746 => to_signed(69, LUT_AMPL_WIDTH),
		32747 => to_signed(66, LUT_AMPL_WIDTH),
		32748 => to_signed(63, LUT_AMPL_WIDTH),
		32749 => to_signed(60, LUT_AMPL_WIDTH),
		32750 => to_signed(57, LUT_AMPL_WIDTH),
		32751 => to_signed(53, LUT_AMPL_WIDTH),
		32752 => to_signed(50, LUT_AMPL_WIDTH),
		32753 => to_signed(47, LUT_AMPL_WIDTH),
		32754 => to_signed(44, LUT_AMPL_WIDTH),
		32755 => to_signed(41, LUT_AMPL_WIDTH),
		32756 => to_signed(38, LUT_AMPL_WIDTH),
		32757 => to_signed(35, LUT_AMPL_WIDTH),
		32758 => to_signed(31, LUT_AMPL_WIDTH),
		32759 => to_signed(28, LUT_AMPL_WIDTH),
		32760 => to_signed(25, LUT_AMPL_WIDTH),
		32761 => to_signed(22, LUT_AMPL_WIDTH),
		32762 => to_signed(19, LUT_AMPL_WIDTH),
		32763 => to_signed(16, LUT_AMPL_WIDTH),
		32764 => to_signed(13, LUT_AMPL_WIDTH),
		32765 => to_signed(9, LUT_AMPL_WIDTH),
		32766 => to_signed(6, LUT_AMPL_WIDTH),
		32767 => to_signed(3, LUT_AMPL_WIDTH),
		others => to_signed(0, LUT_AMPL_WIDTH)
);
end package sine_lut_pkg;

package body sine_lut_pkg is
end package body sine_lut_pkg;
