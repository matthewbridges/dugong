library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package sine_lut_pkg is

constant LUT_AMPL_WIDTH : natural := 16;
constant LUT_ADDR_WIDTH : natural := 15;

type lut_type is array (0 to 2 ** LUT_ADDR_WIDTH - 1) of unsigned(LUT_AMPL_WIDTH - 2 downto 0);
constant sine : lut_type := (
		0 => to_unsigned(0, LUT_AMPL_WIDTH - 1),
		1 => to_unsigned(3, LUT_AMPL_WIDTH - 1),
		2 => to_unsigned(6, LUT_AMPL_WIDTH - 1),
		3 => to_unsigned(9, LUT_AMPL_WIDTH - 1),
		4 => to_unsigned(13, LUT_AMPL_WIDTH - 1),
		5 => to_unsigned(16, LUT_AMPL_WIDTH - 1),
		6 => to_unsigned(19, LUT_AMPL_WIDTH - 1),
		7 => to_unsigned(22, LUT_AMPL_WIDTH - 1),
		8 => to_unsigned(25, LUT_AMPL_WIDTH - 1),
		9 => to_unsigned(28, LUT_AMPL_WIDTH - 1),
		10 => to_unsigned(31, LUT_AMPL_WIDTH - 1),
		11 => to_unsigned(35, LUT_AMPL_WIDTH - 1),
		12 => to_unsigned(38, LUT_AMPL_WIDTH - 1),
		13 => to_unsigned(41, LUT_AMPL_WIDTH - 1),
		14 => to_unsigned(44, LUT_AMPL_WIDTH - 1),
		15 => to_unsigned(47, LUT_AMPL_WIDTH - 1),
		16 => to_unsigned(50, LUT_AMPL_WIDTH - 1),
		17 => to_unsigned(53, LUT_AMPL_WIDTH - 1),
		18 => to_unsigned(57, LUT_AMPL_WIDTH - 1),
		19 => to_unsigned(60, LUT_AMPL_WIDTH - 1),
		20 => to_unsigned(63, LUT_AMPL_WIDTH - 1),
		21 => to_unsigned(66, LUT_AMPL_WIDTH - 1),
		22 => to_unsigned(69, LUT_AMPL_WIDTH - 1),
		23 => to_unsigned(72, LUT_AMPL_WIDTH - 1),
		24 => to_unsigned(75, LUT_AMPL_WIDTH - 1),
		25 => to_unsigned(79, LUT_AMPL_WIDTH - 1),
		26 => to_unsigned(82, LUT_AMPL_WIDTH - 1),
		27 => to_unsigned(85, LUT_AMPL_WIDTH - 1),
		28 => to_unsigned(88, LUT_AMPL_WIDTH - 1),
		29 => to_unsigned(91, LUT_AMPL_WIDTH - 1),
		30 => to_unsigned(94, LUT_AMPL_WIDTH - 1),
		31 => to_unsigned(97, LUT_AMPL_WIDTH - 1),
		32 => to_unsigned(101, LUT_AMPL_WIDTH - 1),
		33 => to_unsigned(104, LUT_AMPL_WIDTH - 1),
		34 => to_unsigned(107, LUT_AMPL_WIDTH - 1),
		35 => to_unsigned(110, LUT_AMPL_WIDTH - 1),
		36 => to_unsigned(113, LUT_AMPL_WIDTH - 1),
		37 => to_unsigned(116, LUT_AMPL_WIDTH - 1),
		38 => to_unsigned(119, LUT_AMPL_WIDTH - 1),
		39 => to_unsigned(123, LUT_AMPL_WIDTH - 1),
		40 => to_unsigned(126, LUT_AMPL_WIDTH - 1),
		41 => to_unsigned(129, LUT_AMPL_WIDTH - 1),
		42 => to_unsigned(132, LUT_AMPL_WIDTH - 1),
		43 => to_unsigned(135, LUT_AMPL_WIDTH - 1),
		44 => to_unsigned(138, LUT_AMPL_WIDTH - 1),
		45 => to_unsigned(141, LUT_AMPL_WIDTH - 1),
		46 => to_unsigned(145, LUT_AMPL_WIDTH - 1),
		47 => to_unsigned(148, LUT_AMPL_WIDTH - 1),
		48 => to_unsigned(151, LUT_AMPL_WIDTH - 1),
		49 => to_unsigned(154, LUT_AMPL_WIDTH - 1),
		50 => to_unsigned(157, LUT_AMPL_WIDTH - 1),
		51 => to_unsigned(160, LUT_AMPL_WIDTH - 1),
		52 => to_unsigned(163, LUT_AMPL_WIDTH - 1),
		53 => to_unsigned(166, LUT_AMPL_WIDTH - 1),
		54 => to_unsigned(170, LUT_AMPL_WIDTH - 1),
		55 => to_unsigned(173, LUT_AMPL_WIDTH - 1),
		56 => to_unsigned(176, LUT_AMPL_WIDTH - 1),
		57 => to_unsigned(179, LUT_AMPL_WIDTH - 1),
		58 => to_unsigned(182, LUT_AMPL_WIDTH - 1),
		59 => to_unsigned(185, LUT_AMPL_WIDTH - 1),
		60 => to_unsigned(188, LUT_AMPL_WIDTH - 1),
		61 => to_unsigned(192, LUT_AMPL_WIDTH - 1),
		62 => to_unsigned(195, LUT_AMPL_WIDTH - 1),
		63 => to_unsigned(198, LUT_AMPL_WIDTH - 1),
		64 => to_unsigned(201, LUT_AMPL_WIDTH - 1),
		65 => to_unsigned(204, LUT_AMPL_WIDTH - 1),
		66 => to_unsigned(207, LUT_AMPL_WIDTH - 1),
		67 => to_unsigned(210, LUT_AMPL_WIDTH - 1),
		68 => to_unsigned(214, LUT_AMPL_WIDTH - 1),
		69 => to_unsigned(217, LUT_AMPL_WIDTH - 1),
		70 => to_unsigned(220, LUT_AMPL_WIDTH - 1),
		71 => to_unsigned(223, LUT_AMPL_WIDTH - 1),
		72 => to_unsigned(226, LUT_AMPL_WIDTH - 1),
		73 => to_unsigned(229, LUT_AMPL_WIDTH - 1),
		74 => to_unsigned(232, LUT_AMPL_WIDTH - 1),
		75 => to_unsigned(236, LUT_AMPL_WIDTH - 1),
		76 => to_unsigned(239, LUT_AMPL_WIDTH - 1),
		77 => to_unsigned(242, LUT_AMPL_WIDTH - 1),
		78 => to_unsigned(245, LUT_AMPL_WIDTH - 1),
		79 => to_unsigned(248, LUT_AMPL_WIDTH - 1),
		80 => to_unsigned(251, LUT_AMPL_WIDTH - 1),
		81 => to_unsigned(254, LUT_AMPL_WIDTH - 1),
		82 => to_unsigned(258, LUT_AMPL_WIDTH - 1),
		83 => to_unsigned(261, LUT_AMPL_WIDTH - 1),
		84 => to_unsigned(264, LUT_AMPL_WIDTH - 1),
		85 => to_unsigned(267, LUT_AMPL_WIDTH - 1),
		86 => to_unsigned(270, LUT_AMPL_WIDTH - 1),
		87 => to_unsigned(273, LUT_AMPL_WIDTH - 1),
		88 => to_unsigned(276, LUT_AMPL_WIDTH - 1),
		89 => to_unsigned(280, LUT_AMPL_WIDTH - 1),
		90 => to_unsigned(283, LUT_AMPL_WIDTH - 1),
		91 => to_unsigned(286, LUT_AMPL_WIDTH - 1),
		92 => to_unsigned(289, LUT_AMPL_WIDTH - 1),
		93 => to_unsigned(292, LUT_AMPL_WIDTH - 1),
		94 => to_unsigned(295, LUT_AMPL_WIDTH - 1),
		95 => to_unsigned(298, LUT_AMPL_WIDTH - 1),
		96 => to_unsigned(302, LUT_AMPL_WIDTH - 1),
		97 => to_unsigned(305, LUT_AMPL_WIDTH - 1),
		98 => to_unsigned(308, LUT_AMPL_WIDTH - 1),
		99 => to_unsigned(311, LUT_AMPL_WIDTH - 1),
		100 => to_unsigned(314, LUT_AMPL_WIDTH - 1),
		101 => to_unsigned(317, LUT_AMPL_WIDTH - 1),
		102 => to_unsigned(320, LUT_AMPL_WIDTH - 1),
		103 => to_unsigned(324, LUT_AMPL_WIDTH - 1),
		104 => to_unsigned(327, LUT_AMPL_WIDTH - 1),
		105 => to_unsigned(330, LUT_AMPL_WIDTH - 1),
		106 => to_unsigned(333, LUT_AMPL_WIDTH - 1),
		107 => to_unsigned(336, LUT_AMPL_WIDTH - 1),
		108 => to_unsigned(339, LUT_AMPL_WIDTH - 1),
		109 => to_unsigned(342, LUT_AMPL_WIDTH - 1),
		110 => to_unsigned(346, LUT_AMPL_WIDTH - 1),
		111 => to_unsigned(349, LUT_AMPL_WIDTH - 1),
		112 => to_unsigned(352, LUT_AMPL_WIDTH - 1),
		113 => to_unsigned(355, LUT_AMPL_WIDTH - 1),
		114 => to_unsigned(358, LUT_AMPL_WIDTH - 1),
		115 => to_unsigned(361, LUT_AMPL_WIDTH - 1),
		116 => to_unsigned(364, LUT_AMPL_WIDTH - 1),
		117 => to_unsigned(368, LUT_AMPL_WIDTH - 1),
		118 => to_unsigned(371, LUT_AMPL_WIDTH - 1),
		119 => to_unsigned(374, LUT_AMPL_WIDTH - 1),
		120 => to_unsigned(377, LUT_AMPL_WIDTH - 1),
		121 => to_unsigned(380, LUT_AMPL_WIDTH - 1),
		122 => to_unsigned(383, LUT_AMPL_WIDTH - 1),
		123 => to_unsigned(386, LUT_AMPL_WIDTH - 1),
		124 => to_unsigned(390, LUT_AMPL_WIDTH - 1),
		125 => to_unsigned(393, LUT_AMPL_WIDTH - 1),
		126 => to_unsigned(396, LUT_AMPL_WIDTH - 1),
		127 => to_unsigned(399, LUT_AMPL_WIDTH - 1),
		128 => to_unsigned(402, LUT_AMPL_WIDTH - 1),
		129 => to_unsigned(405, LUT_AMPL_WIDTH - 1),
		130 => to_unsigned(408, LUT_AMPL_WIDTH - 1),
		131 => to_unsigned(412, LUT_AMPL_WIDTH - 1),
		132 => to_unsigned(415, LUT_AMPL_WIDTH - 1),
		133 => to_unsigned(418, LUT_AMPL_WIDTH - 1),
		134 => to_unsigned(421, LUT_AMPL_WIDTH - 1),
		135 => to_unsigned(424, LUT_AMPL_WIDTH - 1),
		136 => to_unsigned(427, LUT_AMPL_WIDTH - 1),
		137 => to_unsigned(430, LUT_AMPL_WIDTH - 1),
		138 => to_unsigned(434, LUT_AMPL_WIDTH - 1),
		139 => to_unsigned(437, LUT_AMPL_WIDTH - 1),
		140 => to_unsigned(440, LUT_AMPL_WIDTH - 1),
		141 => to_unsigned(443, LUT_AMPL_WIDTH - 1),
		142 => to_unsigned(446, LUT_AMPL_WIDTH - 1),
		143 => to_unsigned(449, LUT_AMPL_WIDTH - 1),
		144 => to_unsigned(452, LUT_AMPL_WIDTH - 1),
		145 => to_unsigned(456, LUT_AMPL_WIDTH - 1),
		146 => to_unsigned(459, LUT_AMPL_WIDTH - 1),
		147 => to_unsigned(462, LUT_AMPL_WIDTH - 1),
		148 => to_unsigned(465, LUT_AMPL_WIDTH - 1),
		149 => to_unsigned(468, LUT_AMPL_WIDTH - 1),
		150 => to_unsigned(471, LUT_AMPL_WIDTH - 1),
		151 => to_unsigned(474, LUT_AMPL_WIDTH - 1),
		152 => to_unsigned(477, LUT_AMPL_WIDTH - 1),
		153 => to_unsigned(481, LUT_AMPL_WIDTH - 1),
		154 => to_unsigned(484, LUT_AMPL_WIDTH - 1),
		155 => to_unsigned(487, LUT_AMPL_WIDTH - 1),
		156 => to_unsigned(490, LUT_AMPL_WIDTH - 1),
		157 => to_unsigned(493, LUT_AMPL_WIDTH - 1),
		158 => to_unsigned(496, LUT_AMPL_WIDTH - 1),
		159 => to_unsigned(499, LUT_AMPL_WIDTH - 1),
		160 => to_unsigned(503, LUT_AMPL_WIDTH - 1),
		161 => to_unsigned(506, LUT_AMPL_WIDTH - 1),
		162 => to_unsigned(509, LUT_AMPL_WIDTH - 1),
		163 => to_unsigned(512, LUT_AMPL_WIDTH - 1),
		164 => to_unsigned(515, LUT_AMPL_WIDTH - 1),
		165 => to_unsigned(518, LUT_AMPL_WIDTH - 1),
		166 => to_unsigned(521, LUT_AMPL_WIDTH - 1),
		167 => to_unsigned(525, LUT_AMPL_WIDTH - 1),
		168 => to_unsigned(528, LUT_AMPL_WIDTH - 1),
		169 => to_unsigned(531, LUT_AMPL_WIDTH - 1),
		170 => to_unsigned(534, LUT_AMPL_WIDTH - 1),
		171 => to_unsigned(537, LUT_AMPL_WIDTH - 1),
		172 => to_unsigned(540, LUT_AMPL_WIDTH - 1),
		173 => to_unsigned(543, LUT_AMPL_WIDTH - 1),
		174 => to_unsigned(547, LUT_AMPL_WIDTH - 1),
		175 => to_unsigned(550, LUT_AMPL_WIDTH - 1),
		176 => to_unsigned(553, LUT_AMPL_WIDTH - 1),
		177 => to_unsigned(556, LUT_AMPL_WIDTH - 1),
		178 => to_unsigned(559, LUT_AMPL_WIDTH - 1),
		179 => to_unsigned(562, LUT_AMPL_WIDTH - 1),
		180 => to_unsigned(565, LUT_AMPL_WIDTH - 1),
		181 => to_unsigned(569, LUT_AMPL_WIDTH - 1),
		182 => to_unsigned(572, LUT_AMPL_WIDTH - 1),
		183 => to_unsigned(575, LUT_AMPL_WIDTH - 1),
		184 => to_unsigned(578, LUT_AMPL_WIDTH - 1),
		185 => to_unsigned(581, LUT_AMPL_WIDTH - 1),
		186 => to_unsigned(584, LUT_AMPL_WIDTH - 1),
		187 => to_unsigned(587, LUT_AMPL_WIDTH - 1),
		188 => to_unsigned(591, LUT_AMPL_WIDTH - 1),
		189 => to_unsigned(594, LUT_AMPL_WIDTH - 1),
		190 => to_unsigned(597, LUT_AMPL_WIDTH - 1),
		191 => to_unsigned(600, LUT_AMPL_WIDTH - 1),
		192 => to_unsigned(603, LUT_AMPL_WIDTH - 1),
		193 => to_unsigned(606, LUT_AMPL_WIDTH - 1),
		194 => to_unsigned(609, LUT_AMPL_WIDTH - 1),
		195 => to_unsigned(613, LUT_AMPL_WIDTH - 1),
		196 => to_unsigned(616, LUT_AMPL_WIDTH - 1),
		197 => to_unsigned(619, LUT_AMPL_WIDTH - 1),
		198 => to_unsigned(622, LUT_AMPL_WIDTH - 1),
		199 => to_unsigned(625, LUT_AMPL_WIDTH - 1),
		200 => to_unsigned(628, LUT_AMPL_WIDTH - 1),
		201 => to_unsigned(631, LUT_AMPL_WIDTH - 1),
		202 => to_unsigned(635, LUT_AMPL_WIDTH - 1),
		203 => to_unsigned(638, LUT_AMPL_WIDTH - 1),
		204 => to_unsigned(641, LUT_AMPL_WIDTH - 1),
		205 => to_unsigned(644, LUT_AMPL_WIDTH - 1),
		206 => to_unsigned(647, LUT_AMPL_WIDTH - 1),
		207 => to_unsigned(650, LUT_AMPL_WIDTH - 1),
		208 => to_unsigned(653, LUT_AMPL_WIDTH - 1),
		209 => to_unsigned(657, LUT_AMPL_WIDTH - 1),
		210 => to_unsigned(660, LUT_AMPL_WIDTH - 1),
		211 => to_unsigned(663, LUT_AMPL_WIDTH - 1),
		212 => to_unsigned(666, LUT_AMPL_WIDTH - 1),
		213 => to_unsigned(669, LUT_AMPL_WIDTH - 1),
		214 => to_unsigned(672, LUT_AMPL_WIDTH - 1),
		215 => to_unsigned(675, LUT_AMPL_WIDTH - 1),
		216 => to_unsigned(679, LUT_AMPL_WIDTH - 1),
		217 => to_unsigned(682, LUT_AMPL_WIDTH - 1),
		218 => to_unsigned(685, LUT_AMPL_WIDTH - 1),
		219 => to_unsigned(688, LUT_AMPL_WIDTH - 1),
		220 => to_unsigned(691, LUT_AMPL_WIDTH - 1),
		221 => to_unsigned(694, LUT_AMPL_WIDTH - 1),
		222 => to_unsigned(697, LUT_AMPL_WIDTH - 1),
		223 => to_unsigned(701, LUT_AMPL_WIDTH - 1),
		224 => to_unsigned(704, LUT_AMPL_WIDTH - 1),
		225 => to_unsigned(707, LUT_AMPL_WIDTH - 1),
		226 => to_unsigned(710, LUT_AMPL_WIDTH - 1),
		227 => to_unsigned(713, LUT_AMPL_WIDTH - 1),
		228 => to_unsigned(716, LUT_AMPL_WIDTH - 1),
		229 => to_unsigned(719, LUT_AMPL_WIDTH - 1),
		230 => to_unsigned(722, LUT_AMPL_WIDTH - 1),
		231 => to_unsigned(726, LUT_AMPL_WIDTH - 1),
		232 => to_unsigned(729, LUT_AMPL_WIDTH - 1),
		233 => to_unsigned(732, LUT_AMPL_WIDTH - 1),
		234 => to_unsigned(735, LUT_AMPL_WIDTH - 1),
		235 => to_unsigned(738, LUT_AMPL_WIDTH - 1),
		236 => to_unsigned(741, LUT_AMPL_WIDTH - 1),
		237 => to_unsigned(744, LUT_AMPL_WIDTH - 1),
		238 => to_unsigned(748, LUT_AMPL_WIDTH - 1),
		239 => to_unsigned(751, LUT_AMPL_WIDTH - 1),
		240 => to_unsigned(754, LUT_AMPL_WIDTH - 1),
		241 => to_unsigned(757, LUT_AMPL_WIDTH - 1),
		242 => to_unsigned(760, LUT_AMPL_WIDTH - 1),
		243 => to_unsigned(763, LUT_AMPL_WIDTH - 1),
		244 => to_unsigned(766, LUT_AMPL_WIDTH - 1),
		245 => to_unsigned(770, LUT_AMPL_WIDTH - 1),
		246 => to_unsigned(773, LUT_AMPL_WIDTH - 1),
		247 => to_unsigned(776, LUT_AMPL_WIDTH - 1),
		248 => to_unsigned(779, LUT_AMPL_WIDTH - 1),
		249 => to_unsigned(782, LUT_AMPL_WIDTH - 1),
		250 => to_unsigned(785, LUT_AMPL_WIDTH - 1),
		251 => to_unsigned(788, LUT_AMPL_WIDTH - 1),
		252 => to_unsigned(792, LUT_AMPL_WIDTH - 1),
		253 => to_unsigned(795, LUT_AMPL_WIDTH - 1),
		254 => to_unsigned(798, LUT_AMPL_WIDTH - 1),
		255 => to_unsigned(801, LUT_AMPL_WIDTH - 1),
		256 => to_unsigned(804, LUT_AMPL_WIDTH - 1),
		257 => to_unsigned(807, LUT_AMPL_WIDTH - 1),
		258 => to_unsigned(810, LUT_AMPL_WIDTH - 1),
		259 => to_unsigned(814, LUT_AMPL_WIDTH - 1),
		260 => to_unsigned(817, LUT_AMPL_WIDTH - 1),
		261 => to_unsigned(820, LUT_AMPL_WIDTH - 1),
		262 => to_unsigned(823, LUT_AMPL_WIDTH - 1),
		263 => to_unsigned(826, LUT_AMPL_WIDTH - 1),
		264 => to_unsigned(829, LUT_AMPL_WIDTH - 1),
		265 => to_unsigned(832, LUT_AMPL_WIDTH - 1),
		266 => to_unsigned(836, LUT_AMPL_WIDTH - 1),
		267 => to_unsigned(839, LUT_AMPL_WIDTH - 1),
		268 => to_unsigned(842, LUT_AMPL_WIDTH - 1),
		269 => to_unsigned(845, LUT_AMPL_WIDTH - 1),
		270 => to_unsigned(848, LUT_AMPL_WIDTH - 1),
		271 => to_unsigned(851, LUT_AMPL_WIDTH - 1),
		272 => to_unsigned(854, LUT_AMPL_WIDTH - 1),
		273 => to_unsigned(858, LUT_AMPL_WIDTH - 1),
		274 => to_unsigned(861, LUT_AMPL_WIDTH - 1),
		275 => to_unsigned(864, LUT_AMPL_WIDTH - 1),
		276 => to_unsigned(867, LUT_AMPL_WIDTH - 1),
		277 => to_unsigned(870, LUT_AMPL_WIDTH - 1),
		278 => to_unsigned(873, LUT_AMPL_WIDTH - 1),
		279 => to_unsigned(876, LUT_AMPL_WIDTH - 1),
		280 => to_unsigned(880, LUT_AMPL_WIDTH - 1),
		281 => to_unsigned(883, LUT_AMPL_WIDTH - 1),
		282 => to_unsigned(886, LUT_AMPL_WIDTH - 1),
		283 => to_unsigned(889, LUT_AMPL_WIDTH - 1),
		284 => to_unsigned(892, LUT_AMPL_WIDTH - 1),
		285 => to_unsigned(895, LUT_AMPL_WIDTH - 1),
		286 => to_unsigned(898, LUT_AMPL_WIDTH - 1),
		287 => to_unsigned(901, LUT_AMPL_WIDTH - 1),
		288 => to_unsigned(905, LUT_AMPL_WIDTH - 1),
		289 => to_unsigned(908, LUT_AMPL_WIDTH - 1),
		290 => to_unsigned(911, LUT_AMPL_WIDTH - 1),
		291 => to_unsigned(914, LUT_AMPL_WIDTH - 1),
		292 => to_unsigned(917, LUT_AMPL_WIDTH - 1),
		293 => to_unsigned(920, LUT_AMPL_WIDTH - 1),
		294 => to_unsigned(923, LUT_AMPL_WIDTH - 1),
		295 => to_unsigned(927, LUT_AMPL_WIDTH - 1),
		296 => to_unsigned(930, LUT_AMPL_WIDTH - 1),
		297 => to_unsigned(933, LUT_AMPL_WIDTH - 1),
		298 => to_unsigned(936, LUT_AMPL_WIDTH - 1),
		299 => to_unsigned(939, LUT_AMPL_WIDTH - 1),
		300 => to_unsigned(942, LUT_AMPL_WIDTH - 1),
		301 => to_unsigned(945, LUT_AMPL_WIDTH - 1),
		302 => to_unsigned(949, LUT_AMPL_WIDTH - 1),
		303 => to_unsigned(952, LUT_AMPL_WIDTH - 1),
		304 => to_unsigned(955, LUT_AMPL_WIDTH - 1),
		305 => to_unsigned(958, LUT_AMPL_WIDTH - 1),
		306 => to_unsigned(961, LUT_AMPL_WIDTH - 1),
		307 => to_unsigned(964, LUT_AMPL_WIDTH - 1),
		308 => to_unsigned(967, LUT_AMPL_WIDTH - 1),
		309 => to_unsigned(971, LUT_AMPL_WIDTH - 1),
		310 => to_unsigned(974, LUT_AMPL_WIDTH - 1),
		311 => to_unsigned(977, LUT_AMPL_WIDTH - 1),
		312 => to_unsigned(980, LUT_AMPL_WIDTH - 1),
		313 => to_unsigned(983, LUT_AMPL_WIDTH - 1),
		314 => to_unsigned(986, LUT_AMPL_WIDTH - 1),
		315 => to_unsigned(989, LUT_AMPL_WIDTH - 1),
		316 => to_unsigned(993, LUT_AMPL_WIDTH - 1),
		317 => to_unsigned(996, LUT_AMPL_WIDTH - 1),
		318 => to_unsigned(999, LUT_AMPL_WIDTH - 1),
		319 => to_unsigned(1002, LUT_AMPL_WIDTH - 1),
		320 => to_unsigned(1005, LUT_AMPL_WIDTH - 1),
		321 => to_unsigned(1008, LUT_AMPL_WIDTH - 1),
		322 => to_unsigned(1011, LUT_AMPL_WIDTH - 1),
		323 => to_unsigned(1015, LUT_AMPL_WIDTH - 1),
		324 => to_unsigned(1018, LUT_AMPL_WIDTH - 1),
		325 => to_unsigned(1021, LUT_AMPL_WIDTH - 1),
		326 => to_unsigned(1024, LUT_AMPL_WIDTH - 1),
		327 => to_unsigned(1027, LUT_AMPL_WIDTH - 1),
		328 => to_unsigned(1030, LUT_AMPL_WIDTH - 1),
		329 => to_unsigned(1033, LUT_AMPL_WIDTH - 1),
		330 => to_unsigned(1037, LUT_AMPL_WIDTH - 1),
		331 => to_unsigned(1040, LUT_AMPL_WIDTH - 1),
		332 => to_unsigned(1043, LUT_AMPL_WIDTH - 1),
		333 => to_unsigned(1046, LUT_AMPL_WIDTH - 1),
		334 => to_unsigned(1049, LUT_AMPL_WIDTH - 1),
		335 => to_unsigned(1052, LUT_AMPL_WIDTH - 1),
		336 => to_unsigned(1055, LUT_AMPL_WIDTH - 1),
		337 => to_unsigned(1059, LUT_AMPL_WIDTH - 1),
		338 => to_unsigned(1062, LUT_AMPL_WIDTH - 1),
		339 => to_unsigned(1065, LUT_AMPL_WIDTH - 1),
		340 => to_unsigned(1068, LUT_AMPL_WIDTH - 1),
		341 => to_unsigned(1071, LUT_AMPL_WIDTH - 1),
		342 => to_unsigned(1074, LUT_AMPL_WIDTH - 1),
		343 => to_unsigned(1077, LUT_AMPL_WIDTH - 1),
		344 => to_unsigned(1080, LUT_AMPL_WIDTH - 1),
		345 => to_unsigned(1084, LUT_AMPL_WIDTH - 1),
		346 => to_unsigned(1087, LUT_AMPL_WIDTH - 1),
		347 => to_unsigned(1090, LUT_AMPL_WIDTH - 1),
		348 => to_unsigned(1093, LUT_AMPL_WIDTH - 1),
		349 => to_unsigned(1096, LUT_AMPL_WIDTH - 1),
		350 => to_unsigned(1099, LUT_AMPL_WIDTH - 1),
		351 => to_unsigned(1102, LUT_AMPL_WIDTH - 1),
		352 => to_unsigned(1106, LUT_AMPL_WIDTH - 1),
		353 => to_unsigned(1109, LUT_AMPL_WIDTH - 1),
		354 => to_unsigned(1112, LUT_AMPL_WIDTH - 1),
		355 => to_unsigned(1115, LUT_AMPL_WIDTH - 1),
		356 => to_unsigned(1118, LUT_AMPL_WIDTH - 1),
		357 => to_unsigned(1121, LUT_AMPL_WIDTH - 1),
		358 => to_unsigned(1124, LUT_AMPL_WIDTH - 1),
		359 => to_unsigned(1128, LUT_AMPL_WIDTH - 1),
		360 => to_unsigned(1131, LUT_AMPL_WIDTH - 1),
		361 => to_unsigned(1134, LUT_AMPL_WIDTH - 1),
		362 => to_unsigned(1137, LUT_AMPL_WIDTH - 1),
		363 => to_unsigned(1140, LUT_AMPL_WIDTH - 1),
		364 => to_unsigned(1143, LUT_AMPL_WIDTH - 1),
		365 => to_unsigned(1146, LUT_AMPL_WIDTH - 1),
		366 => to_unsigned(1150, LUT_AMPL_WIDTH - 1),
		367 => to_unsigned(1153, LUT_AMPL_WIDTH - 1),
		368 => to_unsigned(1156, LUT_AMPL_WIDTH - 1),
		369 => to_unsigned(1159, LUT_AMPL_WIDTH - 1),
		370 => to_unsigned(1162, LUT_AMPL_WIDTH - 1),
		371 => to_unsigned(1165, LUT_AMPL_WIDTH - 1),
		372 => to_unsigned(1168, LUT_AMPL_WIDTH - 1),
		373 => to_unsigned(1172, LUT_AMPL_WIDTH - 1),
		374 => to_unsigned(1175, LUT_AMPL_WIDTH - 1),
		375 => to_unsigned(1178, LUT_AMPL_WIDTH - 1),
		376 => to_unsigned(1181, LUT_AMPL_WIDTH - 1),
		377 => to_unsigned(1184, LUT_AMPL_WIDTH - 1),
		378 => to_unsigned(1187, LUT_AMPL_WIDTH - 1),
		379 => to_unsigned(1190, LUT_AMPL_WIDTH - 1),
		380 => to_unsigned(1194, LUT_AMPL_WIDTH - 1),
		381 => to_unsigned(1197, LUT_AMPL_WIDTH - 1),
		382 => to_unsigned(1200, LUT_AMPL_WIDTH - 1),
		383 => to_unsigned(1203, LUT_AMPL_WIDTH - 1),
		384 => to_unsigned(1206, LUT_AMPL_WIDTH - 1),
		385 => to_unsigned(1209, LUT_AMPL_WIDTH - 1),
		386 => to_unsigned(1212, LUT_AMPL_WIDTH - 1),
		387 => to_unsigned(1215, LUT_AMPL_WIDTH - 1),
		388 => to_unsigned(1219, LUT_AMPL_WIDTH - 1),
		389 => to_unsigned(1222, LUT_AMPL_WIDTH - 1),
		390 => to_unsigned(1225, LUT_AMPL_WIDTH - 1),
		391 => to_unsigned(1228, LUT_AMPL_WIDTH - 1),
		392 => to_unsigned(1231, LUT_AMPL_WIDTH - 1),
		393 => to_unsigned(1234, LUT_AMPL_WIDTH - 1),
		394 => to_unsigned(1237, LUT_AMPL_WIDTH - 1),
		395 => to_unsigned(1241, LUT_AMPL_WIDTH - 1),
		396 => to_unsigned(1244, LUT_AMPL_WIDTH - 1),
		397 => to_unsigned(1247, LUT_AMPL_WIDTH - 1),
		398 => to_unsigned(1250, LUT_AMPL_WIDTH - 1),
		399 => to_unsigned(1253, LUT_AMPL_WIDTH - 1),
		400 => to_unsigned(1256, LUT_AMPL_WIDTH - 1),
		401 => to_unsigned(1259, LUT_AMPL_WIDTH - 1),
		402 => to_unsigned(1263, LUT_AMPL_WIDTH - 1),
		403 => to_unsigned(1266, LUT_AMPL_WIDTH - 1),
		404 => to_unsigned(1269, LUT_AMPL_WIDTH - 1),
		405 => to_unsigned(1272, LUT_AMPL_WIDTH - 1),
		406 => to_unsigned(1275, LUT_AMPL_WIDTH - 1),
		407 => to_unsigned(1278, LUT_AMPL_WIDTH - 1),
		408 => to_unsigned(1281, LUT_AMPL_WIDTH - 1),
		409 => to_unsigned(1285, LUT_AMPL_WIDTH - 1),
		410 => to_unsigned(1288, LUT_AMPL_WIDTH - 1),
		411 => to_unsigned(1291, LUT_AMPL_WIDTH - 1),
		412 => to_unsigned(1294, LUT_AMPL_WIDTH - 1),
		413 => to_unsigned(1297, LUT_AMPL_WIDTH - 1),
		414 => to_unsigned(1300, LUT_AMPL_WIDTH - 1),
		415 => to_unsigned(1303, LUT_AMPL_WIDTH - 1),
		416 => to_unsigned(1307, LUT_AMPL_WIDTH - 1),
		417 => to_unsigned(1310, LUT_AMPL_WIDTH - 1),
		418 => to_unsigned(1313, LUT_AMPL_WIDTH - 1),
		419 => to_unsigned(1316, LUT_AMPL_WIDTH - 1),
		420 => to_unsigned(1319, LUT_AMPL_WIDTH - 1),
		421 => to_unsigned(1322, LUT_AMPL_WIDTH - 1),
		422 => to_unsigned(1325, LUT_AMPL_WIDTH - 1),
		423 => to_unsigned(1328, LUT_AMPL_WIDTH - 1),
		424 => to_unsigned(1332, LUT_AMPL_WIDTH - 1),
		425 => to_unsigned(1335, LUT_AMPL_WIDTH - 1),
		426 => to_unsigned(1338, LUT_AMPL_WIDTH - 1),
		427 => to_unsigned(1341, LUT_AMPL_WIDTH - 1),
		428 => to_unsigned(1344, LUT_AMPL_WIDTH - 1),
		429 => to_unsigned(1347, LUT_AMPL_WIDTH - 1),
		430 => to_unsigned(1350, LUT_AMPL_WIDTH - 1),
		431 => to_unsigned(1354, LUT_AMPL_WIDTH - 1),
		432 => to_unsigned(1357, LUT_AMPL_WIDTH - 1),
		433 => to_unsigned(1360, LUT_AMPL_WIDTH - 1),
		434 => to_unsigned(1363, LUT_AMPL_WIDTH - 1),
		435 => to_unsigned(1366, LUT_AMPL_WIDTH - 1),
		436 => to_unsigned(1369, LUT_AMPL_WIDTH - 1),
		437 => to_unsigned(1372, LUT_AMPL_WIDTH - 1),
		438 => to_unsigned(1376, LUT_AMPL_WIDTH - 1),
		439 => to_unsigned(1379, LUT_AMPL_WIDTH - 1),
		440 => to_unsigned(1382, LUT_AMPL_WIDTH - 1),
		441 => to_unsigned(1385, LUT_AMPL_WIDTH - 1),
		442 => to_unsigned(1388, LUT_AMPL_WIDTH - 1),
		443 => to_unsigned(1391, LUT_AMPL_WIDTH - 1),
		444 => to_unsigned(1394, LUT_AMPL_WIDTH - 1),
		445 => to_unsigned(1398, LUT_AMPL_WIDTH - 1),
		446 => to_unsigned(1401, LUT_AMPL_WIDTH - 1),
		447 => to_unsigned(1404, LUT_AMPL_WIDTH - 1),
		448 => to_unsigned(1407, LUT_AMPL_WIDTH - 1),
		449 => to_unsigned(1410, LUT_AMPL_WIDTH - 1),
		450 => to_unsigned(1413, LUT_AMPL_WIDTH - 1),
		451 => to_unsigned(1416, LUT_AMPL_WIDTH - 1),
		452 => to_unsigned(1420, LUT_AMPL_WIDTH - 1),
		453 => to_unsigned(1423, LUT_AMPL_WIDTH - 1),
		454 => to_unsigned(1426, LUT_AMPL_WIDTH - 1),
		455 => to_unsigned(1429, LUT_AMPL_WIDTH - 1),
		456 => to_unsigned(1432, LUT_AMPL_WIDTH - 1),
		457 => to_unsigned(1435, LUT_AMPL_WIDTH - 1),
		458 => to_unsigned(1438, LUT_AMPL_WIDTH - 1),
		459 => to_unsigned(1441, LUT_AMPL_WIDTH - 1),
		460 => to_unsigned(1445, LUT_AMPL_WIDTH - 1),
		461 => to_unsigned(1448, LUT_AMPL_WIDTH - 1),
		462 => to_unsigned(1451, LUT_AMPL_WIDTH - 1),
		463 => to_unsigned(1454, LUT_AMPL_WIDTH - 1),
		464 => to_unsigned(1457, LUT_AMPL_WIDTH - 1),
		465 => to_unsigned(1460, LUT_AMPL_WIDTH - 1),
		466 => to_unsigned(1463, LUT_AMPL_WIDTH - 1),
		467 => to_unsigned(1467, LUT_AMPL_WIDTH - 1),
		468 => to_unsigned(1470, LUT_AMPL_WIDTH - 1),
		469 => to_unsigned(1473, LUT_AMPL_WIDTH - 1),
		470 => to_unsigned(1476, LUT_AMPL_WIDTH - 1),
		471 => to_unsigned(1479, LUT_AMPL_WIDTH - 1),
		472 => to_unsigned(1482, LUT_AMPL_WIDTH - 1),
		473 => to_unsigned(1485, LUT_AMPL_WIDTH - 1),
		474 => to_unsigned(1489, LUT_AMPL_WIDTH - 1),
		475 => to_unsigned(1492, LUT_AMPL_WIDTH - 1),
		476 => to_unsigned(1495, LUT_AMPL_WIDTH - 1),
		477 => to_unsigned(1498, LUT_AMPL_WIDTH - 1),
		478 => to_unsigned(1501, LUT_AMPL_WIDTH - 1),
		479 => to_unsigned(1504, LUT_AMPL_WIDTH - 1),
		480 => to_unsigned(1507, LUT_AMPL_WIDTH - 1),
		481 => to_unsigned(1511, LUT_AMPL_WIDTH - 1),
		482 => to_unsigned(1514, LUT_AMPL_WIDTH - 1),
		483 => to_unsigned(1517, LUT_AMPL_WIDTH - 1),
		484 => to_unsigned(1520, LUT_AMPL_WIDTH - 1),
		485 => to_unsigned(1523, LUT_AMPL_WIDTH - 1),
		486 => to_unsigned(1526, LUT_AMPL_WIDTH - 1),
		487 => to_unsigned(1529, LUT_AMPL_WIDTH - 1),
		488 => to_unsigned(1532, LUT_AMPL_WIDTH - 1),
		489 => to_unsigned(1536, LUT_AMPL_WIDTH - 1),
		490 => to_unsigned(1539, LUT_AMPL_WIDTH - 1),
		491 => to_unsigned(1542, LUT_AMPL_WIDTH - 1),
		492 => to_unsigned(1545, LUT_AMPL_WIDTH - 1),
		493 => to_unsigned(1548, LUT_AMPL_WIDTH - 1),
		494 => to_unsigned(1551, LUT_AMPL_WIDTH - 1),
		495 => to_unsigned(1554, LUT_AMPL_WIDTH - 1),
		496 => to_unsigned(1558, LUT_AMPL_WIDTH - 1),
		497 => to_unsigned(1561, LUT_AMPL_WIDTH - 1),
		498 => to_unsigned(1564, LUT_AMPL_WIDTH - 1),
		499 => to_unsigned(1567, LUT_AMPL_WIDTH - 1),
		500 => to_unsigned(1570, LUT_AMPL_WIDTH - 1),
		501 => to_unsigned(1573, LUT_AMPL_WIDTH - 1),
		502 => to_unsigned(1576, LUT_AMPL_WIDTH - 1),
		503 => to_unsigned(1580, LUT_AMPL_WIDTH - 1),
		504 => to_unsigned(1583, LUT_AMPL_WIDTH - 1),
		505 => to_unsigned(1586, LUT_AMPL_WIDTH - 1),
		506 => to_unsigned(1589, LUT_AMPL_WIDTH - 1),
		507 => to_unsigned(1592, LUT_AMPL_WIDTH - 1),
		508 => to_unsigned(1595, LUT_AMPL_WIDTH - 1),
		509 => to_unsigned(1598, LUT_AMPL_WIDTH - 1),
		510 => to_unsigned(1602, LUT_AMPL_WIDTH - 1),
		511 => to_unsigned(1605, LUT_AMPL_WIDTH - 1),
		512 => to_unsigned(1608, LUT_AMPL_WIDTH - 1),
		513 => to_unsigned(1611, LUT_AMPL_WIDTH - 1),
		514 => to_unsigned(1614, LUT_AMPL_WIDTH - 1),
		515 => to_unsigned(1617, LUT_AMPL_WIDTH - 1),
		516 => to_unsigned(1620, LUT_AMPL_WIDTH - 1),
		517 => to_unsigned(1623, LUT_AMPL_WIDTH - 1),
		518 => to_unsigned(1627, LUT_AMPL_WIDTH - 1),
		519 => to_unsigned(1630, LUT_AMPL_WIDTH - 1),
		520 => to_unsigned(1633, LUT_AMPL_WIDTH - 1),
		521 => to_unsigned(1636, LUT_AMPL_WIDTH - 1),
		522 => to_unsigned(1639, LUT_AMPL_WIDTH - 1),
		523 => to_unsigned(1642, LUT_AMPL_WIDTH - 1),
		524 => to_unsigned(1645, LUT_AMPL_WIDTH - 1),
		525 => to_unsigned(1649, LUT_AMPL_WIDTH - 1),
		526 => to_unsigned(1652, LUT_AMPL_WIDTH - 1),
		527 => to_unsigned(1655, LUT_AMPL_WIDTH - 1),
		528 => to_unsigned(1658, LUT_AMPL_WIDTH - 1),
		529 => to_unsigned(1661, LUT_AMPL_WIDTH - 1),
		530 => to_unsigned(1664, LUT_AMPL_WIDTH - 1),
		531 => to_unsigned(1667, LUT_AMPL_WIDTH - 1),
		532 => to_unsigned(1671, LUT_AMPL_WIDTH - 1),
		533 => to_unsigned(1674, LUT_AMPL_WIDTH - 1),
		534 => to_unsigned(1677, LUT_AMPL_WIDTH - 1),
		535 => to_unsigned(1680, LUT_AMPL_WIDTH - 1),
		536 => to_unsigned(1683, LUT_AMPL_WIDTH - 1),
		537 => to_unsigned(1686, LUT_AMPL_WIDTH - 1),
		538 => to_unsigned(1689, LUT_AMPL_WIDTH - 1),
		539 => to_unsigned(1693, LUT_AMPL_WIDTH - 1),
		540 => to_unsigned(1696, LUT_AMPL_WIDTH - 1),
		541 => to_unsigned(1699, LUT_AMPL_WIDTH - 1),
		542 => to_unsigned(1702, LUT_AMPL_WIDTH - 1),
		543 => to_unsigned(1705, LUT_AMPL_WIDTH - 1),
		544 => to_unsigned(1708, LUT_AMPL_WIDTH - 1),
		545 => to_unsigned(1711, LUT_AMPL_WIDTH - 1),
		546 => to_unsigned(1714, LUT_AMPL_WIDTH - 1),
		547 => to_unsigned(1718, LUT_AMPL_WIDTH - 1),
		548 => to_unsigned(1721, LUT_AMPL_WIDTH - 1),
		549 => to_unsigned(1724, LUT_AMPL_WIDTH - 1),
		550 => to_unsigned(1727, LUT_AMPL_WIDTH - 1),
		551 => to_unsigned(1730, LUT_AMPL_WIDTH - 1),
		552 => to_unsigned(1733, LUT_AMPL_WIDTH - 1),
		553 => to_unsigned(1736, LUT_AMPL_WIDTH - 1),
		554 => to_unsigned(1740, LUT_AMPL_WIDTH - 1),
		555 => to_unsigned(1743, LUT_AMPL_WIDTH - 1),
		556 => to_unsigned(1746, LUT_AMPL_WIDTH - 1),
		557 => to_unsigned(1749, LUT_AMPL_WIDTH - 1),
		558 => to_unsigned(1752, LUT_AMPL_WIDTH - 1),
		559 => to_unsigned(1755, LUT_AMPL_WIDTH - 1),
		560 => to_unsigned(1758, LUT_AMPL_WIDTH - 1),
		561 => to_unsigned(1762, LUT_AMPL_WIDTH - 1),
		562 => to_unsigned(1765, LUT_AMPL_WIDTH - 1),
		563 => to_unsigned(1768, LUT_AMPL_WIDTH - 1),
		564 => to_unsigned(1771, LUT_AMPL_WIDTH - 1),
		565 => to_unsigned(1774, LUT_AMPL_WIDTH - 1),
		566 => to_unsigned(1777, LUT_AMPL_WIDTH - 1),
		567 => to_unsigned(1780, LUT_AMPL_WIDTH - 1),
		568 => to_unsigned(1783, LUT_AMPL_WIDTH - 1),
		569 => to_unsigned(1787, LUT_AMPL_WIDTH - 1),
		570 => to_unsigned(1790, LUT_AMPL_WIDTH - 1),
		571 => to_unsigned(1793, LUT_AMPL_WIDTH - 1),
		572 => to_unsigned(1796, LUT_AMPL_WIDTH - 1),
		573 => to_unsigned(1799, LUT_AMPL_WIDTH - 1),
		574 => to_unsigned(1802, LUT_AMPL_WIDTH - 1),
		575 => to_unsigned(1805, LUT_AMPL_WIDTH - 1),
		576 => to_unsigned(1809, LUT_AMPL_WIDTH - 1),
		577 => to_unsigned(1812, LUT_AMPL_WIDTH - 1),
		578 => to_unsigned(1815, LUT_AMPL_WIDTH - 1),
		579 => to_unsigned(1818, LUT_AMPL_WIDTH - 1),
		580 => to_unsigned(1821, LUT_AMPL_WIDTH - 1),
		581 => to_unsigned(1824, LUT_AMPL_WIDTH - 1),
		582 => to_unsigned(1827, LUT_AMPL_WIDTH - 1),
		583 => to_unsigned(1831, LUT_AMPL_WIDTH - 1),
		584 => to_unsigned(1834, LUT_AMPL_WIDTH - 1),
		585 => to_unsigned(1837, LUT_AMPL_WIDTH - 1),
		586 => to_unsigned(1840, LUT_AMPL_WIDTH - 1),
		587 => to_unsigned(1843, LUT_AMPL_WIDTH - 1),
		588 => to_unsigned(1846, LUT_AMPL_WIDTH - 1),
		589 => to_unsigned(1849, LUT_AMPL_WIDTH - 1),
		590 => to_unsigned(1852, LUT_AMPL_WIDTH - 1),
		591 => to_unsigned(1856, LUT_AMPL_WIDTH - 1),
		592 => to_unsigned(1859, LUT_AMPL_WIDTH - 1),
		593 => to_unsigned(1862, LUT_AMPL_WIDTH - 1),
		594 => to_unsigned(1865, LUT_AMPL_WIDTH - 1),
		595 => to_unsigned(1868, LUT_AMPL_WIDTH - 1),
		596 => to_unsigned(1871, LUT_AMPL_WIDTH - 1),
		597 => to_unsigned(1874, LUT_AMPL_WIDTH - 1),
		598 => to_unsigned(1878, LUT_AMPL_WIDTH - 1),
		599 => to_unsigned(1881, LUT_AMPL_WIDTH - 1),
		600 => to_unsigned(1884, LUT_AMPL_WIDTH - 1),
		601 => to_unsigned(1887, LUT_AMPL_WIDTH - 1),
		602 => to_unsigned(1890, LUT_AMPL_WIDTH - 1),
		603 => to_unsigned(1893, LUT_AMPL_WIDTH - 1),
		604 => to_unsigned(1896, LUT_AMPL_WIDTH - 1),
		605 => to_unsigned(1900, LUT_AMPL_WIDTH - 1),
		606 => to_unsigned(1903, LUT_AMPL_WIDTH - 1),
		607 => to_unsigned(1906, LUT_AMPL_WIDTH - 1),
		608 => to_unsigned(1909, LUT_AMPL_WIDTH - 1),
		609 => to_unsigned(1912, LUT_AMPL_WIDTH - 1),
		610 => to_unsigned(1915, LUT_AMPL_WIDTH - 1),
		611 => to_unsigned(1918, LUT_AMPL_WIDTH - 1),
		612 => to_unsigned(1921, LUT_AMPL_WIDTH - 1),
		613 => to_unsigned(1925, LUT_AMPL_WIDTH - 1),
		614 => to_unsigned(1928, LUT_AMPL_WIDTH - 1),
		615 => to_unsigned(1931, LUT_AMPL_WIDTH - 1),
		616 => to_unsigned(1934, LUT_AMPL_WIDTH - 1),
		617 => to_unsigned(1937, LUT_AMPL_WIDTH - 1),
		618 => to_unsigned(1940, LUT_AMPL_WIDTH - 1),
		619 => to_unsigned(1943, LUT_AMPL_WIDTH - 1),
		620 => to_unsigned(1947, LUT_AMPL_WIDTH - 1),
		621 => to_unsigned(1950, LUT_AMPL_WIDTH - 1),
		622 => to_unsigned(1953, LUT_AMPL_WIDTH - 1),
		623 => to_unsigned(1956, LUT_AMPL_WIDTH - 1),
		624 => to_unsigned(1959, LUT_AMPL_WIDTH - 1),
		625 => to_unsigned(1962, LUT_AMPL_WIDTH - 1),
		626 => to_unsigned(1965, LUT_AMPL_WIDTH - 1),
		627 => to_unsigned(1969, LUT_AMPL_WIDTH - 1),
		628 => to_unsigned(1972, LUT_AMPL_WIDTH - 1),
		629 => to_unsigned(1975, LUT_AMPL_WIDTH - 1),
		630 => to_unsigned(1978, LUT_AMPL_WIDTH - 1),
		631 => to_unsigned(1981, LUT_AMPL_WIDTH - 1),
		632 => to_unsigned(1984, LUT_AMPL_WIDTH - 1),
		633 => to_unsigned(1987, LUT_AMPL_WIDTH - 1),
		634 => to_unsigned(1990, LUT_AMPL_WIDTH - 1),
		635 => to_unsigned(1994, LUT_AMPL_WIDTH - 1),
		636 => to_unsigned(1997, LUT_AMPL_WIDTH - 1),
		637 => to_unsigned(2000, LUT_AMPL_WIDTH - 1),
		638 => to_unsigned(2003, LUT_AMPL_WIDTH - 1),
		639 => to_unsigned(2006, LUT_AMPL_WIDTH - 1),
		640 => to_unsigned(2009, LUT_AMPL_WIDTH - 1),
		641 => to_unsigned(2012, LUT_AMPL_WIDTH - 1),
		642 => to_unsigned(2016, LUT_AMPL_WIDTH - 1),
		643 => to_unsigned(2019, LUT_AMPL_WIDTH - 1),
		644 => to_unsigned(2022, LUT_AMPL_WIDTH - 1),
		645 => to_unsigned(2025, LUT_AMPL_WIDTH - 1),
		646 => to_unsigned(2028, LUT_AMPL_WIDTH - 1),
		647 => to_unsigned(2031, LUT_AMPL_WIDTH - 1),
		648 => to_unsigned(2034, LUT_AMPL_WIDTH - 1),
		649 => to_unsigned(2038, LUT_AMPL_WIDTH - 1),
		650 => to_unsigned(2041, LUT_AMPL_WIDTH - 1),
		651 => to_unsigned(2044, LUT_AMPL_WIDTH - 1),
		652 => to_unsigned(2047, LUT_AMPL_WIDTH - 1),
		653 => to_unsigned(2050, LUT_AMPL_WIDTH - 1),
		654 => to_unsigned(2053, LUT_AMPL_WIDTH - 1),
		655 => to_unsigned(2056, LUT_AMPL_WIDTH - 1),
		656 => to_unsigned(2059, LUT_AMPL_WIDTH - 1),
		657 => to_unsigned(2063, LUT_AMPL_WIDTH - 1),
		658 => to_unsigned(2066, LUT_AMPL_WIDTH - 1),
		659 => to_unsigned(2069, LUT_AMPL_WIDTH - 1),
		660 => to_unsigned(2072, LUT_AMPL_WIDTH - 1),
		661 => to_unsigned(2075, LUT_AMPL_WIDTH - 1),
		662 => to_unsigned(2078, LUT_AMPL_WIDTH - 1),
		663 => to_unsigned(2081, LUT_AMPL_WIDTH - 1),
		664 => to_unsigned(2085, LUT_AMPL_WIDTH - 1),
		665 => to_unsigned(2088, LUT_AMPL_WIDTH - 1),
		666 => to_unsigned(2091, LUT_AMPL_WIDTH - 1),
		667 => to_unsigned(2094, LUT_AMPL_WIDTH - 1),
		668 => to_unsigned(2097, LUT_AMPL_WIDTH - 1),
		669 => to_unsigned(2100, LUT_AMPL_WIDTH - 1),
		670 => to_unsigned(2103, LUT_AMPL_WIDTH - 1),
		671 => to_unsigned(2106, LUT_AMPL_WIDTH - 1),
		672 => to_unsigned(2110, LUT_AMPL_WIDTH - 1),
		673 => to_unsigned(2113, LUT_AMPL_WIDTH - 1),
		674 => to_unsigned(2116, LUT_AMPL_WIDTH - 1),
		675 => to_unsigned(2119, LUT_AMPL_WIDTH - 1),
		676 => to_unsigned(2122, LUT_AMPL_WIDTH - 1),
		677 => to_unsigned(2125, LUT_AMPL_WIDTH - 1),
		678 => to_unsigned(2128, LUT_AMPL_WIDTH - 1),
		679 => to_unsigned(2132, LUT_AMPL_WIDTH - 1),
		680 => to_unsigned(2135, LUT_AMPL_WIDTH - 1),
		681 => to_unsigned(2138, LUT_AMPL_WIDTH - 1),
		682 => to_unsigned(2141, LUT_AMPL_WIDTH - 1),
		683 => to_unsigned(2144, LUT_AMPL_WIDTH - 1),
		684 => to_unsigned(2147, LUT_AMPL_WIDTH - 1),
		685 => to_unsigned(2150, LUT_AMPL_WIDTH - 1),
		686 => to_unsigned(2154, LUT_AMPL_WIDTH - 1),
		687 => to_unsigned(2157, LUT_AMPL_WIDTH - 1),
		688 => to_unsigned(2160, LUT_AMPL_WIDTH - 1),
		689 => to_unsigned(2163, LUT_AMPL_WIDTH - 1),
		690 => to_unsigned(2166, LUT_AMPL_WIDTH - 1),
		691 => to_unsigned(2169, LUT_AMPL_WIDTH - 1),
		692 => to_unsigned(2172, LUT_AMPL_WIDTH - 1),
		693 => to_unsigned(2175, LUT_AMPL_WIDTH - 1),
		694 => to_unsigned(2179, LUT_AMPL_WIDTH - 1),
		695 => to_unsigned(2182, LUT_AMPL_WIDTH - 1),
		696 => to_unsigned(2185, LUT_AMPL_WIDTH - 1),
		697 => to_unsigned(2188, LUT_AMPL_WIDTH - 1),
		698 => to_unsigned(2191, LUT_AMPL_WIDTH - 1),
		699 => to_unsigned(2194, LUT_AMPL_WIDTH - 1),
		700 => to_unsigned(2197, LUT_AMPL_WIDTH - 1),
		701 => to_unsigned(2201, LUT_AMPL_WIDTH - 1),
		702 => to_unsigned(2204, LUT_AMPL_WIDTH - 1),
		703 => to_unsigned(2207, LUT_AMPL_WIDTH - 1),
		704 => to_unsigned(2210, LUT_AMPL_WIDTH - 1),
		705 => to_unsigned(2213, LUT_AMPL_WIDTH - 1),
		706 => to_unsigned(2216, LUT_AMPL_WIDTH - 1),
		707 => to_unsigned(2219, LUT_AMPL_WIDTH - 1),
		708 => to_unsigned(2222, LUT_AMPL_WIDTH - 1),
		709 => to_unsigned(2226, LUT_AMPL_WIDTH - 1),
		710 => to_unsigned(2229, LUT_AMPL_WIDTH - 1),
		711 => to_unsigned(2232, LUT_AMPL_WIDTH - 1),
		712 => to_unsigned(2235, LUT_AMPL_WIDTH - 1),
		713 => to_unsigned(2238, LUT_AMPL_WIDTH - 1),
		714 => to_unsigned(2241, LUT_AMPL_WIDTH - 1),
		715 => to_unsigned(2244, LUT_AMPL_WIDTH - 1),
		716 => to_unsigned(2248, LUT_AMPL_WIDTH - 1),
		717 => to_unsigned(2251, LUT_AMPL_WIDTH - 1),
		718 => to_unsigned(2254, LUT_AMPL_WIDTH - 1),
		719 => to_unsigned(2257, LUT_AMPL_WIDTH - 1),
		720 => to_unsigned(2260, LUT_AMPL_WIDTH - 1),
		721 => to_unsigned(2263, LUT_AMPL_WIDTH - 1),
		722 => to_unsigned(2266, LUT_AMPL_WIDTH - 1),
		723 => to_unsigned(2269, LUT_AMPL_WIDTH - 1),
		724 => to_unsigned(2273, LUT_AMPL_WIDTH - 1),
		725 => to_unsigned(2276, LUT_AMPL_WIDTH - 1),
		726 => to_unsigned(2279, LUT_AMPL_WIDTH - 1),
		727 => to_unsigned(2282, LUT_AMPL_WIDTH - 1),
		728 => to_unsigned(2285, LUT_AMPL_WIDTH - 1),
		729 => to_unsigned(2288, LUT_AMPL_WIDTH - 1),
		730 => to_unsigned(2291, LUT_AMPL_WIDTH - 1),
		731 => to_unsigned(2295, LUT_AMPL_WIDTH - 1),
		732 => to_unsigned(2298, LUT_AMPL_WIDTH - 1),
		733 => to_unsigned(2301, LUT_AMPL_WIDTH - 1),
		734 => to_unsigned(2304, LUT_AMPL_WIDTH - 1),
		735 => to_unsigned(2307, LUT_AMPL_WIDTH - 1),
		736 => to_unsigned(2310, LUT_AMPL_WIDTH - 1),
		737 => to_unsigned(2313, LUT_AMPL_WIDTH - 1),
		738 => to_unsigned(2316, LUT_AMPL_WIDTH - 1),
		739 => to_unsigned(2320, LUT_AMPL_WIDTH - 1),
		740 => to_unsigned(2323, LUT_AMPL_WIDTH - 1),
		741 => to_unsigned(2326, LUT_AMPL_WIDTH - 1),
		742 => to_unsigned(2329, LUT_AMPL_WIDTH - 1),
		743 => to_unsigned(2332, LUT_AMPL_WIDTH - 1),
		744 => to_unsigned(2335, LUT_AMPL_WIDTH - 1),
		745 => to_unsigned(2338, LUT_AMPL_WIDTH - 1),
		746 => to_unsigned(2342, LUT_AMPL_WIDTH - 1),
		747 => to_unsigned(2345, LUT_AMPL_WIDTH - 1),
		748 => to_unsigned(2348, LUT_AMPL_WIDTH - 1),
		749 => to_unsigned(2351, LUT_AMPL_WIDTH - 1),
		750 => to_unsigned(2354, LUT_AMPL_WIDTH - 1),
		751 => to_unsigned(2357, LUT_AMPL_WIDTH - 1),
		752 => to_unsigned(2360, LUT_AMPL_WIDTH - 1),
		753 => to_unsigned(2363, LUT_AMPL_WIDTH - 1),
		754 => to_unsigned(2367, LUT_AMPL_WIDTH - 1),
		755 => to_unsigned(2370, LUT_AMPL_WIDTH - 1),
		756 => to_unsigned(2373, LUT_AMPL_WIDTH - 1),
		757 => to_unsigned(2376, LUT_AMPL_WIDTH - 1),
		758 => to_unsigned(2379, LUT_AMPL_WIDTH - 1),
		759 => to_unsigned(2382, LUT_AMPL_WIDTH - 1),
		760 => to_unsigned(2385, LUT_AMPL_WIDTH - 1),
		761 => to_unsigned(2389, LUT_AMPL_WIDTH - 1),
		762 => to_unsigned(2392, LUT_AMPL_WIDTH - 1),
		763 => to_unsigned(2395, LUT_AMPL_WIDTH - 1),
		764 => to_unsigned(2398, LUT_AMPL_WIDTH - 1),
		765 => to_unsigned(2401, LUT_AMPL_WIDTH - 1),
		766 => to_unsigned(2404, LUT_AMPL_WIDTH - 1),
		767 => to_unsigned(2407, LUT_AMPL_WIDTH - 1),
		768 => to_unsigned(2410, LUT_AMPL_WIDTH - 1),
		769 => to_unsigned(2414, LUT_AMPL_WIDTH - 1),
		770 => to_unsigned(2417, LUT_AMPL_WIDTH - 1),
		771 => to_unsigned(2420, LUT_AMPL_WIDTH - 1),
		772 => to_unsigned(2423, LUT_AMPL_WIDTH - 1),
		773 => to_unsigned(2426, LUT_AMPL_WIDTH - 1),
		774 => to_unsigned(2429, LUT_AMPL_WIDTH - 1),
		775 => to_unsigned(2432, LUT_AMPL_WIDTH - 1),
		776 => to_unsigned(2436, LUT_AMPL_WIDTH - 1),
		777 => to_unsigned(2439, LUT_AMPL_WIDTH - 1),
		778 => to_unsigned(2442, LUT_AMPL_WIDTH - 1),
		779 => to_unsigned(2445, LUT_AMPL_WIDTH - 1),
		780 => to_unsigned(2448, LUT_AMPL_WIDTH - 1),
		781 => to_unsigned(2451, LUT_AMPL_WIDTH - 1),
		782 => to_unsigned(2454, LUT_AMPL_WIDTH - 1),
		783 => to_unsigned(2457, LUT_AMPL_WIDTH - 1),
		784 => to_unsigned(2461, LUT_AMPL_WIDTH - 1),
		785 => to_unsigned(2464, LUT_AMPL_WIDTH - 1),
		786 => to_unsigned(2467, LUT_AMPL_WIDTH - 1),
		787 => to_unsigned(2470, LUT_AMPL_WIDTH - 1),
		788 => to_unsigned(2473, LUT_AMPL_WIDTH - 1),
		789 => to_unsigned(2476, LUT_AMPL_WIDTH - 1),
		790 => to_unsigned(2479, LUT_AMPL_WIDTH - 1),
		791 => to_unsigned(2483, LUT_AMPL_WIDTH - 1),
		792 => to_unsigned(2486, LUT_AMPL_WIDTH - 1),
		793 => to_unsigned(2489, LUT_AMPL_WIDTH - 1),
		794 => to_unsigned(2492, LUT_AMPL_WIDTH - 1),
		795 => to_unsigned(2495, LUT_AMPL_WIDTH - 1),
		796 => to_unsigned(2498, LUT_AMPL_WIDTH - 1),
		797 => to_unsigned(2501, LUT_AMPL_WIDTH - 1),
		798 => to_unsigned(2504, LUT_AMPL_WIDTH - 1),
		799 => to_unsigned(2508, LUT_AMPL_WIDTH - 1),
		800 => to_unsigned(2511, LUT_AMPL_WIDTH - 1),
		801 => to_unsigned(2514, LUT_AMPL_WIDTH - 1),
		802 => to_unsigned(2517, LUT_AMPL_WIDTH - 1),
		803 => to_unsigned(2520, LUT_AMPL_WIDTH - 1),
		804 => to_unsigned(2523, LUT_AMPL_WIDTH - 1),
		805 => to_unsigned(2526, LUT_AMPL_WIDTH - 1),
		806 => to_unsigned(2530, LUT_AMPL_WIDTH - 1),
		807 => to_unsigned(2533, LUT_AMPL_WIDTH - 1),
		808 => to_unsigned(2536, LUT_AMPL_WIDTH - 1),
		809 => to_unsigned(2539, LUT_AMPL_WIDTH - 1),
		810 => to_unsigned(2542, LUT_AMPL_WIDTH - 1),
		811 => to_unsigned(2545, LUT_AMPL_WIDTH - 1),
		812 => to_unsigned(2548, LUT_AMPL_WIDTH - 1),
		813 => to_unsigned(2551, LUT_AMPL_WIDTH - 1),
		814 => to_unsigned(2555, LUT_AMPL_WIDTH - 1),
		815 => to_unsigned(2558, LUT_AMPL_WIDTH - 1),
		816 => to_unsigned(2561, LUT_AMPL_WIDTH - 1),
		817 => to_unsigned(2564, LUT_AMPL_WIDTH - 1),
		818 => to_unsigned(2567, LUT_AMPL_WIDTH - 1),
		819 => to_unsigned(2570, LUT_AMPL_WIDTH - 1),
		820 => to_unsigned(2573, LUT_AMPL_WIDTH - 1),
		821 => to_unsigned(2577, LUT_AMPL_WIDTH - 1),
		822 => to_unsigned(2580, LUT_AMPL_WIDTH - 1),
		823 => to_unsigned(2583, LUT_AMPL_WIDTH - 1),
		824 => to_unsigned(2586, LUT_AMPL_WIDTH - 1),
		825 => to_unsigned(2589, LUT_AMPL_WIDTH - 1),
		826 => to_unsigned(2592, LUT_AMPL_WIDTH - 1),
		827 => to_unsigned(2595, LUT_AMPL_WIDTH - 1),
		828 => to_unsigned(2598, LUT_AMPL_WIDTH - 1),
		829 => to_unsigned(2602, LUT_AMPL_WIDTH - 1),
		830 => to_unsigned(2605, LUT_AMPL_WIDTH - 1),
		831 => to_unsigned(2608, LUT_AMPL_WIDTH - 1),
		832 => to_unsigned(2611, LUT_AMPL_WIDTH - 1),
		833 => to_unsigned(2614, LUT_AMPL_WIDTH - 1),
		834 => to_unsigned(2617, LUT_AMPL_WIDTH - 1),
		835 => to_unsigned(2620, LUT_AMPL_WIDTH - 1),
		836 => to_unsigned(2623, LUT_AMPL_WIDTH - 1),
		837 => to_unsigned(2627, LUT_AMPL_WIDTH - 1),
		838 => to_unsigned(2630, LUT_AMPL_WIDTH - 1),
		839 => to_unsigned(2633, LUT_AMPL_WIDTH - 1),
		840 => to_unsigned(2636, LUT_AMPL_WIDTH - 1),
		841 => to_unsigned(2639, LUT_AMPL_WIDTH - 1),
		842 => to_unsigned(2642, LUT_AMPL_WIDTH - 1),
		843 => to_unsigned(2645, LUT_AMPL_WIDTH - 1),
		844 => to_unsigned(2649, LUT_AMPL_WIDTH - 1),
		845 => to_unsigned(2652, LUT_AMPL_WIDTH - 1),
		846 => to_unsigned(2655, LUT_AMPL_WIDTH - 1),
		847 => to_unsigned(2658, LUT_AMPL_WIDTH - 1),
		848 => to_unsigned(2661, LUT_AMPL_WIDTH - 1),
		849 => to_unsigned(2664, LUT_AMPL_WIDTH - 1),
		850 => to_unsigned(2667, LUT_AMPL_WIDTH - 1),
		851 => to_unsigned(2670, LUT_AMPL_WIDTH - 1),
		852 => to_unsigned(2674, LUT_AMPL_WIDTH - 1),
		853 => to_unsigned(2677, LUT_AMPL_WIDTH - 1),
		854 => to_unsigned(2680, LUT_AMPL_WIDTH - 1),
		855 => to_unsigned(2683, LUT_AMPL_WIDTH - 1),
		856 => to_unsigned(2686, LUT_AMPL_WIDTH - 1),
		857 => to_unsigned(2689, LUT_AMPL_WIDTH - 1),
		858 => to_unsigned(2692, LUT_AMPL_WIDTH - 1),
		859 => to_unsigned(2695, LUT_AMPL_WIDTH - 1),
		860 => to_unsigned(2699, LUT_AMPL_WIDTH - 1),
		861 => to_unsigned(2702, LUT_AMPL_WIDTH - 1),
		862 => to_unsigned(2705, LUT_AMPL_WIDTH - 1),
		863 => to_unsigned(2708, LUT_AMPL_WIDTH - 1),
		864 => to_unsigned(2711, LUT_AMPL_WIDTH - 1),
		865 => to_unsigned(2714, LUT_AMPL_WIDTH - 1),
		866 => to_unsigned(2717, LUT_AMPL_WIDTH - 1),
		867 => to_unsigned(2721, LUT_AMPL_WIDTH - 1),
		868 => to_unsigned(2724, LUT_AMPL_WIDTH - 1),
		869 => to_unsigned(2727, LUT_AMPL_WIDTH - 1),
		870 => to_unsigned(2730, LUT_AMPL_WIDTH - 1),
		871 => to_unsigned(2733, LUT_AMPL_WIDTH - 1),
		872 => to_unsigned(2736, LUT_AMPL_WIDTH - 1),
		873 => to_unsigned(2739, LUT_AMPL_WIDTH - 1),
		874 => to_unsigned(2742, LUT_AMPL_WIDTH - 1),
		875 => to_unsigned(2746, LUT_AMPL_WIDTH - 1),
		876 => to_unsigned(2749, LUT_AMPL_WIDTH - 1),
		877 => to_unsigned(2752, LUT_AMPL_WIDTH - 1),
		878 => to_unsigned(2755, LUT_AMPL_WIDTH - 1),
		879 => to_unsigned(2758, LUT_AMPL_WIDTH - 1),
		880 => to_unsigned(2761, LUT_AMPL_WIDTH - 1),
		881 => to_unsigned(2764, LUT_AMPL_WIDTH - 1),
		882 => to_unsigned(2767, LUT_AMPL_WIDTH - 1),
		883 => to_unsigned(2771, LUT_AMPL_WIDTH - 1),
		884 => to_unsigned(2774, LUT_AMPL_WIDTH - 1),
		885 => to_unsigned(2777, LUT_AMPL_WIDTH - 1),
		886 => to_unsigned(2780, LUT_AMPL_WIDTH - 1),
		887 => to_unsigned(2783, LUT_AMPL_WIDTH - 1),
		888 => to_unsigned(2786, LUT_AMPL_WIDTH - 1),
		889 => to_unsigned(2789, LUT_AMPL_WIDTH - 1),
		890 => to_unsigned(2793, LUT_AMPL_WIDTH - 1),
		891 => to_unsigned(2796, LUT_AMPL_WIDTH - 1),
		892 => to_unsigned(2799, LUT_AMPL_WIDTH - 1),
		893 => to_unsigned(2802, LUT_AMPL_WIDTH - 1),
		894 => to_unsigned(2805, LUT_AMPL_WIDTH - 1),
		895 => to_unsigned(2808, LUT_AMPL_WIDTH - 1),
		896 => to_unsigned(2811, LUT_AMPL_WIDTH - 1),
		897 => to_unsigned(2814, LUT_AMPL_WIDTH - 1),
		898 => to_unsigned(2818, LUT_AMPL_WIDTH - 1),
		899 => to_unsigned(2821, LUT_AMPL_WIDTH - 1),
		900 => to_unsigned(2824, LUT_AMPL_WIDTH - 1),
		901 => to_unsigned(2827, LUT_AMPL_WIDTH - 1),
		902 => to_unsigned(2830, LUT_AMPL_WIDTH - 1),
		903 => to_unsigned(2833, LUT_AMPL_WIDTH - 1),
		904 => to_unsigned(2836, LUT_AMPL_WIDTH - 1),
		905 => to_unsigned(2839, LUT_AMPL_WIDTH - 1),
		906 => to_unsigned(2843, LUT_AMPL_WIDTH - 1),
		907 => to_unsigned(2846, LUT_AMPL_WIDTH - 1),
		908 => to_unsigned(2849, LUT_AMPL_WIDTH - 1),
		909 => to_unsigned(2852, LUT_AMPL_WIDTH - 1),
		910 => to_unsigned(2855, LUT_AMPL_WIDTH - 1),
		911 => to_unsigned(2858, LUT_AMPL_WIDTH - 1),
		912 => to_unsigned(2861, LUT_AMPL_WIDTH - 1),
		913 => to_unsigned(2865, LUT_AMPL_WIDTH - 1),
		914 => to_unsigned(2868, LUT_AMPL_WIDTH - 1),
		915 => to_unsigned(2871, LUT_AMPL_WIDTH - 1),
		916 => to_unsigned(2874, LUT_AMPL_WIDTH - 1),
		917 => to_unsigned(2877, LUT_AMPL_WIDTH - 1),
		918 => to_unsigned(2880, LUT_AMPL_WIDTH - 1),
		919 => to_unsigned(2883, LUT_AMPL_WIDTH - 1),
		920 => to_unsigned(2886, LUT_AMPL_WIDTH - 1),
		921 => to_unsigned(2890, LUT_AMPL_WIDTH - 1),
		922 => to_unsigned(2893, LUT_AMPL_WIDTH - 1),
		923 => to_unsigned(2896, LUT_AMPL_WIDTH - 1),
		924 => to_unsigned(2899, LUT_AMPL_WIDTH - 1),
		925 => to_unsigned(2902, LUT_AMPL_WIDTH - 1),
		926 => to_unsigned(2905, LUT_AMPL_WIDTH - 1),
		927 => to_unsigned(2908, LUT_AMPL_WIDTH - 1),
		928 => to_unsigned(2911, LUT_AMPL_WIDTH - 1),
		929 => to_unsigned(2915, LUT_AMPL_WIDTH - 1),
		930 => to_unsigned(2918, LUT_AMPL_WIDTH - 1),
		931 => to_unsigned(2921, LUT_AMPL_WIDTH - 1),
		932 => to_unsigned(2924, LUT_AMPL_WIDTH - 1),
		933 => to_unsigned(2927, LUT_AMPL_WIDTH - 1),
		934 => to_unsigned(2930, LUT_AMPL_WIDTH - 1),
		935 => to_unsigned(2933, LUT_AMPL_WIDTH - 1),
		936 => to_unsigned(2936, LUT_AMPL_WIDTH - 1),
		937 => to_unsigned(2940, LUT_AMPL_WIDTH - 1),
		938 => to_unsigned(2943, LUT_AMPL_WIDTH - 1),
		939 => to_unsigned(2946, LUT_AMPL_WIDTH - 1),
		940 => to_unsigned(2949, LUT_AMPL_WIDTH - 1),
		941 => to_unsigned(2952, LUT_AMPL_WIDTH - 1),
		942 => to_unsigned(2955, LUT_AMPL_WIDTH - 1),
		943 => to_unsigned(2958, LUT_AMPL_WIDTH - 1),
		944 => to_unsigned(2962, LUT_AMPL_WIDTH - 1),
		945 => to_unsigned(2965, LUT_AMPL_WIDTH - 1),
		946 => to_unsigned(2968, LUT_AMPL_WIDTH - 1),
		947 => to_unsigned(2971, LUT_AMPL_WIDTH - 1),
		948 => to_unsigned(2974, LUT_AMPL_WIDTH - 1),
		949 => to_unsigned(2977, LUT_AMPL_WIDTH - 1),
		950 => to_unsigned(2980, LUT_AMPL_WIDTH - 1),
		951 => to_unsigned(2983, LUT_AMPL_WIDTH - 1),
		952 => to_unsigned(2987, LUT_AMPL_WIDTH - 1),
		953 => to_unsigned(2990, LUT_AMPL_WIDTH - 1),
		954 => to_unsigned(2993, LUT_AMPL_WIDTH - 1),
		955 => to_unsigned(2996, LUT_AMPL_WIDTH - 1),
		956 => to_unsigned(2999, LUT_AMPL_WIDTH - 1),
		957 => to_unsigned(3002, LUT_AMPL_WIDTH - 1),
		958 => to_unsigned(3005, LUT_AMPL_WIDTH - 1),
		959 => to_unsigned(3008, LUT_AMPL_WIDTH - 1),
		960 => to_unsigned(3012, LUT_AMPL_WIDTH - 1),
		961 => to_unsigned(3015, LUT_AMPL_WIDTH - 1),
		962 => to_unsigned(3018, LUT_AMPL_WIDTH - 1),
		963 => to_unsigned(3021, LUT_AMPL_WIDTH - 1),
		964 => to_unsigned(3024, LUT_AMPL_WIDTH - 1),
		965 => to_unsigned(3027, LUT_AMPL_WIDTH - 1),
		966 => to_unsigned(3030, LUT_AMPL_WIDTH - 1),
		967 => to_unsigned(3033, LUT_AMPL_WIDTH - 1),
		968 => to_unsigned(3037, LUT_AMPL_WIDTH - 1),
		969 => to_unsigned(3040, LUT_AMPL_WIDTH - 1),
		970 => to_unsigned(3043, LUT_AMPL_WIDTH - 1),
		971 => to_unsigned(3046, LUT_AMPL_WIDTH - 1),
		972 => to_unsigned(3049, LUT_AMPL_WIDTH - 1),
		973 => to_unsigned(3052, LUT_AMPL_WIDTH - 1),
		974 => to_unsigned(3055, LUT_AMPL_WIDTH - 1),
		975 => to_unsigned(3059, LUT_AMPL_WIDTH - 1),
		976 => to_unsigned(3062, LUT_AMPL_WIDTH - 1),
		977 => to_unsigned(3065, LUT_AMPL_WIDTH - 1),
		978 => to_unsigned(3068, LUT_AMPL_WIDTH - 1),
		979 => to_unsigned(3071, LUT_AMPL_WIDTH - 1),
		980 => to_unsigned(3074, LUT_AMPL_WIDTH - 1),
		981 => to_unsigned(3077, LUT_AMPL_WIDTH - 1),
		982 => to_unsigned(3080, LUT_AMPL_WIDTH - 1),
		983 => to_unsigned(3084, LUT_AMPL_WIDTH - 1),
		984 => to_unsigned(3087, LUT_AMPL_WIDTH - 1),
		985 => to_unsigned(3090, LUT_AMPL_WIDTH - 1),
		986 => to_unsigned(3093, LUT_AMPL_WIDTH - 1),
		987 => to_unsigned(3096, LUT_AMPL_WIDTH - 1),
		988 => to_unsigned(3099, LUT_AMPL_WIDTH - 1),
		989 => to_unsigned(3102, LUT_AMPL_WIDTH - 1),
		990 => to_unsigned(3105, LUT_AMPL_WIDTH - 1),
		991 => to_unsigned(3109, LUT_AMPL_WIDTH - 1),
		992 => to_unsigned(3112, LUT_AMPL_WIDTH - 1),
		993 => to_unsigned(3115, LUT_AMPL_WIDTH - 1),
		994 => to_unsigned(3118, LUT_AMPL_WIDTH - 1),
		995 => to_unsigned(3121, LUT_AMPL_WIDTH - 1),
		996 => to_unsigned(3124, LUT_AMPL_WIDTH - 1),
		997 => to_unsigned(3127, LUT_AMPL_WIDTH - 1),
		998 => to_unsigned(3130, LUT_AMPL_WIDTH - 1),
		999 => to_unsigned(3134, LUT_AMPL_WIDTH - 1),
		1000 => to_unsigned(3137, LUT_AMPL_WIDTH - 1),
		1001 => to_unsigned(3140, LUT_AMPL_WIDTH - 1),
		1002 => to_unsigned(3143, LUT_AMPL_WIDTH - 1),
		1003 => to_unsigned(3146, LUT_AMPL_WIDTH - 1),
		1004 => to_unsigned(3149, LUT_AMPL_WIDTH - 1),
		1005 => to_unsigned(3152, LUT_AMPL_WIDTH - 1),
		1006 => to_unsigned(3155, LUT_AMPL_WIDTH - 1),
		1007 => to_unsigned(3159, LUT_AMPL_WIDTH - 1),
		1008 => to_unsigned(3162, LUT_AMPL_WIDTH - 1),
		1009 => to_unsigned(3165, LUT_AMPL_WIDTH - 1),
		1010 => to_unsigned(3168, LUT_AMPL_WIDTH - 1),
		1011 => to_unsigned(3171, LUT_AMPL_WIDTH - 1),
		1012 => to_unsigned(3174, LUT_AMPL_WIDTH - 1),
		1013 => to_unsigned(3177, LUT_AMPL_WIDTH - 1),
		1014 => to_unsigned(3180, LUT_AMPL_WIDTH - 1),
		1015 => to_unsigned(3184, LUT_AMPL_WIDTH - 1),
		1016 => to_unsigned(3187, LUT_AMPL_WIDTH - 1),
		1017 => to_unsigned(3190, LUT_AMPL_WIDTH - 1),
		1018 => to_unsigned(3193, LUT_AMPL_WIDTH - 1),
		1019 => to_unsigned(3196, LUT_AMPL_WIDTH - 1),
		1020 => to_unsigned(3199, LUT_AMPL_WIDTH - 1),
		1021 => to_unsigned(3202, LUT_AMPL_WIDTH - 1),
		1022 => to_unsigned(3205, LUT_AMPL_WIDTH - 1),
		1023 => to_unsigned(3209, LUT_AMPL_WIDTH - 1),
		1024 => to_unsigned(3212, LUT_AMPL_WIDTH - 1),
		1025 => to_unsigned(3215, LUT_AMPL_WIDTH - 1),
		1026 => to_unsigned(3218, LUT_AMPL_WIDTH - 1),
		1027 => to_unsigned(3221, LUT_AMPL_WIDTH - 1),
		1028 => to_unsigned(3224, LUT_AMPL_WIDTH - 1),
		1029 => to_unsigned(3227, LUT_AMPL_WIDTH - 1),
		1030 => to_unsigned(3230, LUT_AMPL_WIDTH - 1),
		1031 => to_unsigned(3234, LUT_AMPL_WIDTH - 1),
		1032 => to_unsigned(3237, LUT_AMPL_WIDTH - 1),
		1033 => to_unsigned(3240, LUT_AMPL_WIDTH - 1),
		1034 => to_unsigned(3243, LUT_AMPL_WIDTH - 1),
		1035 => to_unsigned(3246, LUT_AMPL_WIDTH - 1),
		1036 => to_unsigned(3249, LUT_AMPL_WIDTH - 1),
		1037 => to_unsigned(3252, LUT_AMPL_WIDTH - 1),
		1038 => to_unsigned(3255, LUT_AMPL_WIDTH - 1),
		1039 => to_unsigned(3259, LUT_AMPL_WIDTH - 1),
		1040 => to_unsigned(3262, LUT_AMPL_WIDTH - 1),
		1041 => to_unsigned(3265, LUT_AMPL_WIDTH - 1),
		1042 => to_unsigned(3268, LUT_AMPL_WIDTH - 1),
		1043 => to_unsigned(3271, LUT_AMPL_WIDTH - 1),
		1044 => to_unsigned(3274, LUT_AMPL_WIDTH - 1),
		1045 => to_unsigned(3277, LUT_AMPL_WIDTH - 1),
		1046 => to_unsigned(3281, LUT_AMPL_WIDTH - 1),
		1047 => to_unsigned(3284, LUT_AMPL_WIDTH - 1),
		1048 => to_unsigned(3287, LUT_AMPL_WIDTH - 1),
		1049 => to_unsigned(3290, LUT_AMPL_WIDTH - 1),
		1050 => to_unsigned(3293, LUT_AMPL_WIDTH - 1),
		1051 => to_unsigned(3296, LUT_AMPL_WIDTH - 1),
		1052 => to_unsigned(3299, LUT_AMPL_WIDTH - 1),
		1053 => to_unsigned(3302, LUT_AMPL_WIDTH - 1),
		1054 => to_unsigned(3306, LUT_AMPL_WIDTH - 1),
		1055 => to_unsigned(3309, LUT_AMPL_WIDTH - 1),
		1056 => to_unsigned(3312, LUT_AMPL_WIDTH - 1),
		1057 => to_unsigned(3315, LUT_AMPL_WIDTH - 1),
		1058 => to_unsigned(3318, LUT_AMPL_WIDTH - 1),
		1059 => to_unsigned(3321, LUT_AMPL_WIDTH - 1),
		1060 => to_unsigned(3324, LUT_AMPL_WIDTH - 1),
		1061 => to_unsigned(3327, LUT_AMPL_WIDTH - 1),
		1062 => to_unsigned(3331, LUT_AMPL_WIDTH - 1),
		1063 => to_unsigned(3334, LUT_AMPL_WIDTH - 1),
		1064 => to_unsigned(3337, LUT_AMPL_WIDTH - 1),
		1065 => to_unsigned(3340, LUT_AMPL_WIDTH - 1),
		1066 => to_unsigned(3343, LUT_AMPL_WIDTH - 1),
		1067 => to_unsigned(3346, LUT_AMPL_WIDTH - 1),
		1068 => to_unsigned(3349, LUT_AMPL_WIDTH - 1),
		1069 => to_unsigned(3352, LUT_AMPL_WIDTH - 1),
		1070 => to_unsigned(3356, LUT_AMPL_WIDTH - 1),
		1071 => to_unsigned(3359, LUT_AMPL_WIDTH - 1),
		1072 => to_unsigned(3362, LUT_AMPL_WIDTH - 1),
		1073 => to_unsigned(3365, LUT_AMPL_WIDTH - 1),
		1074 => to_unsigned(3368, LUT_AMPL_WIDTH - 1),
		1075 => to_unsigned(3371, LUT_AMPL_WIDTH - 1),
		1076 => to_unsigned(3374, LUT_AMPL_WIDTH - 1),
		1077 => to_unsigned(3377, LUT_AMPL_WIDTH - 1),
		1078 => to_unsigned(3381, LUT_AMPL_WIDTH - 1),
		1079 => to_unsigned(3384, LUT_AMPL_WIDTH - 1),
		1080 => to_unsigned(3387, LUT_AMPL_WIDTH - 1),
		1081 => to_unsigned(3390, LUT_AMPL_WIDTH - 1),
		1082 => to_unsigned(3393, LUT_AMPL_WIDTH - 1),
		1083 => to_unsigned(3396, LUT_AMPL_WIDTH - 1),
		1084 => to_unsigned(3399, LUT_AMPL_WIDTH - 1),
		1085 => to_unsigned(3402, LUT_AMPL_WIDTH - 1),
		1086 => to_unsigned(3406, LUT_AMPL_WIDTH - 1),
		1087 => to_unsigned(3409, LUT_AMPL_WIDTH - 1),
		1088 => to_unsigned(3412, LUT_AMPL_WIDTH - 1),
		1089 => to_unsigned(3415, LUT_AMPL_WIDTH - 1),
		1090 => to_unsigned(3418, LUT_AMPL_WIDTH - 1),
		1091 => to_unsigned(3421, LUT_AMPL_WIDTH - 1),
		1092 => to_unsigned(3424, LUT_AMPL_WIDTH - 1),
		1093 => to_unsigned(3427, LUT_AMPL_WIDTH - 1),
		1094 => to_unsigned(3430, LUT_AMPL_WIDTH - 1),
		1095 => to_unsigned(3434, LUT_AMPL_WIDTH - 1),
		1096 => to_unsigned(3437, LUT_AMPL_WIDTH - 1),
		1097 => to_unsigned(3440, LUT_AMPL_WIDTH - 1),
		1098 => to_unsigned(3443, LUT_AMPL_WIDTH - 1),
		1099 => to_unsigned(3446, LUT_AMPL_WIDTH - 1),
		1100 => to_unsigned(3449, LUT_AMPL_WIDTH - 1),
		1101 => to_unsigned(3452, LUT_AMPL_WIDTH - 1),
		1102 => to_unsigned(3455, LUT_AMPL_WIDTH - 1),
		1103 => to_unsigned(3459, LUT_AMPL_WIDTH - 1),
		1104 => to_unsigned(3462, LUT_AMPL_WIDTH - 1),
		1105 => to_unsigned(3465, LUT_AMPL_WIDTH - 1),
		1106 => to_unsigned(3468, LUT_AMPL_WIDTH - 1),
		1107 => to_unsigned(3471, LUT_AMPL_WIDTH - 1),
		1108 => to_unsigned(3474, LUT_AMPL_WIDTH - 1),
		1109 => to_unsigned(3477, LUT_AMPL_WIDTH - 1),
		1110 => to_unsigned(3480, LUT_AMPL_WIDTH - 1),
		1111 => to_unsigned(3484, LUT_AMPL_WIDTH - 1),
		1112 => to_unsigned(3487, LUT_AMPL_WIDTH - 1),
		1113 => to_unsigned(3490, LUT_AMPL_WIDTH - 1),
		1114 => to_unsigned(3493, LUT_AMPL_WIDTH - 1),
		1115 => to_unsigned(3496, LUT_AMPL_WIDTH - 1),
		1116 => to_unsigned(3499, LUT_AMPL_WIDTH - 1),
		1117 => to_unsigned(3502, LUT_AMPL_WIDTH - 1),
		1118 => to_unsigned(3505, LUT_AMPL_WIDTH - 1),
		1119 => to_unsigned(3509, LUT_AMPL_WIDTH - 1),
		1120 => to_unsigned(3512, LUT_AMPL_WIDTH - 1),
		1121 => to_unsigned(3515, LUT_AMPL_WIDTH - 1),
		1122 => to_unsigned(3518, LUT_AMPL_WIDTH - 1),
		1123 => to_unsigned(3521, LUT_AMPL_WIDTH - 1),
		1124 => to_unsigned(3524, LUT_AMPL_WIDTH - 1),
		1125 => to_unsigned(3527, LUT_AMPL_WIDTH - 1),
		1126 => to_unsigned(3530, LUT_AMPL_WIDTH - 1),
		1127 => to_unsigned(3534, LUT_AMPL_WIDTH - 1),
		1128 => to_unsigned(3537, LUT_AMPL_WIDTH - 1),
		1129 => to_unsigned(3540, LUT_AMPL_WIDTH - 1),
		1130 => to_unsigned(3543, LUT_AMPL_WIDTH - 1),
		1131 => to_unsigned(3546, LUT_AMPL_WIDTH - 1),
		1132 => to_unsigned(3549, LUT_AMPL_WIDTH - 1),
		1133 => to_unsigned(3552, LUT_AMPL_WIDTH - 1),
		1134 => to_unsigned(3555, LUT_AMPL_WIDTH - 1),
		1135 => to_unsigned(3559, LUT_AMPL_WIDTH - 1),
		1136 => to_unsigned(3562, LUT_AMPL_WIDTH - 1),
		1137 => to_unsigned(3565, LUT_AMPL_WIDTH - 1),
		1138 => to_unsigned(3568, LUT_AMPL_WIDTH - 1),
		1139 => to_unsigned(3571, LUT_AMPL_WIDTH - 1),
		1140 => to_unsigned(3574, LUT_AMPL_WIDTH - 1),
		1141 => to_unsigned(3577, LUT_AMPL_WIDTH - 1),
		1142 => to_unsigned(3580, LUT_AMPL_WIDTH - 1),
		1143 => to_unsigned(3584, LUT_AMPL_WIDTH - 1),
		1144 => to_unsigned(3587, LUT_AMPL_WIDTH - 1),
		1145 => to_unsigned(3590, LUT_AMPL_WIDTH - 1),
		1146 => to_unsigned(3593, LUT_AMPL_WIDTH - 1),
		1147 => to_unsigned(3596, LUT_AMPL_WIDTH - 1),
		1148 => to_unsigned(3599, LUT_AMPL_WIDTH - 1),
		1149 => to_unsigned(3602, LUT_AMPL_WIDTH - 1),
		1150 => to_unsigned(3605, LUT_AMPL_WIDTH - 1),
		1151 => to_unsigned(3609, LUT_AMPL_WIDTH - 1),
		1152 => to_unsigned(3612, LUT_AMPL_WIDTH - 1),
		1153 => to_unsigned(3615, LUT_AMPL_WIDTH - 1),
		1154 => to_unsigned(3618, LUT_AMPL_WIDTH - 1),
		1155 => to_unsigned(3621, LUT_AMPL_WIDTH - 1),
		1156 => to_unsigned(3624, LUT_AMPL_WIDTH - 1),
		1157 => to_unsigned(3627, LUT_AMPL_WIDTH - 1),
		1158 => to_unsigned(3630, LUT_AMPL_WIDTH - 1),
		1159 => to_unsigned(3634, LUT_AMPL_WIDTH - 1),
		1160 => to_unsigned(3637, LUT_AMPL_WIDTH - 1),
		1161 => to_unsigned(3640, LUT_AMPL_WIDTH - 1),
		1162 => to_unsigned(3643, LUT_AMPL_WIDTH - 1),
		1163 => to_unsigned(3646, LUT_AMPL_WIDTH - 1),
		1164 => to_unsigned(3649, LUT_AMPL_WIDTH - 1),
		1165 => to_unsigned(3652, LUT_AMPL_WIDTH - 1),
		1166 => to_unsigned(3655, LUT_AMPL_WIDTH - 1),
		1167 => to_unsigned(3658, LUT_AMPL_WIDTH - 1),
		1168 => to_unsigned(3662, LUT_AMPL_WIDTH - 1),
		1169 => to_unsigned(3665, LUT_AMPL_WIDTH - 1),
		1170 => to_unsigned(3668, LUT_AMPL_WIDTH - 1),
		1171 => to_unsigned(3671, LUT_AMPL_WIDTH - 1),
		1172 => to_unsigned(3674, LUT_AMPL_WIDTH - 1),
		1173 => to_unsigned(3677, LUT_AMPL_WIDTH - 1),
		1174 => to_unsigned(3680, LUT_AMPL_WIDTH - 1),
		1175 => to_unsigned(3683, LUT_AMPL_WIDTH - 1),
		1176 => to_unsigned(3687, LUT_AMPL_WIDTH - 1),
		1177 => to_unsigned(3690, LUT_AMPL_WIDTH - 1),
		1178 => to_unsigned(3693, LUT_AMPL_WIDTH - 1),
		1179 => to_unsigned(3696, LUT_AMPL_WIDTH - 1),
		1180 => to_unsigned(3699, LUT_AMPL_WIDTH - 1),
		1181 => to_unsigned(3702, LUT_AMPL_WIDTH - 1),
		1182 => to_unsigned(3705, LUT_AMPL_WIDTH - 1),
		1183 => to_unsigned(3708, LUT_AMPL_WIDTH - 1),
		1184 => to_unsigned(3712, LUT_AMPL_WIDTH - 1),
		1185 => to_unsigned(3715, LUT_AMPL_WIDTH - 1),
		1186 => to_unsigned(3718, LUT_AMPL_WIDTH - 1),
		1187 => to_unsigned(3721, LUT_AMPL_WIDTH - 1),
		1188 => to_unsigned(3724, LUT_AMPL_WIDTH - 1),
		1189 => to_unsigned(3727, LUT_AMPL_WIDTH - 1),
		1190 => to_unsigned(3730, LUT_AMPL_WIDTH - 1),
		1191 => to_unsigned(3733, LUT_AMPL_WIDTH - 1),
		1192 => to_unsigned(3737, LUT_AMPL_WIDTH - 1),
		1193 => to_unsigned(3740, LUT_AMPL_WIDTH - 1),
		1194 => to_unsigned(3743, LUT_AMPL_WIDTH - 1),
		1195 => to_unsigned(3746, LUT_AMPL_WIDTH - 1),
		1196 => to_unsigned(3749, LUT_AMPL_WIDTH - 1),
		1197 => to_unsigned(3752, LUT_AMPL_WIDTH - 1),
		1198 => to_unsigned(3755, LUT_AMPL_WIDTH - 1),
		1199 => to_unsigned(3758, LUT_AMPL_WIDTH - 1),
		1200 => to_unsigned(3761, LUT_AMPL_WIDTH - 1),
		1201 => to_unsigned(3765, LUT_AMPL_WIDTH - 1),
		1202 => to_unsigned(3768, LUT_AMPL_WIDTH - 1),
		1203 => to_unsigned(3771, LUT_AMPL_WIDTH - 1),
		1204 => to_unsigned(3774, LUT_AMPL_WIDTH - 1),
		1205 => to_unsigned(3777, LUT_AMPL_WIDTH - 1),
		1206 => to_unsigned(3780, LUT_AMPL_WIDTH - 1),
		1207 => to_unsigned(3783, LUT_AMPL_WIDTH - 1),
		1208 => to_unsigned(3786, LUT_AMPL_WIDTH - 1),
		1209 => to_unsigned(3790, LUT_AMPL_WIDTH - 1),
		1210 => to_unsigned(3793, LUT_AMPL_WIDTH - 1),
		1211 => to_unsigned(3796, LUT_AMPL_WIDTH - 1),
		1212 => to_unsigned(3799, LUT_AMPL_WIDTH - 1),
		1213 => to_unsigned(3802, LUT_AMPL_WIDTH - 1),
		1214 => to_unsigned(3805, LUT_AMPL_WIDTH - 1),
		1215 => to_unsigned(3808, LUT_AMPL_WIDTH - 1),
		1216 => to_unsigned(3811, LUT_AMPL_WIDTH - 1),
		1217 => to_unsigned(3815, LUT_AMPL_WIDTH - 1),
		1218 => to_unsigned(3818, LUT_AMPL_WIDTH - 1),
		1219 => to_unsigned(3821, LUT_AMPL_WIDTH - 1),
		1220 => to_unsigned(3824, LUT_AMPL_WIDTH - 1),
		1221 => to_unsigned(3827, LUT_AMPL_WIDTH - 1),
		1222 => to_unsigned(3830, LUT_AMPL_WIDTH - 1),
		1223 => to_unsigned(3833, LUT_AMPL_WIDTH - 1),
		1224 => to_unsigned(3836, LUT_AMPL_WIDTH - 1),
		1225 => to_unsigned(3839, LUT_AMPL_WIDTH - 1),
		1226 => to_unsigned(3843, LUT_AMPL_WIDTH - 1),
		1227 => to_unsigned(3846, LUT_AMPL_WIDTH - 1),
		1228 => to_unsigned(3849, LUT_AMPL_WIDTH - 1),
		1229 => to_unsigned(3852, LUT_AMPL_WIDTH - 1),
		1230 => to_unsigned(3855, LUT_AMPL_WIDTH - 1),
		1231 => to_unsigned(3858, LUT_AMPL_WIDTH - 1),
		1232 => to_unsigned(3861, LUT_AMPL_WIDTH - 1),
		1233 => to_unsigned(3864, LUT_AMPL_WIDTH - 1),
		1234 => to_unsigned(3868, LUT_AMPL_WIDTH - 1),
		1235 => to_unsigned(3871, LUT_AMPL_WIDTH - 1),
		1236 => to_unsigned(3874, LUT_AMPL_WIDTH - 1),
		1237 => to_unsigned(3877, LUT_AMPL_WIDTH - 1),
		1238 => to_unsigned(3880, LUT_AMPL_WIDTH - 1),
		1239 => to_unsigned(3883, LUT_AMPL_WIDTH - 1),
		1240 => to_unsigned(3886, LUT_AMPL_WIDTH - 1),
		1241 => to_unsigned(3889, LUT_AMPL_WIDTH - 1),
		1242 => to_unsigned(3893, LUT_AMPL_WIDTH - 1),
		1243 => to_unsigned(3896, LUT_AMPL_WIDTH - 1),
		1244 => to_unsigned(3899, LUT_AMPL_WIDTH - 1),
		1245 => to_unsigned(3902, LUT_AMPL_WIDTH - 1),
		1246 => to_unsigned(3905, LUT_AMPL_WIDTH - 1),
		1247 => to_unsigned(3908, LUT_AMPL_WIDTH - 1),
		1248 => to_unsigned(3911, LUT_AMPL_WIDTH - 1),
		1249 => to_unsigned(3914, LUT_AMPL_WIDTH - 1),
		1250 => to_unsigned(3917, LUT_AMPL_WIDTH - 1),
		1251 => to_unsigned(3921, LUT_AMPL_WIDTH - 1),
		1252 => to_unsigned(3924, LUT_AMPL_WIDTH - 1),
		1253 => to_unsigned(3927, LUT_AMPL_WIDTH - 1),
		1254 => to_unsigned(3930, LUT_AMPL_WIDTH - 1),
		1255 => to_unsigned(3933, LUT_AMPL_WIDTH - 1),
		1256 => to_unsigned(3936, LUT_AMPL_WIDTH - 1),
		1257 => to_unsigned(3939, LUT_AMPL_WIDTH - 1),
		1258 => to_unsigned(3942, LUT_AMPL_WIDTH - 1),
		1259 => to_unsigned(3946, LUT_AMPL_WIDTH - 1),
		1260 => to_unsigned(3949, LUT_AMPL_WIDTH - 1),
		1261 => to_unsigned(3952, LUT_AMPL_WIDTH - 1),
		1262 => to_unsigned(3955, LUT_AMPL_WIDTH - 1),
		1263 => to_unsigned(3958, LUT_AMPL_WIDTH - 1),
		1264 => to_unsigned(3961, LUT_AMPL_WIDTH - 1),
		1265 => to_unsigned(3964, LUT_AMPL_WIDTH - 1),
		1266 => to_unsigned(3967, LUT_AMPL_WIDTH - 1),
		1267 => to_unsigned(3970, LUT_AMPL_WIDTH - 1),
		1268 => to_unsigned(3974, LUT_AMPL_WIDTH - 1),
		1269 => to_unsigned(3977, LUT_AMPL_WIDTH - 1),
		1270 => to_unsigned(3980, LUT_AMPL_WIDTH - 1),
		1271 => to_unsigned(3983, LUT_AMPL_WIDTH - 1),
		1272 => to_unsigned(3986, LUT_AMPL_WIDTH - 1),
		1273 => to_unsigned(3989, LUT_AMPL_WIDTH - 1),
		1274 => to_unsigned(3992, LUT_AMPL_WIDTH - 1),
		1275 => to_unsigned(3995, LUT_AMPL_WIDTH - 1),
		1276 => to_unsigned(3999, LUT_AMPL_WIDTH - 1),
		1277 => to_unsigned(4002, LUT_AMPL_WIDTH - 1),
		1278 => to_unsigned(4005, LUT_AMPL_WIDTH - 1),
		1279 => to_unsigned(4008, LUT_AMPL_WIDTH - 1),
		1280 => to_unsigned(4011, LUT_AMPL_WIDTH - 1),
		1281 => to_unsigned(4014, LUT_AMPL_WIDTH - 1),
		1282 => to_unsigned(4017, LUT_AMPL_WIDTH - 1),
		1283 => to_unsigned(4020, LUT_AMPL_WIDTH - 1),
		1284 => to_unsigned(4024, LUT_AMPL_WIDTH - 1),
		1285 => to_unsigned(4027, LUT_AMPL_WIDTH - 1),
		1286 => to_unsigned(4030, LUT_AMPL_WIDTH - 1),
		1287 => to_unsigned(4033, LUT_AMPL_WIDTH - 1),
		1288 => to_unsigned(4036, LUT_AMPL_WIDTH - 1),
		1289 => to_unsigned(4039, LUT_AMPL_WIDTH - 1),
		1290 => to_unsigned(4042, LUT_AMPL_WIDTH - 1),
		1291 => to_unsigned(4045, LUT_AMPL_WIDTH - 1),
		1292 => to_unsigned(4048, LUT_AMPL_WIDTH - 1),
		1293 => to_unsigned(4052, LUT_AMPL_WIDTH - 1),
		1294 => to_unsigned(4055, LUT_AMPL_WIDTH - 1),
		1295 => to_unsigned(4058, LUT_AMPL_WIDTH - 1),
		1296 => to_unsigned(4061, LUT_AMPL_WIDTH - 1),
		1297 => to_unsigned(4064, LUT_AMPL_WIDTH - 1),
		1298 => to_unsigned(4067, LUT_AMPL_WIDTH - 1),
		1299 => to_unsigned(4070, LUT_AMPL_WIDTH - 1),
		1300 => to_unsigned(4073, LUT_AMPL_WIDTH - 1),
		1301 => to_unsigned(4076, LUT_AMPL_WIDTH - 1),
		1302 => to_unsigned(4080, LUT_AMPL_WIDTH - 1),
		1303 => to_unsigned(4083, LUT_AMPL_WIDTH - 1),
		1304 => to_unsigned(4086, LUT_AMPL_WIDTH - 1),
		1305 => to_unsigned(4089, LUT_AMPL_WIDTH - 1),
		1306 => to_unsigned(4092, LUT_AMPL_WIDTH - 1),
		1307 => to_unsigned(4095, LUT_AMPL_WIDTH - 1),
		1308 => to_unsigned(4098, LUT_AMPL_WIDTH - 1),
		1309 => to_unsigned(4101, LUT_AMPL_WIDTH - 1),
		1310 => to_unsigned(4105, LUT_AMPL_WIDTH - 1),
		1311 => to_unsigned(4108, LUT_AMPL_WIDTH - 1),
		1312 => to_unsigned(4111, LUT_AMPL_WIDTH - 1),
		1313 => to_unsigned(4114, LUT_AMPL_WIDTH - 1),
		1314 => to_unsigned(4117, LUT_AMPL_WIDTH - 1),
		1315 => to_unsigned(4120, LUT_AMPL_WIDTH - 1),
		1316 => to_unsigned(4123, LUT_AMPL_WIDTH - 1),
		1317 => to_unsigned(4126, LUT_AMPL_WIDTH - 1),
		1318 => to_unsigned(4129, LUT_AMPL_WIDTH - 1),
		1319 => to_unsigned(4133, LUT_AMPL_WIDTH - 1),
		1320 => to_unsigned(4136, LUT_AMPL_WIDTH - 1),
		1321 => to_unsigned(4139, LUT_AMPL_WIDTH - 1),
		1322 => to_unsigned(4142, LUT_AMPL_WIDTH - 1),
		1323 => to_unsigned(4145, LUT_AMPL_WIDTH - 1),
		1324 => to_unsigned(4148, LUT_AMPL_WIDTH - 1),
		1325 => to_unsigned(4151, LUT_AMPL_WIDTH - 1),
		1326 => to_unsigned(4154, LUT_AMPL_WIDTH - 1),
		1327 => to_unsigned(4158, LUT_AMPL_WIDTH - 1),
		1328 => to_unsigned(4161, LUT_AMPL_WIDTH - 1),
		1329 => to_unsigned(4164, LUT_AMPL_WIDTH - 1),
		1330 => to_unsigned(4167, LUT_AMPL_WIDTH - 1),
		1331 => to_unsigned(4170, LUT_AMPL_WIDTH - 1),
		1332 => to_unsigned(4173, LUT_AMPL_WIDTH - 1),
		1333 => to_unsigned(4176, LUT_AMPL_WIDTH - 1),
		1334 => to_unsigned(4179, LUT_AMPL_WIDTH - 1),
		1335 => to_unsigned(4182, LUT_AMPL_WIDTH - 1),
		1336 => to_unsigned(4186, LUT_AMPL_WIDTH - 1),
		1337 => to_unsigned(4189, LUT_AMPL_WIDTH - 1),
		1338 => to_unsigned(4192, LUT_AMPL_WIDTH - 1),
		1339 => to_unsigned(4195, LUT_AMPL_WIDTH - 1),
		1340 => to_unsigned(4198, LUT_AMPL_WIDTH - 1),
		1341 => to_unsigned(4201, LUT_AMPL_WIDTH - 1),
		1342 => to_unsigned(4204, LUT_AMPL_WIDTH - 1),
		1343 => to_unsigned(4207, LUT_AMPL_WIDTH - 1),
		1344 => to_unsigned(4210, LUT_AMPL_WIDTH - 1),
		1345 => to_unsigned(4214, LUT_AMPL_WIDTH - 1),
		1346 => to_unsigned(4217, LUT_AMPL_WIDTH - 1),
		1347 => to_unsigned(4220, LUT_AMPL_WIDTH - 1),
		1348 => to_unsigned(4223, LUT_AMPL_WIDTH - 1),
		1349 => to_unsigned(4226, LUT_AMPL_WIDTH - 1),
		1350 => to_unsigned(4229, LUT_AMPL_WIDTH - 1),
		1351 => to_unsigned(4232, LUT_AMPL_WIDTH - 1),
		1352 => to_unsigned(4235, LUT_AMPL_WIDTH - 1),
		1353 => to_unsigned(4239, LUT_AMPL_WIDTH - 1),
		1354 => to_unsigned(4242, LUT_AMPL_WIDTH - 1),
		1355 => to_unsigned(4245, LUT_AMPL_WIDTH - 1),
		1356 => to_unsigned(4248, LUT_AMPL_WIDTH - 1),
		1357 => to_unsigned(4251, LUT_AMPL_WIDTH - 1),
		1358 => to_unsigned(4254, LUT_AMPL_WIDTH - 1),
		1359 => to_unsigned(4257, LUT_AMPL_WIDTH - 1),
		1360 => to_unsigned(4260, LUT_AMPL_WIDTH - 1),
		1361 => to_unsigned(4263, LUT_AMPL_WIDTH - 1),
		1362 => to_unsigned(4267, LUT_AMPL_WIDTH - 1),
		1363 => to_unsigned(4270, LUT_AMPL_WIDTH - 1),
		1364 => to_unsigned(4273, LUT_AMPL_WIDTH - 1),
		1365 => to_unsigned(4276, LUT_AMPL_WIDTH - 1),
		1366 => to_unsigned(4279, LUT_AMPL_WIDTH - 1),
		1367 => to_unsigned(4282, LUT_AMPL_WIDTH - 1),
		1368 => to_unsigned(4285, LUT_AMPL_WIDTH - 1),
		1369 => to_unsigned(4288, LUT_AMPL_WIDTH - 1),
		1370 => to_unsigned(4291, LUT_AMPL_WIDTH - 1),
		1371 => to_unsigned(4295, LUT_AMPL_WIDTH - 1),
		1372 => to_unsigned(4298, LUT_AMPL_WIDTH - 1),
		1373 => to_unsigned(4301, LUT_AMPL_WIDTH - 1),
		1374 => to_unsigned(4304, LUT_AMPL_WIDTH - 1),
		1375 => to_unsigned(4307, LUT_AMPL_WIDTH - 1),
		1376 => to_unsigned(4310, LUT_AMPL_WIDTH - 1),
		1377 => to_unsigned(4313, LUT_AMPL_WIDTH - 1),
		1378 => to_unsigned(4316, LUT_AMPL_WIDTH - 1),
		1379 => to_unsigned(4320, LUT_AMPL_WIDTH - 1),
		1380 => to_unsigned(4323, LUT_AMPL_WIDTH - 1),
		1381 => to_unsigned(4326, LUT_AMPL_WIDTH - 1),
		1382 => to_unsigned(4329, LUT_AMPL_WIDTH - 1),
		1383 => to_unsigned(4332, LUT_AMPL_WIDTH - 1),
		1384 => to_unsigned(4335, LUT_AMPL_WIDTH - 1),
		1385 => to_unsigned(4338, LUT_AMPL_WIDTH - 1),
		1386 => to_unsigned(4341, LUT_AMPL_WIDTH - 1),
		1387 => to_unsigned(4344, LUT_AMPL_WIDTH - 1),
		1388 => to_unsigned(4348, LUT_AMPL_WIDTH - 1),
		1389 => to_unsigned(4351, LUT_AMPL_WIDTH - 1),
		1390 => to_unsigned(4354, LUT_AMPL_WIDTH - 1),
		1391 => to_unsigned(4357, LUT_AMPL_WIDTH - 1),
		1392 => to_unsigned(4360, LUT_AMPL_WIDTH - 1),
		1393 => to_unsigned(4363, LUT_AMPL_WIDTH - 1),
		1394 => to_unsigned(4366, LUT_AMPL_WIDTH - 1),
		1395 => to_unsigned(4369, LUT_AMPL_WIDTH - 1),
		1396 => to_unsigned(4372, LUT_AMPL_WIDTH - 1),
		1397 => to_unsigned(4376, LUT_AMPL_WIDTH - 1),
		1398 => to_unsigned(4379, LUT_AMPL_WIDTH - 1),
		1399 => to_unsigned(4382, LUT_AMPL_WIDTH - 1),
		1400 => to_unsigned(4385, LUT_AMPL_WIDTH - 1),
		1401 => to_unsigned(4388, LUT_AMPL_WIDTH - 1),
		1402 => to_unsigned(4391, LUT_AMPL_WIDTH - 1),
		1403 => to_unsigned(4394, LUT_AMPL_WIDTH - 1),
		1404 => to_unsigned(4397, LUT_AMPL_WIDTH - 1),
		1405 => to_unsigned(4400, LUT_AMPL_WIDTH - 1),
		1406 => to_unsigned(4404, LUT_AMPL_WIDTH - 1),
		1407 => to_unsigned(4407, LUT_AMPL_WIDTH - 1),
		1408 => to_unsigned(4410, LUT_AMPL_WIDTH - 1),
		1409 => to_unsigned(4413, LUT_AMPL_WIDTH - 1),
		1410 => to_unsigned(4416, LUT_AMPL_WIDTH - 1),
		1411 => to_unsigned(4419, LUT_AMPL_WIDTH - 1),
		1412 => to_unsigned(4422, LUT_AMPL_WIDTH - 1),
		1413 => to_unsigned(4425, LUT_AMPL_WIDTH - 1),
		1414 => to_unsigned(4428, LUT_AMPL_WIDTH - 1),
		1415 => to_unsigned(4432, LUT_AMPL_WIDTH - 1),
		1416 => to_unsigned(4435, LUT_AMPL_WIDTH - 1),
		1417 => to_unsigned(4438, LUT_AMPL_WIDTH - 1),
		1418 => to_unsigned(4441, LUT_AMPL_WIDTH - 1),
		1419 => to_unsigned(4444, LUT_AMPL_WIDTH - 1),
		1420 => to_unsigned(4447, LUT_AMPL_WIDTH - 1),
		1421 => to_unsigned(4450, LUT_AMPL_WIDTH - 1),
		1422 => to_unsigned(4453, LUT_AMPL_WIDTH - 1),
		1423 => to_unsigned(4456, LUT_AMPL_WIDTH - 1),
		1424 => to_unsigned(4460, LUT_AMPL_WIDTH - 1),
		1425 => to_unsigned(4463, LUT_AMPL_WIDTH - 1),
		1426 => to_unsigned(4466, LUT_AMPL_WIDTH - 1),
		1427 => to_unsigned(4469, LUT_AMPL_WIDTH - 1),
		1428 => to_unsigned(4472, LUT_AMPL_WIDTH - 1),
		1429 => to_unsigned(4475, LUT_AMPL_WIDTH - 1),
		1430 => to_unsigned(4478, LUT_AMPL_WIDTH - 1),
		1431 => to_unsigned(4481, LUT_AMPL_WIDTH - 1),
		1432 => to_unsigned(4485, LUT_AMPL_WIDTH - 1),
		1433 => to_unsigned(4488, LUT_AMPL_WIDTH - 1),
		1434 => to_unsigned(4491, LUT_AMPL_WIDTH - 1),
		1435 => to_unsigned(4494, LUT_AMPL_WIDTH - 1),
		1436 => to_unsigned(4497, LUT_AMPL_WIDTH - 1),
		1437 => to_unsigned(4500, LUT_AMPL_WIDTH - 1),
		1438 => to_unsigned(4503, LUT_AMPL_WIDTH - 1),
		1439 => to_unsigned(4506, LUT_AMPL_WIDTH - 1),
		1440 => to_unsigned(4509, LUT_AMPL_WIDTH - 1),
		1441 => to_unsigned(4513, LUT_AMPL_WIDTH - 1),
		1442 => to_unsigned(4516, LUT_AMPL_WIDTH - 1),
		1443 => to_unsigned(4519, LUT_AMPL_WIDTH - 1),
		1444 => to_unsigned(4522, LUT_AMPL_WIDTH - 1),
		1445 => to_unsigned(4525, LUT_AMPL_WIDTH - 1),
		1446 => to_unsigned(4528, LUT_AMPL_WIDTH - 1),
		1447 => to_unsigned(4531, LUT_AMPL_WIDTH - 1),
		1448 => to_unsigned(4534, LUT_AMPL_WIDTH - 1),
		1449 => to_unsigned(4537, LUT_AMPL_WIDTH - 1),
		1450 => to_unsigned(4541, LUT_AMPL_WIDTH - 1),
		1451 => to_unsigned(4544, LUT_AMPL_WIDTH - 1),
		1452 => to_unsigned(4547, LUT_AMPL_WIDTH - 1),
		1453 => to_unsigned(4550, LUT_AMPL_WIDTH - 1),
		1454 => to_unsigned(4553, LUT_AMPL_WIDTH - 1),
		1455 => to_unsigned(4556, LUT_AMPL_WIDTH - 1),
		1456 => to_unsigned(4559, LUT_AMPL_WIDTH - 1),
		1457 => to_unsigned(4562, LUT_AMPL_WIDTH - 1),
		1458 => to_unsigned(4565, LUT_AMPL_WIDTH - 1),
		1459 => to_unsigned(4569, LUT_AMPL_WIDTH - 1),
		1460 => to_unsigned(4572, LUT_AMPL_WIDTH - 1),
		1461 => to_unsigned(4575, LUT_AMPL_WIDTH - 1),
		1462 => to_unsigned(4578, LUT_AMPL_WIDTH - 1),
		1463 => to_unsigned(4581, LUT_AMPL_WIDTH - 1),
		1464 => to_unsigned(4584, LUT_AMPL_WIDTH - 1),
		1465 => to_unsigned(4587, LUT_AMPL_WIDTH - 1),
		1466 => to_unsigned(4590, LUT_AMPL_WIDTH - 1),
		1467 => to_unsigned(4593, LUT_AMPL_WIDTH - 1),
		1468 => to_unsigned(4597, LUT_AMPL_WIDTH - 1),
		1469 => to_unsigned(4600, LUT_AMPL_WIDTH - 1),
		1470 => to_unsigned(4603, LUT_AMPL_WIDTH - 1),
		1471 => to_unsigned(4606, LUT_AMPL_WIDTH - 1),
		1472 => to_unsigned(4609, LUT_AMPL_WIDTH - 1),
		1473 => to_unsigned(4612, LUT_AMPL_WIDTH - 1),
		1474 => to_unsigned(4615, LUT_AMPL_WIDTH - 1),
		1475 => to_unsigned(4618, LUT_AMPL_WIDTH - 1),
		1476 => to_unsigned(4621, LUT_AMPL_WIDTH - 1),
		1477 => to_unsigned(4624, LUT_AMPL_WIDTH - 1),
		1478 => to_unsigned(4628, LUT_AMPL_WIDTH - 1),
		1479 => to_unsigned(4631, LUT_AMPL_WIDTH - 1),
		1480 => to_unsigned(4634, LUT_AMPL_WIDTH - 1),
		1481 => to_unsigned(4637, LUT_AMPL_WIDTH - 1),
		1482 => to_unsigned(4640, LUT_AMPL_WIDTH - 1),
		1483 => to_unsigned(4643, LUT_AMPL_WIDTH - 1),
		1484 => to_unsigned(4646, LUT_AMPL_WIDTH - 1),
		1485 => to_unsigned(4649, LUT_AMPL_WIDTH - 1),
		1486 => to_unsigned(4652, LUT_AMPL_WIDTH - 1),
		1487 => to_unsigned(4656, LUT_AMPL_WIDTH - 1),
		1488 => to_unsigned(4659, LUT_AMPL_WIDTH - 1),
		1489 => to_unsigned(4662, LUT_AMPL_WIDTH - 1),
		1490 => to_unsigned(4665, LUT_AMPL_WIDTH - 1),
		1491 => to_unsigned(4668, LUT_AMPL_WIDTH - 1),
		1492 => to_unsigned(4671, LUT_AMPL_WIDTH - 1),
		1493 => to_unsigned(4674, LUT_AMPL_WIDTH - 1),
		1494 => to_unsigned(4677, LUT_AMPL_WIDTH - 1),
		1495 => to_unsigned(4680, LUT_AMPL_WIDTH - 1),
		1496 => to_unsigned(4684, LUT_AMPL_WIDTH - 1),
		1497 => to_unsigned(4687, LUT_AMPL_WIDTH - 1),
		1498 => to_unsigned(4690, LUT_AMPL_WIDTH - 1),
		1499 => to_unsigned(4693, LUT_AMPL_WIDTH - 1),
		1500 => to_unsigned(4696, LUT_AMPL_WIDTH - 1),
		1501 => to_unsigned(4699, LUT_AMPL_WIDTH - 1),
		1502 => to_unsigned(4702, LUT_AMPL_WIDTH - 1),
		1503 => to_unsigned(4705, LUT_AMPL_WIDTH - 1),
		1504 => to_unsigned(4708, LUT_AMPL_WIDTH - 1),
		1505 => to_unsigned(4712, LUT_AMPL_WIDTH - 1),
		1506 => to_unsigned(4715, LUT_AMPL_WIDTH - 1),
		1507 => to_unsigned(4718, LUT_AMPL_WIDTH - 1),
		1508 => to_unsigned(4721, LUT_AMPL_WIDTH - 1),
		1509 => to_unsigned(4724, LUT_AMPL_WIDTH - 1),
		1510 => to_unsigned(4727, LUT_AMPL_WIDTH - 1),
		1511 => to_unsigned(4730, LUT_AMPL_WIDTH - 1),
		1512 => to_unsigned(4733, LUT_AMPL_WIDTH - 1),
		1513 => to_unsigned(4736, LUT_AMPL_WIDTH - 1),
		1514 => to_unsigned(4740, LUT_AMPL_WIDTH - 1),
		1515 => to_unsigned(4743, LUT_AMPL_WIDTH - 1),
		1516 => to_unsigned(4746, LUT_AMPL_WIDTH - 1),
		1517 => to_unsigned(4749, LUT_AMPL_WIDTH - 1),
		1518 => to_unsigned(4752, LUT_AMPL_WIDTH - 1),
		1519 => to_unsigned(4755, LUT_AMPL_WIDTH - 1),
		1520 => to_unsigned(4758, LUT_AMPL_WIDTH - 1),
		1521 => to_unsigned(4761, LUT_AMPL_WIDTH - 1),
		1522 => to_unsigned(4764, LUT_AMPL_WIDTH - 1),
		1523 => to_unsigned(4768, LUT_AMPL_WIDTH - 1),
		1524 => to_unsigned(4771, LUT_AMPL_WIDTH - 1),
		1525 => to_unsigned(4774, LUT_AMPL_WIDTH - 1),
		1526 => to_unsigned(4777, LUT_AMPL_WIDTH - 1),
		1527 => to_unsigned(4780, LUT_AMPL_WIDTH - 1),
		1528 => to_unsigned(4783, LUT_AMPL_WIDTH - 1),
		1529 => to_unsigned(4786, LUT_AMPL_WIDTH - 1),
		1530 => to_unsigned(4789, LUT_AMPL_WIDTH - 1),
		1531 => to_unsigned(4792, LUT_AMPL_WIDTH - 1),
		1532 => to_unsigned(4795, LUT_AMPL_WIDTH - 1),
		1533 => to_unsigned(4799, LUT_AMPL_WIDTH - 1),
		1534 => to_unsigned(4802, LUT_AMPL_WIDTH - 1),
		1535 => to_unsigned(4805, LUT_AMPL_WIDTH - 1),
		1536 => to_unsigned(4808, LUT_AMPL_WIDTH - 1),
		1537 => to_unsigned(4811, LUT_AMPL_WIDTH - 1),
		1538 => to_unsigned(4814, LUT_AMPL_WIDTH - 1),
		1539 => to_unsigned(4817, LUT_AMPL_WIDTH - 1),
		1540 => to_unsigned(4820, LUT_AMPL_WIDTH - 1),
		1541 => to_unsigned(4823, LUT_AMPL_WIDTH - 1),
		1542 => to_unsigned(4827, LUT_AMPL_WIDTH - 1),
		1543 => to_unsigned(4830, LUT_AMPL_WIDTH - 1),
		1544 => to_unsigned(4833, LUT_AMPL_WIDTH - 1),
		1545 => to_unsigned(4836, LUT_AMPL_WIDTH - 1),
		1546 => to_unsigned(4839, LUT_AMPL_WIDTH - 1),
		1547 => to_unsigned(4842, LUT_AMPL_WIDTH - 1),
		1548 => to_unsigned(4845, LUT_AMPL_WIDTH - 1),
		1549 => to_unsigned(4848, LUT_AMPL_WIDTH - 1),
		1550 => to_unsigned(4851, LUT_AMPL_WIDTH - 1),
		1551 => to_unsigned(4855, LUT_AMPL_WIDTH - 1),
		1552 => to_unsigned(4858, LUT_AMPL_WIDTH - 1),
		1553 => to_unsigned(4861, LUT_AMPL_WIDTH - 1),
		1554 => to_unsigned(4864, LUT_AMPL_WIDTH - 1),
		1555 => to_unsigned(4867, LUT_AMPL_WIDTH - 1),
		1556 => to_unsigned(4870, LUT_AMPL_WIDTH - 1),
		1557 => to_unsigned(4873, LUT_AMPL_WIDTH - 1),
		1558 => to_unsigned(4876, LUT_AMPL_WIDTH - 1),
		1559 => to_unsigned(4879, LUT_AMPL_WIDTH - 1),
		1560 => to_unsigned(4882, LUT_AMPL_WIDTH - 1),
		1561 => to_unsigned(4886, LUT_AMPL_WIDTH - 1),
		1562 => to_unsigned(4889, LUT_AMPL_WIDTH - 1),
		1563 => to_unsigned(4892, LUT_AMPL_WIDTH - 1),
		1564 => to_unsigned(4895, LUT_AMPL_WIDTH - 1),
		1565 => to_unsigned(4898, LUT_AMPL_WIDTH - 1),
		1566 => to_unsigned(4901, LUT_AMPL_WIDTH - 1),
		1567 => to_unsigned(4904, LUT_AMPL_WIDTH - 1),
		1568 => to_unsigned(4907, LUT_AMPL_WIDTH - 1),
		1569 => to_unsigned(4910, LUT_AMPL_WIDTH - 1),
		1570 => to_unsigned(4914, LUT_AMPL_WIDTH - 1),
		1571 => to_unsigned(4917, LUT_AMPL_WIDTH - 1),
		1572 => to_unsigned(4920, LUT_AMPL_WIDTH - 1),
		1573 => to_unsigned(4923, LUT_AMPL_WIDTH - 1),
		1574 => to_unsigned(4926, LUT_AMPL_WIDTH - 1),
		1575 => to_unsigned(4929, LUT_AMPL_WIDTH - 1),
		1576 => to_unsigned(4932, LUT_AMPL_WIDTH - 1),
		1577 => to_unsigned(4935, LUT_AMPL_WIDTH - 1),
		1578 => to_unsigned(4938, LUT_AMPL_WIDTH - 1),
		1579 => to_unsigned(4941, LUT_AMPL_WIDTH - 1),
		1580 => to_unsigned(4945, LUT_AMPL_WIDTH - 1),
		1581 => to_unsigned(4948, LUT_AMPL_WIDTH - 1),
		1582 => to_unsigned(4951, LUT_AMPL_WIDTH - 1),
		1583 => to_unsigned(4954, LUT_AMPL_WIDTH - 1),
		1584 => to_unsigned(4957, LUT_AMPL_WIDTH - 1),
		1585 => to_unsigned(4960, LUT_AMPL_WIDTH - 1),
		1586 => to_unsigned(4963, LUT_AMPL_WIDTH - 1),
		1587 => to_unsigned(4966, LUT_AMPL_WIDTH - 1),
		1588 => to_unsigned(4969, LUT_AMPL_WIDTH - 1),
		1589 => to_unsigned(4973, LUT_AMPL_WIDTH - 1),
		1590 => to_unsigned(4976, LUT_AMPL_WIDTH - 1),
		1591 => to_unsigned(4979, LUT_AMPL_WIDTH - 1),
		1592 => to_unsigned(4982, LUT_AMPL_WIDTH - 1),
		1593 => to_unsigned(4985, LUT_AMPL_WIDTH - 1),
		1594 => to_unsigned(4988, LUT_AMPL_WIDTH - 1),
		1595 => to_unsigned(4991, LUT_AMPL_WIDTH - 1),
		1596 => to_unsigned(4994, LUT_AMPL_WIDTH - 1),
		1597 => to_unsigned(4997, LUT_AMPL_WIDTH - 1),
		1598 => to_unsigned(5000, LUT_AMPL_WIDTH - 1),
		1599 => to_unsigned(5004, LUT_AMPL_WIDTH - 1),
		1600 => to_unsigned(5007, LUT_AMPL_WIDTH - 1),
		1601 => to_unsigned(5010, LUT_AMPL_WIDTH - 1),
		1602 => to_unsigned(5013, LUT_AMPL_WIDTH - 1),
		1603 => to_unsigned(5016, LUT_AMPL_WIDTH - 1),
		1604 => to_unsigned(5019, LUT_AMPL_WIDTH - 1),
		1605 => to_unsigned(5022, LUT_AMPL_WIDTH - 1),
		1606 => to_unsigned(5025, LUT_AMPL_WIDTH - 1),
		1607 => to_unsigned(5028, LUT_AMPL_WIDTH - 1),
		1608 => to_unsigned(5032, LUT_AMPL_WIDTH - 1),
		1609 => to_unsigned(5035, LUT_AMPL_WIDTH - 1),
		1610 => to_unsigned(5038, LUT_AMPL_WIDTH - 1),
		1611 => to_unsigned(5041, LUT_AMPL_WIDTH - 1),
		1612 => to_unsigned(5044, LUT_AMPL_WIDTH - 1),
		1613 => to_unsigned(5047, LUT_AMPL_WIDTH - 1),
		1614 => to_unsigned(5050, LUT_AMPL_WIDTH - 1),
		1615 => to_unsigned(5053, LUT_AMPL_WIDTH - 1),
		1616 => to_unsigned(5056, LUT_AMPL_WIDTH - 1),
		1617 => to_unsigned(5059, LUT_AMPL_WIDTH - 1),
		1618 => to_unsigned(5063, LUT_AMPL_WIDTH - 1),
		1619 => to_unsigned(5066, LUT_AMPL_WIDTH - 1),
		1620 => to_unsigned(5069, LUT_AMPL_WIDTH - 1),
		1621 => to_unsigned(5072, LUT_AMPL_WIDTH - 1),
		1622 => to_unsigned(5075, LUT_AMPL_WIDTH - 1),
		1623 => to_unsigned(5078, LUT_AMPL_WIDTH - 1),
		1624 => to_unsigned(5081, LUT_AMPL_WIDTH - 1),
		1625 => to_unsigned(5084, LUT_AMPL_WIDTH - 1),
		1626 => to_unsigned(5087, LUT_AMPL_WIDTH - 1),
		1627 => to_unsigned(5091, LUT_AMPL_WIDTH - 1),
		1628 => to_unsigned(5094, LUT_AMPL_WIDTH - 1),
		1629 => to_unsigned(5097, LUT_AMPL_WIDTH - 1),
		1630 => to_unsigned(5100, LUT_AMPL_WIDTH - 1),
		1631 => to_unsigned(5103, LUT_AMPL_WIDTH - 1),
		1632 => to_unsigned(5106, LUT_AMPL_WIDTH - 1),
		1633 => to_unsigned(5109, LUT_AMPL_WIDTH - 1),
		1634 => to_unsigned(5112, LUT_AMPL_WIDTH - 1),
		1635 => to_unsigned(5115, LUT_AMPL_WIDTH - 1),
		1636 => to_unsigned(5118, LUT_AMPL_WIDTH - 1),
		1637 => to_unsigned(5122, LUT_AMPL_WIDTH - 1),
		1638 => to_unsigned(5125, LUT_AMPL_WIDTH - 1),
		1639 => to_unsigned(5128, LUT_AMPL_WIDTH - 1),
		1640 => to_unsigned(5131, LUT_AMPL_WIDTH - 1),
		1641 => to_unsigned(5134, LUT_AMPL_WIDTH - 1),
		1642 => to_unsigned(5137, LUT_AMPL_WIDTH - 1),
		1643 => to_unsigned(5140, LUT_AMPL_WIDTH - 1),
		1644 => to_unsigned(5143, LUT_AMPL_WIDTH - 1),
		1645 => to_unsigned(5146, LUT_AMPL_WIDTH - 1),
		1646 => to_unsigned(5149, LUT_AMPL_WIDTH - 1),
		1647 => to_unsigned(5153, LUT_AMPL_WIDTH - 1),
		1648 => to_unsigned(5156, LUT_AMPL_WIDTH - 1),
		1649 => to_unsigned(5159, LUT_AMPL_WIDTH - 1),
		1650 => to_unsigned(5162, LUT_AMPL_WIDTH - 1),
		1651 => to_unsigned(5165, LUT_AMPL_WIDTH - 1),
		1652 => to_unsigned(5168, LUT_AMPL_WIDTH - 1),
		1653 => to_unsigned(5171, LUT_AMPL_WIDTH - 1),
		1654 => to_unsigned(5174, LUT_AMPL_WIDTH - 1),
		1655 => to_unsigned(5177, LUT_AMPL_WIDTH - 1),
		1656 => to_unsigned(5180, LUT_AMPL_WIDTH - 1),
		1657 => to_unsigned(5184, LUT_AMPL_WIDTH - 1),
		1658 => to_unsigned(5187, LUT_AMPL_WIDTH - 1),
		1659 => to_unsigned(5190, LUT_AMPL_WIDTH - 1),
		1660 => to_unsigned(5193, LUT_AMPL_WIDTH - 1),
		1661 => to_unsigned(5196, LUT_AMPL_WIDTH - 1),
		1662 => to_unsigned(5199, LUT_AMPL_WIDTH - 1),
		1663 => to_unsigned(5202, LUT_AMPL_WIDTH - 1),
		1664 => to_unsigned(5205, LUT_AMPL_WIDTH - 1),
		1665 => to_unsigned(5208, LUT_AMPL_WIDTH - 1),
		1666 => to_unsigned(5212, LUT_AMPL_WIDTH - 1),
		1667 => to_unsigned(5215, LUT_AMPL_WIDTH - 1),
		1668 => to_unsigned(5218, LUT_AMPL_WIDTH - 1),
		1669 => to_unsigned(5221, LUT_AMPL_WIDTH - 1),
		1670 => to_unsigned(5224, LUT_AMPL_WIDTH - 1),
		1671 => to_unsigned(5227, LUT_AMPL_WIDTH - 1),
		1672 => to_unsigned(5230, LUT_AMPL_WIDTH - 1),
		1673 => to_unsigned(5233, LUT_AMPL_WIDTH - 1),
		1674 => to_unsigned(5236, LUT_AMPL_WIDTH - 1),
		1675 => to_unsigned(5239, LUT_AMPL_WIDTH - 1),
		1676 => to_unsigned(5243, LUT_AMPL_WIDTH - 1),
		1677 => to_unsigned(5246, LUT_AMPL_WIDTH - 1),
		1678 => to_unsigned(5249, LUT_AMPL_WIDTH - 1),
		1679 => to_unsigned(5252, LUT_AMPL_WIDTH - 1),
		1680 => to_unsigned(5255, LUT_AMPL_WIDTH - 1),
		1681 => to_unsigned(5258, LUT_AMPL_WIDTH - 1),
		1682 => to_unsigned(5261, LUT_AMPL_WIDTH - 1),
		1683 => to_unsigned(5264, LUT_AMPL_WIDTH - 1),
		1684 => to_unsigned(5267, LUT_AMPL_WIDTH - 1),
		1685 => to_unsigned(5270, LUT_AMPL_WIDTH - 1),
		1686 => to_unsigned(5274, LUT_AMPL_WIDTH - 1),
		1687 => to_unsigned(5277, LUT_AMPL_WIDTH - 1),
		1688 => to_unsigned(5280, LUT_AMPL_WIDTH - 1),
		1689 => to_unsigned(5283, LUT_AMPL_WIDTH - 1),
		1690 => to_unsigned(5286, LUT_AMPL_WIDTH - 1),
		1691 => to_unsigned(5289, LUT_AMPL_WIDTH - 1),
		1692 => to_unsigned(5292, LUT_AMPL_WIDTH - 1),
		1693 => to_unsigned(5295, LUT_AMPL_WIDTH - 1),
		1694 => to_unsigned(5298, LUT_AMPL_WIDTH - 1),
		1695 => to_unsigned(5301, LUT_AMPL_WIDTH - 1),
		1696 => to_unsigned(5305, LUT_AMPL_WIDTH - 1),
		1697 => to_unsigned(5308, LUT_AMPL_WIDTH - 1),
		1698 => to_unsigned(5311, LUT_AMPL_WIDTH - 1),
		1699 => to_unsigned(5314, LUT_AMPL_WIDTH - 1),
		1700 => to_unsigned(5317, LUT_AMPL_WIDTH - 1),
		1701 => to_unsigned(5320, LUT_AMPL_WIDTH - 1),
		1702 => to_unsigned(5323, LUT_AMPL_WIDTH - 1),
		1703 => to_unsigned(5326, LUT_AMPL_WIDTH - 1),
		1704 => to_unsigned(5329, LUT_AMPL_WIDTH - 1),
		1705 => to_unsigned(5332, LUT_AMPL_WIDTH - 1),
		1706 => to_unsigned(5336, LUT_AMPL_WIDTH - 1),
		1707 => to_unsigned(5339, LUT_AMPL_WIDTH - 1),
		1708 => to_unsigned(5342, LUT_AMPL_WIDTH - 1),
		1709 => to_unsigned(5345, LUT_AMPL_WIDTH - 1),
		1710 => to_unsigned(5348, LUT_AMPL_WIDTH - 1),
		1711 => to_unsigned(5351, LUT_AMPL_WIDTH - 1),
		1712 => to_unsigned(5354, LUT_AMPL_WIDTH - 1),
		1713 => to_unsigned(5357, LUT_AMPL_WIDTH - 1),
		1714 => to_unsigned(5360, LUT_AMPL_WIDTH - 1),
		1715 => to_unsigned(5363, LUT_AMPL_WIDTH - 1),
		1716 => to_unsigned(5367, LUT_AMPL_WIDTH - 1),
		1717 => to_unsigned(5370, LUT_AMPL_WIDTH - 1),
		1718 => to_unsigned(5373, LUT_AMPL_WIDTH - 1),
		1719 => to_unsigned(5376, LUT_AMPL_WIDTH - 1),
		1720 => to_unsigned(5379, LUT_AMPL_WIDTH - 1),
		1721 => to_unsigned(5382, LUT_AMPL_WIDTH - 1),
		1722 => to_unsigned(5385, LUT_AMPL_WIDTH - 1),
		1723 => to_unsigned(5388, LUT_AMPL_WIDTH - 1),
		1724 => to_unsigned(5391, LUT_AMPL_WIDTH - 1),
		1725 => to_unsigned(5394, LUT_AMPL_WIDTH - 1),
		1726 => to_unsigned(5398, LUT_AMPL_WIDTH - 1),
		1727 => to_unsigned(5401, LUT_AMPL_WIDTH - 1),
		1728 => to_unsigned(5404, LUT_AMPL_WIDTH - 1),
		1729 => to_unsigned(5407, LUT_AMPL_WIDTH - 1),
		1730 => to_unsigned(5410, LUT_AMPL_WIDTH - 1),
		1731 => to_unsigned(5413, LUT_AMPL_WIDTH - 1),
		1732 => to_unsigned(5416, LUT_AMPL_WIDTH - 1),
		1733 => to_unsigned(5419, LUT_AMPL_WIDTH - 1),
		1734 => to_unsigned(5422, LUT_AMPL_WIDTH - 1),
		1735 => to_unsigned(5425, LUT_AMPL_WIDTH - 1),
		1736 => to_unsigned(5428, LUT_AMPL_WIDTH - 1),
		1737 => to_unsigned(5432, LUT_AMPL_WIDTH - 1),
		1738 => to_unsigned(5435, LUT_AMPL_WIDTH - 1),
		1739 => to_unsigned(5438, LUT_AMPL_WIDTH - 1),
		1740 => to_unsigned(5441, LUT_AMPL_WIDTH - 1),
		1741 => to_unsigned(5444, LUT_AMPL_WIDTH - 1),
		1742 => to_unsigned(5447, LUT_AMPL_WIDTH - 1),
		1743 => to_unsigned(5450, LUT_AMPL_WIDTH - 1),
		1744 => to_unsigned(5453, LUT_AMPL_WIDTH - 1),
		1745 => to_unsigned(5456, LUT_AMPL_WIDTH - 1),
		1746 => to_unsigned(5459, LUT_AMPL_WIDTH - 1),
		1747 => to_unsigned(5463, LUT_AMPL_WIDTH - 1),
		1748 => to_unsigned(5466, LUT_AMPL_WIDTH - 1),
		1749 => to_unsigned(5469, LUT_AMPL_WIDTH - 1),
		1750 => to_unsigned(5472, LUT_AMPL_WIDTH - 1),
		1751 => to_unsigned(5475, LUT_AMPL_WIDTH - 1),
		1752 => to_unsigned(5478, LUT_AMPL_WIDTH - 1),
		1753 => to_unsigned(5481, LUT_AMPL_WIDTH - 1),
		1754 => to_unsigned(5484, LUT_AMPL_WIDTH - 1),
		1755 => to_unsigned(5487, LUT_AMPL_WIDTH - 1),
		1756 => to_unsigned(5490, LUT_AMPL_WIDTH - 1),
		1757 => to_unsigned(5494, LUT_AMPL_WIDTH - 1),
		1758 => to_unsigned(5497, LUT_AMPL_WIDTH - 1),
		1759 => to_unsigned(5500, LUT_AMPL_WIDTH - 1),
		1760 => to_unsigned(5503, LUT_AMPL_WIDTH - 1),
		1761 => to_unsigned(5506, LUT_AMPL_WIDTH - 1),
		1762 => to_unsigned(5509, LUT_AMPL_WIDTH - 1),
		1763 => to_unsigned(5512, LUT_AMPL_WIDTH - 1),
		1764 => to_unsigned(5515, LUT_AMPL_WIDTH - 1),
		1765 => to_unsigned(5518, LUT_AMPL_WIDTH - 1),
		1766 => to_unsigned(5521, LUT_AMPL_WIDTH - 1),
		1767 => to_unsigned(5525, LUT_AMPL_WIDTH - 1),
		1768 => to_unsigned(5528, LUT_AMPL_WIDTH - 1),
		1769 => to_unsigned(5531, LUT_AMPL_WIDTH - 1),
		1770 => to_unsigned(5534, LUT_AMPL_WIDTH - 1),
		1771 => to_unsigned(5537, LUT_AMPL_WIDTH - 1),
		1772 => to_unsigned(5540, LUT_AMPL_WIDTH - 1),
		1773 => to_unsigned(5543, LUT_AMPL_WIDTH - 1),
		1774 => to_unsigned(5546, LUT_AMPL_WIDTH - 1),
		1775 => to_unsigned(5549, LUT_AMPL_WIDTH - 1),
		1776 => to_unsigned(5552, LUT_AMPL_WIDTH - 1),
		1777 => to_unsigned(5555, LUT_AMPL_WIDTH - 1),
		1778 => to_unsigned(5559, LUT_AMPL_WIDTH - 1),
		1779 => to_unsigned(5562, LUT_AMPL_WIDTH - 1),
		1780 => to_unsigned(5565, LUT_AMPL_WIDTH - 1),
		1781 => to_unsigned(5568, LUT_AMPL_WIDTH - 1),
		1782 => to_unsigned(5571, LUT_AMPL_WIDTH - 1),
		1783 => to_unsigned(5574, LUT_AMPL_WIDTH - 1),
		1784 => to_unsigned(5577, LUT_AMPL_WIDTH - 1),
		1785 => to_unsigned(5580, LUT_AMPL_WIDTH - 1),
		1786 => to_unsigned(5583, LUT_AMPL_WIDTH - 1),
		1787 => to_unsigned(5586, LUT_AMPL_WIDTH - 1),
		1788 => to_unsigned(5590, LUT_AMPL_WIDTH - 1),
		1789 => to_unsigned(5593, LUT_AMPL_WIDTH - 1),
		1790 => to_unsigned(5596, LUT_AMPL_WIDTH - 1),
		1791 => to_unsigned(5599, LUT_AMPL_WIDTH - 1),
		1792 => to_unsigned(5602, LUT_AMPL_WIDTH - 1),
		1793 => to_unsigned(5605, LUT_AMPL_WIDTH - 1),
		1794 => to_unsigned(5608, LUT_AMPL_WIDTH - 1),
		1795 => to_unsigned(5611, LUT_AMPL_WIDTH - 1),
		1796 => to_unsigned(5614, LUT_AMPL_WIDTH - 1),
		1797 => to_unsigned(5617, LUT_AMPL_WIDTH - 1),
		1798 => to_unsigned(5620, LUT_AMPL_WIDTH - 1),
		1799 => to_unsigned(5624, LUT_AMPL_WIDTH - 1),
		1800 => to_unsigned(5627, LUT_AMPL_WIDTH - 1),
		1801 => to_unsigned(5630, LUT_AMPL_WIDTH - 1),
		1802 => to_unsigned(5633, LUT_AMPL_WIDTH - 1),
		1803 => to_unsigned(5636, LUT_AMPL_WIDTH - 1),
		1804 => to_unsigned(5639, LUT_AMPL_WIDTH - 1),
		1805 => to_unsigned(5642, LUT_AMPL_WIDTH - 1),
		1806 => to_unsigned(5645, LUT_AMPL_WIDTH - 1),
		1807 => to_unsigned(5648, LUT_AMPL_WIDTH - 1),
		1808 => to_unsigned(5651, LUT_AMPL_WIDTH - 1),
		1809 => to_unsigned(5655, LUT_AMPL_WIDTH - 1),
		1810 => to_unsigned(5658, LUT_AMPL_WIDTH - 1),
		1811 => to_unsigned(5661, LUT_AMPL_WIDTH - 1),
		1812 => to_unsigned(5664, LUT_AMPL_WIDTH - 1),
		1813 => to_unsigned(5667, LUT_AMPL_WIDTH - 1),
		1814 => to_unsigned(5670, LUT_AMPL_WIDTH - 1),
		1815 => to_unsigned(5673, LUT_AMPL_WIDTH - 1),
		1816 => to_unsigned(5676, LUT_AMPL_WIDTH - 1),
		1817 => to_unsigned(5679, LUT_AMPL_WIDTH - 1),
		1818 => to_unsigned(5682, LUT_AMPL_WIDTH - 1),
		1819 => to_unsigned(5685, LUT_AMPL_WIDTH - 1),
		1820 => to_unsigned(5689, LUT_AMPL_WIDTH - 1),
		1821 => to_unsigned(5692, LUT_AMPL_WIDTH - 1),
		1822 => to_unsigned(5695, LUT_AMPL_WIDTH - 1),
		1823 => to_unsigned(5698, LUT_AMPL_WIDTH - 1),
		1824 => to_unsigned(5701, LUT_AMPL_WIDTH - 1),
		1825 => to_unsigned(5704, LUT_AMPL_WIDTH - 1),
		1826 => to_unsigned(5707, LUT_AMPL_WIDTH - 1),
		1827 => to_unsigned(5710, LUT_AMPL_WIDTH - 1),
		1828 => to_unsigned(5713, LUT_AMPL_WIDTH - 1),
		1829 => to_unsigned(5716, LUT_AMPL_WIDTH - 1),
		1830 => to_unsigned(5719, LUT_AMPL_WIDTH - 1),
		1831 => to_unsigned(5723, LUT_AMPL_WIDTH - 1),
		1832 => to_unsigned(5726, LUT_AMPL_WIDTH - 1),
		1833 => to_unsigned(5729, LUT_AMPL_WIDTH - 1),
		1834 => to_unsigned(5732, LUT_AMPL_WIDTH - 1),
		1835 => to_unsigned(5735, LUT_AMPL_WIDTH - 1),
		1836 => to_unsigned(5738, LUT_AMPL_WIDTH - 1),
		1837 => to_unsigned(5741, LUT_AMPL_WIDTH - 1),
		1838 => to_unsigned(5744, LUT_AMPL_WIDTH - 1),
		1839 => to_unsigned(5747, LUT_AMPL_WIDTH - 1),
		1840 => to_unsigned(5750, LUT_AMPL_WIDTH - 1),
		1841 => to_unsigned(5754, LUT_AMPL_WIDTH - 1),
		1842 => to_unsigned(5757, LUT_AMPL_WIDTH - 1),
		1843 => to_unsigned(5760, LUT_AMPL_WIDTH - 1),
		1844 => to_unsigned(5763, LUT_AMPL_WIDTH - 1),
		1845 => to_unsigned(5766, LUT_AMPL_WIDTH - 1),
		1846 => to_unsigned(5769, LUT_AMPL_WIDTH - 1),
		1847 => to_unsigned(5772, LUT_AMPL_WIDTH - 1),
		1848 => to_unsigned(5775, LUT_AMPL_WIDTH - 1),
		1849 => to_unsigned(5778, LUT_AMPL_WIDTH - 1),
		1850 => to_unsigned(5781, LUT_AMPL_WIDTH - 1),
		1851 => to_unsigned(5784, LUT_AMPL_WIDTH - 1),
		1852 => to_unsigned(5788, LUT_AMPL_WIDTH - 1),
		1853 => to_unsigned(5791, LUT_AMPL_WIDTH - 1),
		1854 => to_unsigned(5794, LUT_AMPL_WIDTH - 1),
		1855 => to_unsigned(5797, LUT_AMPL_WIDTH - 1),
		1856 => to_unsigned(5800, LUT_AMPL_WIDTH - 1),
		1857 => to_unsigned(5803, LUT_AMPL_WIDTH - 1),
		1858 => to_unsigned(5806, LUT_AMPL_WIDTH - 1),
		1859 => to_unsigned(5809, LUT_AMPL_WIDTH - 1),
		1860 => to_unsigned(5812, LUT_AMPL_WIDTH - 1),
		1861 => to_unsigned(5815, LUT_AMPL_WIDTH - 1),
		1862 => to_unsigned(5818, LUT_AMPL_WIDTH - 1),
		1863 => to_unsigned(5822, LUT_AMPL_WIDTH - 1),
		1864 => to_unsigned(5825, LUT_AMPL_WIDTH - 1),
		1865 => to_unsigned(5828, LUT_AMPL_WIDTH - 1),
		1866 => to_unsigned(5831, LUT_AMPL_WIDTH - 1),
		1867 => to_unsigned(5834, LUT_AMPL_WIDTH - 1),
		1868 => to_unsigned(5837, LUT_AMPL_WIDTH - 1),
		1869 => to_unsigned(5840, LUT_AMPL_WIDTH - 1),
		1870 => to_unsigned(5843, LUT_AMPL_WIDTH - 1),
		1871 => to_unsigned(5846, LUT_AMPL_WIDTH - 1),
		1872 => to_unsigned(5849, LUT_AMPL_WIDTH - 1),
		1873 => to_unsigned(5852, LUT_AMPL_WIDTH - 1),
		1874 => to_unsigned(5856, LUT_AMPL_WIDTH - 1),
		1875 => to_unsigned(5859, LUT_AMPL_WIDTH - 1),
		1876 => to_unsigned(5862, LUT_AMPL_WIDTH - 1),
		1877 => to_unsigned(5865, LUT_AMPL_WIDTH - 1),
		1878 => to_unsigned(5868, LUT_AMPL_WIDTH - 1),
		1879 => to_unsigned(5871, LUT_AMPL_WIDTH - 1),
		1880 => to_unsigned(5874, LUT_AMPL_WIDTH - 1),
		1881 => to_unsigned(5877, LUT_AMPL_WIDTH - 1),
		1882 => to_unsigned(5880, LUT_AMPL_WIDTH - 1),
		1883 => to_unsigned(5883, LUT_AMPL_WIDTH - 1),
		1884 => to_unsigned(5886, LUT_AMPL_WIDTH - 1),
		1885 => to_unsigned(5890, LUT_AMPL_WIDTH - 1),
		1886 => to_unsigned(5893, LUT_AMPL_WIDTH - 1),
		1887 => to_unsigned(5896, LUT_AMPL_WIDTH - 1),
		1888 => to_unsigned(5899, LUT_AMPL_WIDTH - 1),
		1889 => to_unsigned(5902, LUT_AMPL_WIDTH - 1),
		1890 => to_unsigned(5905, LUT_AMPL_WIDTH - 1),
		1891 => to_unsigned(5908, LUT_AMPL_WIDTH - 1),
		1892 => to_unsigned(5911, LUT_AMPL_WIDTH - 1),
		1893 => to_unsigned(5914, LUT_AMPL_WIDTH - 1),
		1894 => to_unsigned(5917, LUT_AMPL_WIDTH - 1),
		1895 => to_unsigned(5920, LUT_AMPL_WIDTH - 1),
		1896 => to_unsigned(5924, LUT_AMPL_WIDTH - 1),
		1897 => to_unsigned(5927, LUT_AMPL_WIDTH - 1),
		1898 => to_unsigned(5930, LUT_AMPL_WIDTH - 1),
		1899 => to_unsigned(5933, LUT_AMPL_WIDTH - 1),
		1900 => to_unsigned(5936, LUT_AMPL_WIDTH - 1),
		1901 => to_unsigned(5939, LUT_AMPL_WIDTH - 1),
		1902 => to_unsigned(5942, LUT_AMPL_WIDTH - 1),
		1903 => to_unsigned(5945, LUT_AMPL_WIDTH - 1),
		1904 => to_unsigned(5948, LUT_AMPL_WIDTH - 1),
		1905 => to_unsigned(5951, LUT_AMPL_WIDTH - 1),
		1906 => to_unsigned(5954, LUT_AMPL_WIDTH - 1),
		1907 => to_unsigned(5958, LUT_AMPL_WIDTH - 1),
		1908 => to_unsigned(5961, LUT_AMPL_WIDTH - 1),
		1909 => to_unsigned(5964, LUT_AMPL_WIDTH - 1),
		1910 => to_unsigned(5967, LUT_AMPL_WIDTH - 1),
		1911 => to_unsigned(5970, LUT_AMPL_WIDTH - 1),
		1912 => to_unsigned(5973, LUT_AMPL_WIDTH - 1),
		1913 => to_unsigned(5976, LUT_AMPL_WIDTH - 1),
		1914 => to_unsigned(5979, LUT_AMPL_WIDTH - 1),
		1915 => to_unsigned(5982, LUT_AMPL_WIDTH - 1),
		1916 => to_unsigned(5985, LUT_AMPL_WIDTH - 1),
		1917 => to_unsigned(5988, LUT_AMPL_WIDTH - 1),
		1918 => to_unsigned(5991, LUT_AMPL_WIDTH - 1),
		1919 => to_unsigned(5995, LUT_AMPL_WIDTH - 1),
		1920 => to_unsigned(5998, LUT_AMPL_WIDTH - 1),
		1921 => to_unsigned(6001, LUT_AMPL_WIDTH - 1),
		1922 => to_unsigned(6004, LUT_AMPL_WIDTH - 1),
		1923 => to_unsigned(6007, LUT_AMPL_WIDTH - 1),
		1924 => to_unsigned(6010, LUT_AMPL_WIDTH - 1),
		1925 => to_unsigned(6013, LUT_AMPL_WIDTH - 1),
		1926 => to_unsigned(6016, LUT_AMPL_WIDTH - 1),
		1927 => to_unsigned(6019, LUT_AMPL_WIDTH - 1),
		1928 => to_unsigned(6022, LUT_AMPL_WIDTH - 1),
		1929 => to_unsigned(6025, LUT_AMPL_WIDTH - 1),
		1930 => to_unsigned(6029, LUT_AMPL_WIDTH - 1),
		1931 => to_unsigned(6032, LUT_AMPL_WIDTH - 1),
		1932 => to_unsigned(6035, LUT_AMPL_WIDTH - 1),
		1933 => to_unsigned(6038, LUT_AMPL_WIDTH - 1),
		1934 => to_unsigned(6041, LUT_AMPL_WIDTH - 1),
		1935 => to_unsigned(6044, LUT_AMPL_WIDTH - 1),
		1936 => to_unsigned(6047, LUT_AMPL_WIDTH - 1),
		1937 => to_unsigned(6050, LUT_AMPL_WIDTH - 1),
		1938 => to_unsigned(6053, LUT_AMPL_WIDTH - 1),
		1939 => to_unsigned(6056, LUT_AMPL_WIDTH - 1),
		1940 => to_unsigned(6059, LUT_AMPL_WIDTH - 1),
		1941 => to_unsigned(6063, LUT_AMPL_WIDTH - 1),
		1942 => to_unsigned(6066, LUT_AMPL_WIDTH - 1),
		1943 => to_unsigned(6069, LUT_AMPL_WIDTH - 1),
		1944 => to_unsigned(6072, LUT_AMPL_WIDTH - 1),
		1945 => to_unsigned(6075, LUT_AMPL_WIDTH - 1),
		1946 => to_unsigned(6078, LUT_AMPL_WIDTH - 1),
		1947 => to_unsigned(6081, LUT_AMPL_WIDTH - 1),
		1948 => to_unsigned(6084, LUT_AMPL_WIDTH - 1),
		1949 => to_unsigned(6087, LUT_AMPL_WIDTH - 1),
		1950 => to_unsigned(6090, LUT_AMPL_WIDTH - 1),
		1951 => to_unsigned(6093, LUT_AMPL_WIDTH - 1),
		1952 => to_unsigned(6096, LUT_AMPL_WIDTH - 1),
		1953 => to_unsigned(6100, LUT_AMPL_WIDTH - 1),
		1954 => to_unsigned(6103, LUT_AMPL_WIDTH - 1),
		1955 => to_unsigned(6106, LUT_AMPL_WIDTH - 1),
		1956 => to_unsigned(6109, LUT_AMPL_WIDTH - 1),
		1957 => to_unsigned(6112, LUT_AMPL_WIDTH - 1),
		1958 => to_unsigned(6115, LUT_AMPL_WIDTH - 1),
		1959 => to_unsigned(6118, LUT_AMPL_WIDTH - 1),
		1960 => to_unsigned(6121, LUT_AMPL_WIDTH - 1),
		1961 => to_unsigned(6124, LUT_AMPL_WIDTH - 1),
		1962 => to_unsigned(6127, LUT_AMPL_WIDTH - 1),
		1963 => to_unsigned(6130, LUT_AMPL_WIDTH - 1),
		1964 => to_unsigned(6134, LUT_AMPL_WIDTH - 1),
		1965 => to_unsigned(6137, LUT_AMPL_WIDTH - 1),
		1966 => to_unsigned(6140, LUT_AMPL_WIDTH - 1),
		1967 => to_unsigned(6143, LUT_AMPL_WIDTH - 1),
		1968 => to_unsigned(6146, LUT_AMPL_WIDTH - 1),
		1969 => to_unsigned(6149, LUT_AMPL_WIDTH - 1),
		1970 => to_unsigned(6152, LUT_AMPL_WIDTH - 1),
		1971 => to_unsigned(6155, LUT_AMPL_WIDTH - 1),
		1972 => to_unsigned(6158, LUT_AMPL_WIDTH - 1),
		1973 => to_unsigned(6161, LUT_AMPL_WIDTH - 1),
		1974 => to_unsigned(6164, LUT_AMPL_WIDTH - 1),
		1975 => to_unsigned(6167, LUT_AMPL_WIDTH - 1),
		1976 => to_unsigned(6171, LUT_AMPL_WIDTH - 1),
		1977 => to_unsigned(6174, LUT_AMPL_WIDTH - 1),
		1978 => to_unsigned(6177, LUT_AMPL_WIDTH - 1),
		1979 => to_unsigned(6180, LUT_AMPL_WIDTH - 1),
		1980 => to_unsigned(6183, LUT_AMPL_WIDTH - 1),
		1981 => to_unsigned(6186, LUT_AMPL_WIDTH - 1),
		1982 => to_unsigned(6189, LUT_AMPL_WIDTH - 1),
		1983 => to_unsigned(6192, LUT_AMPL_WIDTH - 1),
		1984 => to_unsigned(6195, LUT_AMPL_WIDTH - 1),
		1985 => to_unsigned(6198, LUT_AMPL_WIDTH - 1),
		1986 => to_unsigned(6201, LUT_AMPL_WIDTH - 1),
		1987 => to_unsigned(6204, LUT_AMPL_WIDTH - 1),
		1988 => to_unsigned(6208, LUT_AMPL_WIDTH - 1),
		1989 => to_unsigned(6211, LUT_AMPL_WIDTH - 1),
		1990 => to_unsigned(6214, LUT_AMPL_WIDTH - 1),
		1991 => to_unsigned(6217, LUT_AMPL_WIDTH - 1),
		1992 => to_unsigned(6220, LUT_AMPL_WIDTH - 1),
		1993 => to_unsigned(6223, LUT_AMPL_WIDTH - 1),
		1994 => to_unsigned(6226, LUT_AMPL_WIDTH - 1),
		1995 => to_unsigned(6229, LUT_AMPL_WIDTH - 1),
		1996 => to_unsigned(6232, LUT_AMPL_WIDTH - 1),
		1997 => to_unsigned(6235, LUT_AMPL_WIDTH - 1),
		1998 => to_unsigned(6238, LUT_AMPL_WIDTH - 1),
		1999 => to_unsigned(6241, LUT_AMPL_WIDTH - 1),
		2000 => to_unsigned(6245, LUT_AMPL_WIDTH - 1),
		2001 => to_unsigned(6248, LUT_AMPL_WIDTH - 1),
		2002 => to_unsigned(6251, LUT_AMPL_WIDTH - 1),
		2003 => to_unsigned(6254, LUT_AMPL_WIDTH - 1),
		2004 => to_unsigned(6257, LUT_AMPL_WIDTH - 1),
		2005 => to_unsigned(6260, LUT_AMPL_WIDTH - 1),
		2006 => to_unsigned(6263, LUT_AMPL_WIDTH - 1),
		2007 => to_unsigned(6266, LUT_AMPL_WIDTH - 1),
		2008 => to_unsigned(6269, LUT_AMPL_WIDTH - 1),
		2009 => to_unsigned(6272, LUT_AMPL_WIDTH - 1),
		2010 => to_unsigned(6275, LUT_AMPL_WIDTH - 1),
		2011 => to_unsigned(6278, LUT_AMPL_WIDTH - 1),
		2012 => to_unsigned(6282, LUT_AMPL_WIDTH - 1),
		2013 => to_unsigned(6285, LUT_AMPL_WIDTH - 1),
		2014 => to_unsigned(6288, LUT_AMPL_WIDTH - 1),
		2015 => to_unsigned(6291, LUT_AMPL_WIDTH - 1),
		2016 => to_unsigned(6294, LUT_AMPL_WIDTH - 1),
		2017 => to_unsigned(6297, LUT_AMPL_WIDTH - 1),
		2018 => to_unsigned(6300, LUT_AMPL_WIDTH - 1),
		2019 => to_unsigned(6303, LUT_AMPL_WIDTH - 1),
		2020 => to_unsigned(6306, LUT_AMPL_WIDTH - 1),
		2021 => to_unsigned(6309, LUT_AMPL_WIDTH - 1),
		2022 => to_unsigned(6312, LUT_AMPL_WIDTH - 1),
		2023 => to_unsigned(6315, LUT_AMPL_WIDTH - 1),
		2024 => to_unsigned(6319, LUT_AMPL_WIDTH - 1),
		2025 => to_unsigned(6322, LUT_AMPL_WIDTH - 1),
		2026 => to_unsigned(6325, LUT_AMPL_WIDTH - 1),
		2027 => to_unsigned(6328, LUT_AMPL_WIDTH - 1),
		2028 => to_unsigned(6331, LUT_AMPL_WIDTH - 1),
		2029 => to_unsigned(6334, LUT_AMPL_WIDTH - 1),
		2030 => to_unsigned(6337, LUT_AMPL_WIDTH - 1),
		2031 => to_unsigned(6340, LUT_AMPL_WIDTH - 1),
		2032 => to_unsigned(6343, LUT_AMPL_WIDTH - 1),
		2033 => to_unsigned(6346, LUT_AMPL_WIDTH - 1),
		2034 => to_unsigned(6349, LUT_AMPL_WIDTH - 1),
		2035 => to_unsigned(6352, LUT_AMPL_WIDTH - 1),
		2036 => to_unsigned(6356, LUT_AMPL_WIDTH - 1),
		2037 => to_unsigned(6359, LUT_AMPL_WIDTH - 1),
		2038 => to_unsigned(6362, LUT_AMPL_WIDTH - 1),
		2039 => to_unsigned(6365, LUT_AMPL_WIDTH - 1),
		2040 => to_unsigned(6368, LUT_AMPL_WIDTH - 1),
		2041 => to_unsigned(6371, LUT_AMPL_WIDTH - 1),
		2042 => to_unsigned(6374, LUT_AMPL_WIDTH - 1),
		2043 => to_unsigned(6377, LUT_AMPL_WIDTH - 1),
		2044 => to_unsigned(6380, LUT_AMPL_WIDTH - 1),
		2045 => to_unsigned(6383, LUT_AMPL_WIDTH - 1),
		2046 => to_unsigned(6386, LUT_AMPL_WIDTH - 1),
		2047 => to_unsigned(6389, LUT_AMPL_WIDTH - 1),
		2048 => to_unsigned(6393, LUT_AMPL_WIDTH - 1),
		2049 => to_unsigned(6396, LUT_AMPL_WIDTH - 1),
		2050 => to_unsigned(6399, LUT_AMPL_WIDTH - 1),
		2051 => to_unsigned(6402, LUT_AMPL_WIDTH - 1),
		2052 => to_unsigned(6405, LUT_AMPL_WIDTH - 1),
		2053 => to_unsigned(6408, LUT_AMPL_WIDTH - 1),
		2054 => to_unsigned(6411, LUT_AMPL_WIDTH - 1),
		2055 => to_unsigned(6414, LUT_AMPL_WIDTH - 1),
		2056 => to_unsigned(6417, LUT_AMPL_WIDTH - 1),
		2057 => to_unsigned(6420, LUT_AMPL_WIDTH - 1),
		2058 => to_unsigned(6423, LUT_AMPL_WIDTH - 1),
		2059 => to_unsigned(6426, LUT_AMPL_WIDTH - 1),
		2060 => to_unsigned(6429, LUT_AMPL_WIDTH - 1),
		2061 => to_unsigned(6433, LUT_AMPL_WIDTH - 1),
		2062 => to_unsigned(6436, LUT_AMPL_WIDTH - 1),
		2063 => to_unsigned(6439, LUT_AMPL_WIDTH - 1),
		2064 => to_unsigned(6442, LUT_AMPL_WIDTH - 1),
		2065 => to_unsigned(6445, LUT_AMPL_WIDTH - 1),
		2066 => to_unsigned(6448, LUT_AMPL_WIDTH - 1),
		2067 => to_unsigned(6451, LUT_AMPL_WIDTH - 1),
		2068 => to_unsigned(6454, LUT_AMPL_WIDTH - 1),
		2069 => to_unsigned(6457, LUT_AMPL_WIDTH - 1),
		2070 => to_unsigned(6460, LUT_AMPL_WIDTH - 1),
		2071 => to_unsigned(6463, LUT_AMPL_WIDTH - 1),
		2072 => to_unsigned(6466, LUT_AMPL_WIDTH - 1),
		2073 => to_unsigned(6470, LUT_AMPL_WIDTH - 1),
		2074 => to_unsigned(6473, LUT_AMPL_WIDTH - 1),
		2075 => to_unsigned(6476, LUT_AMPL_WIDTH - 1),
		2076 => to_unsigned(6479, LUT_AMPL_WIDTH - 1),
		2077 => to_unsigned(6482, LUT_AMPL_WIDTH - 1),
		2078 => to_unsigned(6485, LUT_AMPL_WIDTH - 1),
		2079 => to_unsigned(6488, LUT_AMPL_WIDTH - 1),
		2080 => to_unsigned(6491, LUT_AMPL_WIDTH - 1),
		2081 => to_unsigned(6494, LUT_AMPL_WIDTH - 1),
		2082 => to_unsigned(6497, LUT_AMPL_WIDTH - 1),
		2083 => to_unsigned(6500, LUT_AMPL_WIDTH - 1),
		2084 => to_unsigned(6503, LUT_AMPL_WIDTH - 1),
		2085 => to_unsigned(6506, LUT_AMPL_WIDTH - 1),
		2086 => to_unsigned(6510, LUT_AMPL_WIDTH - 1),
		2087 => to_unsigned(6513, LUT_AMPL_WIDTH - 1),
		2088 => to_unsigned(6516, LUT_AMPL_WIDTH - 1),
		2089 => to_unsigned(6519, LUT_AMPL_WIDTH - 1),
		2090 => to_unsigned(6522, LUT_AMPL_WIDTH - 1),
		2091 => to_unsigned(6525, LUT_AMPL_WIDTH - 1),
		2092 => to_unsigned(6528, LUT_AMPL_WIDTH - 1),
		2093 => to_unsigned(6531, LUT_AMPL_WIDTH - 1),
		2094 => to_unsigned(6534, LUT_AMPL_WIDTH - 1),
		2095 => to_unsigned(6537, LUT_AMPL_WIDTH - 1),
		2096 => to_unsigned(6540, LUT_AMPL_WIDTH - 1),
		2097 => to_unsigned(6543, LUT_AMPL_WIDTH - 1),
		2098 => to_unsigned(6547, LUT_AMPL_WIDTH - 1),
		2099 => to_unsigned(6550, LUT_AMPL_WIDTH - 1),
		2100 => to_unsigned(6553, LUT_AMPL_WIDTH - 1),
		2101 => to_unsigned(6556, LUT_AMPL_WIDTH - 1),
		2102 => to_unsigned(6559, LUT_AMPL_WIDTH - 1),
		2103 => to_unsigned(6562, LUT_AMPL_WIDTH - 1),
		2104 => to_unsigned(6565, LUT_AMPL_WIDTH - 1),
		2105 => to_unsigned(6568, LUT_AMPL_WIDTH - 1),
		2106 => to_unsigned(6571, LUT_AMPL_WIDTH - 1),
		2107 => to_unsigned(6574, LUT_AMPL_WIDTH - 1),
		2108 => to_unsigned(6577, LUT_AMPL_WIDTH - 1),
		2109 => to_unsigned(6580, LUT_AMPL_WIDTH - 1),
		2110 => to_unsigned(6583, LUT_AMPL_WIDTH - 1),
		2111 => to_unsigned(6587, LUT_AMPL_WIDTH - 1),
		2112 => to_unsigned(6590, LUT_AMPL_WIDTH - 1),
		2113 => to_unsigned(6593, LUT_AMPL_WIDTH - 1),
		2114 => to_unsigned(6596, LUT_AMPL_WIDTH - 1),
		2115 => to_unsigned(6599, LUT_AMPL_WIDTH - 1),
		2116 => to_unsigned(6602, LUT_AMPL_WIDTH - 1),
		2117 => to_unsigned(6605, LUT_AMPL_WIDTH - 1),
		2118 => to_unsigned(6608, LUT_AMPL_WIDTH - 1),
		2119 => to_unsigned(6611, LUT_AMPL_WIDTH - 1),
		2120 => to_unsigned(6614, LUT_AMPL_WIDTH - 1),
		2121 => to_unsigned(6617, LUT_AMPL_WIDTH - 1),
		2122 => to_unsigned(6620, LUT_AMPL_WIDTH - 1),
		2123 => to_unsigned(6623, LUT_AMPL_WIDTH - 1),
		2124 => to_unsigned(6627, LUT_AMPL_WIDTH - 1),
		2125 => to_unsigned(6630, LUT_AMPL_WIDTH - 1),
		2126 => to_unsigned(6633, LUT_AMPL_WIDTH - 1),
		2127 => to_unsigned(6636, LUT_AMPL_WIDTH - 1),
		2128 => to_unsigned(6639, LUT_AMPL_WIDTH - 1),
		2129 => to_unsigned(6642, LUT_AMPL_WIDTH - 1),
		2130 => to_unsigned(6645, LUT_AMPL_WIDTH - 1),
		2131 => to_unsigned(6648, LUT_AMPL_WIDTH - 1),
		2132 => to_unsigned(6651, LUT_AMPL_WIDTH - 1),
		2133 => to_unsigned(6654, LUT_AMPL_WIDTH - 1),
		2134 => to_unsigned(6657, LUT_AMPL_WIDTH - 1),
		2135 => to_unsigned(6660, LUT_AMPL_WIDTH - 1),
		2136 => to_unsigned(6663, LUT_AMPL_WIDTH - 1),
		2137 => to_unsigned(6667, LUT_AMPL_WIDTH - 1),
		2138 => to_unsigned(6670, LUT_AMPL_WIDTH - 1),
		2139 => to_unsigned(6673, LUT_AMPL_WIDTH - 1),
		2140 => to_unsigned(6676, LUT_AMPL_WIDTH - 1),
		2141 => to_unsigned(6679, LUT_AMPL_WIDTH - 1),
		2142 => to_unsigned(6682, LUT_AMPL_WIDTH - 1),
		2143 => to_unsigned(6685, LUT_AMPL_WIDTH - 1),
		2144 => to_unsigned(6688, LUT_AMPL_WIDTH - 1),
		2145 => to_unsigned(6691, LUT_AMPL_WIDTH - 1),
		2146 => to_unsigned(6694, LUT_AMPL_WIDTH - 1),
		2147 => to_unsigned(6697, LUT_AMPL_WIDTH - 1),
		2148 => to_unsigned(6700, LUT_AMPL_WIDTH - 1),
		2149 => to_unsigned(6703, LUT_AMPL_WIDTH - 1),
		2150 => to_unsigned(6706, LUT_AMPL_WIDTH - 1),
		2151 => to_unsigned(6710, LUT_AMPL_WIDTH - 1),
		2152 => to_unsigned(6713, LUT_AMPL_WIDTH - 1),
		2153 => to_unsigned(6716, LUT_AMPL_WIDTH - 1),
		2154 => to_unsigned(6719, LUT_AMPL_WIDTH - 1),
		2155 => to_unsigned(6722, LUT_AMPL_WIDTH - 1),
		2156 => to_unsigned(6725, LUT_AMPL_WIDTH - 1),
		2157 => to_unsigned(6728, LUT_AMPL_WIDTH - 1),
		2158 => to_unsigned(6731, LUT_AMPL_WIDTH - 1),
		2159 => to_unsigned(6734, LUT_AMPL_WIDTH - 1),
		2160 => to_unsigned(6737, LUT_AMPL_WIDTH - 1),
		2161 => to_unsigned(6740, LUT_AMPL_WIDTH - 1),
		2162 => to_unsigned(6743, LUT_AMPL_WIDTH - 1),
		2163 => to_unsigned(6746, LUT_AMPL_WIDTH - 1),
		2164 => to_unsigned(6750, LUT_AMPL_WIDTH - 1),
		2165 => to_unsigned(6753, LUT_AMPL_WIDTH - 1),
		2166 => to_unsigned(6756, LUT_AMPL_WIDTH - 1),
		2167 => to_unsigned(6759, LUT_AMPL_WIDTH - 1),
		2168 => to_unsigned(6762, LUT_AMPL_WIDTH - 1),
		2169 => to_unsigned(6765, LUT_AMPL_WIDTH - 1),
		2170 => to_unsigned(6768, LUT_AMPL_WIDTH - 1),
		2171 => to_unsigned(6771, LUT_AMPL_WIDTH - 1),
		2172 => to_unsigned(6774, LUT_AMPL_WIDTH - 1),
		2173 => to_unsigned(6777, LUT_AMPL_WIDTH - 1),
		2174 => to_unsigned(6780, LUT_AMPL_WIDTH - 1),
		2175 => to_unsigned(6783, LUT_AMPL_WIDTH - 1),
		2176 => to_unsigned(6786, LUT_AMPL_WIDTH - 1),
		2177 => to_unsigned(6789, LUT_AMPL_WIDTH - 1),
		2178 => to_unsigned(6793, LUT_AMPL_WIDTH - 1),
		2179 => to_unsigned(6796, LUT_AMPL_WIDTH - 1),
		2180 => to_unsigned(6799, LUT_AMPL_WIDTH - 1),
		2181 => to_unsigned(6802, LUT_AMPL_WIDTH - 1),
		2182 => to_unsigned(6805, LUT_AMPL_WIDTH - 1),
		2183 => to_unsigned(6808, LUT_AMPL_WIDTH - 1),
		2184 => to_unsigned(6811, LUT_AMPL_WIDTH - 1),
		2185 => to_unsigned(6814, LUT_AMPL_WIDTH - 1),
		2186 => to_unsigned(6817, LUT_AMPL_WIDTH - 1),
		2187 => to_unsigned(6820, LUT_AMPL_WIDTH - 1),
		2188 => to_unsigned(6823, LUT_AMPL_WIDTH - 1),
		2189 => to_unsigned(6826, LUT_AMPL_WIDTH - 1),
		2190 => to_unsigned(6829, LUT_AMPL_WIDTH - 1),
		2191 => to_unsigned(6833, LUT_AMPL_WIDTH - 1),
		2192 => to_unsigned(6836, LUT_AMPL_WIDTH - 1),
		2193 => to_unsigned(6839, LUT_AMPL_WIDTH - 1),
		2194 => to_unsigned(6842, LUT_AMPL_WIDTH - 1),
		2195 => to_unsigned(6845, LUT_AMPL_WIDTH - 1),
		2196 => to_unsigned(6848, LUT_AMPL_WIDTH - 1),
		2197 => to_unsigned(6851, LUT_AMPL_WIDTH - 1),
		2198 => to_unsigned(6854, LUT_AMPL_WIDTH - 1),
		2199 => to_unsigned(6857, LUT_AMPL_WIDTH - 1),
		2200 => to_unsigned(6860, LUT_AMPL_WIDTH - 1),
		2201 => to_unsigned(6863, LUT_AMPL_WIDTH - 1),
		2202 => to_unsigned(6866, LUT_AMPL_WIDTH - 1),
		2203 => to_unsigned(6869, LUT_AMPL_WIDTH - 1),
		2204 => to_unsigned(6872, LUT_AMPL_WIDTH - 1),
		2205 => to_unsigned(6876, LUT_AMPL_WIDTH - 1),
		2206 => to_unsigned(6879, LUT_AMPL_WIDTH - 1),
		2207 => to_unsigned(6882, LUT_AMPL_WIDTH - 1),
		2208 => to_unsigned(6885, LUT_AMPL_WIDTH - 1),
		2209 => to_unsigned(6888, LUT_AMPL_WIDTH - 1),
		2210 => to_unsigned(6891, LUT_AMPL_WIDTH - 1),
		2211 => to_unsigned(6894, LUT_AMPL_WIDTH - 1),
		2212 => to_unsigned(6897, LUT_AMPL_WIDTH - 1),
		2213 => to_unsigned(6900, LUT_AMPL_WIDTH - 1),
		2214 => to_unsigned(6903, LUT_AMPL_WIDTH - 1),
		2215 => to_unsigned(6906, LUT_AMPL_WIDTH - 1),
		2216 => to_unsigned(6909, LUT_AMPL_WIDTH - 1),
		2217 => to_unsigned(6912, LUT_AMPL_WIDTH - 1),
		2218 => to_unsigned(6915, LUT_AMPL_WIDTH - 1),
		2219 => to_unsigned(6919, LUT_AMPL_WIDTH - 1),
		2220 => to_unsigned(6922, LUT_AMPL_WIDTH - 1),
		2221 => to_unsigned(6925, LUT_AMPL_WIDTH - 1),
		2222 => to_unsigned(6928, LUT_AMPL_WIDTH - 1),
		2223 => to_unsigned(6931, LUT_AMPL_WIDTH - 1),
		2224 => to_unsigned(6934, LUT_AMPL_WIDTH - 1),
		2225 => to_unsigned(6937, LUT_AMPL_WIDTH - 1),
		2226 => to_unsigned(6940, LUT_AMPL_WIDTH - 1),
		2227 => to_unsigned(6943, LUT_AMPL_WIDTH - 1),
		2228 => to_unsigned(6946, LUT_AMPL_WIDTH - 1),
		2229 => to_unsigned(6949, LUT_AMPL_WIDTH - 1),
		2230 => to_unsigned(6952, LUT_AMPL_WIDTH - 1),
		2231 => to_unsigned(6955, LUT_AMPL_WIDTH - 1),
		2232 => to_unsigned(6958, LUT_AMPL_WIDTH - 1),
		2233 => to_unsigned(6961, LUT_AMPL_WIDTH - 1),
		2234 => to_unsigned(6965, LUT_AMPL_WIDTH - 1),
		2235 => to_unsigned(6968, LUT_AMPL_WIDTH - 1),
		2236 => to_unsigned(6971, LUT_AMPL_WIDTH - 1),
		2237 => to_unsigned(6974, LUT_AMPL_WIDTH - 1),
		2238 => to_unsigned(6977, LUT_AMPL_WIDTH - 1),
		2239 => to_unsigned(6980, LUT_AMPL_WIDTH - 1),
		2240 => to_unsigned(6983, LUT_AMPL_WIDTH - 1),
		2241 => to_unsigned(6986, LUT_AMPL_WIDTH - 1),
		2242 => to_unsigned(6989, LUT_AMPL_WIDTH - 1),
		2243 => to_unsigned(6992, LUT_AMPL_WIDTH - 1),
		2244 => to_unsigned(6995, LUT_AMPL_WIDTH - 1),
		2245 => to_unsigned(6998, LUT_AMPL_WIDTH - 1),
		2246 => to_unsigned(7001, LUT_AMPL_WIDTH - 1),
		2247 => to_unsigned(7004, LUT_AMPL_WIDTH - 1),
		2248 => to_unsigned(7008, LUT_AMPL_WIDTH - 1),
		2249 => to_unsigned(7011, LUT_AMPL_WIDTH - 1),
		2250 => to_unsigned(7014, LUT_AMPL_WIDTH - 1),
		2251 => to_unsigned(7017, LUT_AMPL_WIDTH - 1),
		2252 => to_unsigned(7020, LUT_AMPL_WIDTH - 1),
		2253 => to_unsigned(7023, LUT_AMPL_WIDTH - 1),
		2254 => to_unsigned(7026, LUT_AMPL_WIDTH - 1),
		2255 => to_unsigned(7029, LUT_AMPL_WIDTH - 1),
		2256 => to_unsigned(7032, LUT_AMPL_WIDTH - 1),
		2257 => to_unsigned(7035, LUT_AMPL_WIDTH - 1),
		2258 => to_unsigned(7038, LUT_AMPL_WIDTH - 1),
		2259 => to_unsigned(7041, LUT_AMPL_WIDTH - 1),
		2260 => to_unsigned(7044, LUT_AMPL_WIDTH - 1),
		2261 => to_unsigned(7047, LUT_AMPL_WIDTH - 1),
		2262 => to_unsigned(7050, LUT_AMPL_WIDTH - 1),
		2263 => to_unsigned(7054, LUT_AMPL_WIDTH - 1),
		2264 => to_unsigned(7057, LUT_AMPL_WIDTH - 1),
		2265 => to_unsigned(7060, LUT_AMPL_WIDTH - 1),
		2266 => to_unsigned(7063, LUT_AMPL_WIDTH - 1),
		2267 => to_unsigned(7066, LUT_AMPL_WIDTH - 1),
		2268 => to_unsigned(7069, LUT_AMPL_WIDTH - 1),
		2269 => to_unsigned(7072, LUT_AMPL_WIDTH - 1),
		2270 => to_unsigned(7075, LUT_AMPL_WIDTH - 1),
		2271 => to_unsigned(7078, LUT_AMPL_WIDTH - 1),
		2272 => to_unsigned(7081, LUT_AMPL_WIDTH - 1),
		2273 => to_unsigned(7084, LUT_AMPL_WIDTH - 1),
		2274 => to_unsigned(7087, LUT_AMPL_WIDTH - 1),
		2275 => to_unsigned(7090, LUT_AMPL_WIDTH - 1),
		2276 => to_unsigned(7093, LUT_AMPL_WIDTH - 1),
		2277 => to_unsigned(7097, LUT_AMPL_WIDTH - 1),
		2278 => to_unsigned(7100, LUT_AMPL_WIDTH - 1),
		2279 => to_unsigned(7103, LUT_AMPL_WIDTH - 1),
		2280 => to_unsigned(7106, LUT_AMPL_WIDTH - 1),
		2281 => to_unsigned(7109, LUT_AMPL_WIDTH - 1),
		2282 => to_unsigned(7112, LUT_AMPL_WIDTH - 1),
		2283 => to_unsigned(7115, LUT_AMPL_WIDTH - 1),
		2284 => to_unsigned(7118, LUT_AMPL_WIDTH - 1),
		2285 => to_unsigned(7121, LUT_AMPL_WIDTH - 1),
		2286 => to_unsigned(7124, LUT_AMPL_WIDTH - 1),
		2287 => to_unsigned(7127, LUT_AMPL_WIDTH - 1),
		2288 => to_unsigned(7130, LUT_AMPL_WIDTH - 1),
		2289 => to_unsigned(7133, LUT_AMPL_WIDTH - 1),
		2290 => to_unsigned(7136, LUT_AMPL_WIDTH - 1),
		2291 => to_unsigned(7139, LUT_AMPL_WIDTH - 1),
		2292 => to_unsigned(7143, LUT_AMPL_WIDTH - 1),
		2293 => to_unsigned(7146, LUT_AMPL_WIDTH - 1),
		2294 => to_unsigned(7149, LUT_AMPL_WIDTH - 1),
		2295 => to_unsigned(7152, LUT_AMPL_WIDTH - 1),
		2296 => to_unsigned(7155, LUT_AMPL_WIDTH - 1),
		2297 => to_unsigned(7158, LUT_AMPL_WIDTH - 1),
		2298 => to_unsigned(7161, LUT_AMPL_WIDTH - 1),
		2299 => to_unsigned(7164, LUT_AMPL_WIDTH - 1),
		2300 => to_unsigned(7167, LUT_AMPL_WIDTH - 1),
		2301 => to_unsigned(7170, LUT_AMPL_WIDTH - 1),
		2302 => to_unsigned(7173, LUT_AMPL_WIDTH - 1),
		2303 => to_unsigned(7176, LUT_AMPL_WIDTH - 1),
		2304 => to_unsigned(7179, LUT_AMPL_WIDTH - 1),
		2305 => to_unsigned(7182, LUT_AMPL_WIDTH - 1),
		2306 => to_unsigned(7185, LUT_AMPL_WIDTH - 1),
		2307 => to_unsigned(7188, LUT_AMPL_WIDTH - 1),
		2308 => to_unsigned(7192, LUT_AMPL_WIDTH - 1),
		2309 => to_unsigned(7195, LUT_AMPL_WIDTH - 1),
		2310 => to_unsigned(7198, LUT_AMPL_WIDTH - 1),
		2311 => to_unsigned(7201, LUT_AMPL_WIDTH - 1),
		2312 => to_unsigned(7204, LUT_AMPL_WIDTH - 1),
		2313 => to_unsigned(7207, LUT_AMPL_WIDTH - 1),
		2314 => to_unsigned(7210, LUT_AMPL_WIDTH - 1),
		2315 => to_unsigned(7213, LUT_AMPL_WIDTH - 1),
		2316 => to_unsigned(7216, LUT_AMPL_WIDTH - 1),
		2317 => to_unsigned(7219, LUT_AMPL_WIDTH - 1),
		2318 => to_unsigned(7222, LUT_AMPL_WIDTH - 1),
		2319 => to_unsigned(7225, LUT_AMPL_WIDTH - 1),
		2320 => to_unsigned(7228, LUT_AMPL_WIDTH - 1),
		2321 => to_unsigned(7231, LUT_AMPL_WIDTH - 1),
		2322 => to_unsigned(7234, LUT_AMPL_WIDTH - 1),
		2323 => to_unsigned(7238, LUT_AMPL_WIDTH - 1),
		2324 => to_unsigned(7241, LUT_AMPL_WIDTH - 1),
		2325 => to_unsigned(7244, LUT_AMPL_WIDTH - 1),
		2326 => to_unsigned(7247, LUT_AMPL_WIDTH - 1),
		2327 => to_unsigned(7250, LUT_AMPL_WIDTH - 1),
		2328 => to_unsigned(7253, LUT_AMPL_WIDTH - 1),
		2329 => to_unsigned(7256, LUT_AMPL_WIDTH - 1),
		2330 => to_unsigned(7259, LUT_AMPL_WIDTH - 1),
		2331 => to_unsigned(7262, LUT_AMPL_WIDTH - 1),
		2332 => to_unsigned(7265, LUT_AMPL_WIDTH - 1),
		2333 => to_unsigned(7268, LUT_AMPL_WIDTH - 1),
		2334 => to_unsigned(7271, LUT_AMPL_WIDTH - 1),
		2335 => to_unsigned(7274, LUT_AMPL_WIDTH - 1),
		2336 => to_unsigned(7277, LUT_AMPL_WIDTH - 1),
		2337 => to_unsigned(7280, LUT_AMPL_WIDTH - 1),
		2338 => to_unsigned(7283, LUT_AMPL_WIDTH - 1),
		2339 => to_unsigned(7287, LUT_AMPL_WIDTH - 1),
		2340 => to_unsigned(7290, LUT_AMPL_WIDTH - 1),
		2341 => to_unsigned(7293, LUT_AMPL_WIDTH - 1),
		2342 => to_unsigned(7296, LUT_AMPL_WIDTH - 1),
		2343 => to_unsigned(7299, LUT_AMPL_WIDTH - 1),
		2344 => to_unsigned(7302, LUT_AMPL_WIDTH - 1),
		2345 => to_unsigned(7305, LUT_AMPL_WIDTH - 1),
		2346 => to_unsigned(7308, LUT_AMPL_WIDTH - 1),
		2347 => to_unsigned(7311, LUT_AMPL_WIDTH - 1),
		2348 => to_unsigned(7314, LUT_AMPL_WIDTH - 1),
		2349 => to_unsigned(7317, LUT_AMPL_WIDTH - 1),
		2350 => to_unsigned(7320, LUT_AMPL_WIDTH - 1),
		2351 => to_unsigned(7323, LUT_AMPL_WIDTH - 1),
		2352 => to_unsigned(7326, LUT_AMPL_WIDTH - 1),
		2353 => to_unsigned(7329, LUT_AMPL_WIDTH - 1),
		2354 => to_unsigned(7332, LUT_AMPL_WIDTH - 1),
		2355 => to_unsigned(7336, LUT_AMPL_WIDTH - 1),
		2356 => to_unsigned(7339, LUT_AMPL_WIDTH - 1),
		2357 => to_unsigned(7342, LUT_AMPL_WIDTH - 1),
		2358 => to_unsigned(7345, LUT_AMPL_WIDTH - 1),
		2359 => to_unsigned(7348, LUT_AMPL_WIDTH - 1),
		2360 => to_unsigned(7351, LUT_AMPL_WIDTH - 1),
		2361 => to_unsigned(7354, LUT_AMPL_WIDTH - 1),
		2362 => to_unsigned(7357, LUT_AMPL_WIDTH - 1),
		2363 => to_unsigned(7360, LUT_AMPL_WIDTH - 1),
		2364 => to_unsigned(7363, LUT_AMPL_WIDTH - 1),
		2365 => to_unsigned(7366, LUT_AMPL_WIDTH - 1),
		2366 => to_unsigned(7369, LUT_AMPL_WIDTH - 1),
		2367 => to_unsigned(7372, LUT_AMPL_WIDTH - 1),
		2368 => to_unsigned(7375, LUT_AMPL_WIDTH - 1),
		2369 => to_unsigned(7378, LUT_AMPL_WIDTH - 1),
		2370 => to_unsigned(7381, LUT_AMPL_WIDTH - 1),
		2371 => to_unsigned(7385, LUT_AMPL_WIDTH - 1),
		2372 => to_unsigned(7388, LUT_AMPL_WIDTH - 1),
		2373 => to_unsigned(7391, LUT_AMPL_WIDTH - 1),
		2374 => to_unsigned(7394, LUT_AMPL_WIDTH - 1),
		2375 => to_unsigned(7397, LUT_AMPL_WIDTH - 1),
		2376 => to_unsigned(7400, LUT_AMPL_WIDTH - 1),
		2377 => to_unsigned(7403, LUT_AMPL_WIDTH - 1),
		2378 => to_unsigned(7406, LUT_AMPL_WIDTH - 1),
		2379 => to_unsigned(7409, LUT_AMPL_WIDTH - 1),
		2380 => to_unsigned(7412, LUT_AMPL_WIDTH - 1),
		2381 => to_unsigned(7415, LUT_AMPL_WIDTH - 1),
		2382 => to_unsigned(7418, LUT_AMPL_WIDTH - 1),
		2383 => to_unsigned(7421, LUT_AMPL_WIDTH - 1),
		2384 => to_unsigned(7424, LUT_AMPL_WIDTH - 1),
		2385 => to_unsigned(7427, LUT_AMPL_WIDTH - 1),
		2386 => to_unsigned(7430, LUT_AMPL_WIDTH - 1),
		2387 => to_unsigned(7433, LUT_AMPL_WIDTH - 1),
		2388 => to_unsigned(7437, LUT_AMPL_WIDTH - 1),
		2389 => to_unsigned(7440, LUT_AMPL_WIDTH - 1),
		2390 => to_unsigned(7443, LUT_AMPL_WIDTH - 1),
		2391 => to_unsigned(7446, LUT_AMPL_WIDTH - 1),
		2392 => to_unsigned(7449, LUT_AMPL_WIDTH - 1),
		2393 => to_unsigned(7452, LUT_AMPL_WIDTH - 1),
		2394 => to_unsigned(7455, LUT_AMPL_WIDTH - 1),
		2395 => to_unsigned(7458, LUT_AMPL_WIDTH - 1),
		2396 => to_unsigned(7461, LUT_AMPL_WIDTH - 1),
		2397 => to_unsigned(7464, LUT_AMPL_WIDTH - 1),
		2398 => to_unsigned(7467, LUT_AMPL_WIDTH - 1),
		2399 => to_unsigned(7470, LUT_AMPL_WIDTH - 1),
		2400 => to_unsigned(7473, LUT_AMPL_WIDTH - 1),
		2401 => to_unsigned(7476, LUT_AMPL_WIDTH - 1),
		2402 => to_unsigned(7479, LUT_AMPL_WIDTH - 1),
		2403 => to_unsigned(7482, LUT_AMPL_WIDTH - 1),
		2404 => to_unsigned(7485, LUT_AMPL_WIDTH - 1),
		2405 => to_unsigned(7489, LUT_AMPL_WIDTH - 1),
		2406 => to_unsigned(7492, LUT_AMPL_WIDTH - 1),
		2407 => to_unsigned(7495, LUT_AMPL_WIDTH - 1),
		2408 => to_unsigned(7498, LUT_AMPL_WIDTH - 1),
		2409 => to_unsigned(7501, LUT_AMPL_WIDTH - 1),
		2410 => to_unsigned(7504, LUT_AMPL_WIDTH - 1),
		2411 => to_unsigned(7507, LUT_AMPL_WIDTH - 1),
		2412 => to_unsigned(7510, LUT_AMPL_WIDTH - 1),
		2413 => to_unsigned(7513, LUT_AMPL_WIDTH - 1),
		2414 => to_unsigned(7516, LUT_AMPL_WIDTH - 1),
		2415 => to_unsigned(7519, LUT_AMPL_WIDTH - 1),
		2416 => to_unsigned(7522, LUT_AMPL_WIDTH - 1),
		2417 => to_unsigned(7525, LUT_AMPL_WIDTH - 1),
		2418 => to_unsigned(7528, LUT_AMPL_WIDTH - 1),
		2419 => to_unsigned(7531, LUT_AMPL_WIDTH - 1),
		2420 => to_unsigned(7534, LUT_AMPL_WIDTH - 1),
		2421 => to_unsigned(7537, LUT_AMPL_WIDTH - 1),
		2422 => to_unsigned(7541, LUT_AMPL_WIDTH - 1),
		2423 => to_unsigned(7544, LUT_AMPL_WIDTH - 1),
		2424 => to_unsigned(7547, LUT_AMPL_WIDTH - 1),
		2425 => to_unsigned(7550, LUT_AMPL_WIDTH - 1),
		2426 => to_unsigned(7553, LUT_AMPL_WIDTH - 1),
		2427 => to_unsigned(7556, LUT_AMPL_WIDTH - 1),
		2428 => to_unsigned(7559, LUT_AMPL_WIDTH - 1),
		2429 => to_unsigned(7562, LUT_AMPL_WIDTH - 1),
		2430 => to_unsigned(7565, LUT_AMPL_WIDTH - 1),
		2431 => to_unsigned(7568, LUT_AMPL_WIDTH - 1),
		2432 => to_unsigned(7571, LUT_AMPL_WIDTH - 1),
		2433 => to_unsigned(7574, LUT_AMPL_WIDTH - 1),
		2434 => to_unsigned(7577, LUT_AMPL_WIDTH - 1),
		2435 => to_unsigned(7580, LUT_AMPL_WIDTH - 1),
		2436 => to_unsigned(7583, LUT_AMPL_WIDTH - 1),
		2437 => to_unsigned(7586, LUT_AMPL_WIDTH - 1),
		2438 => to_unsigned(7589, LUT_AMPL_WIDTH - 1),
		2439 => to_unsigned(7592, LUT_AMPL_WIDTH - 1),
		2440 => to_unsigned(7596, LUT_AMPL_WIDTH - 1),
		2441 => to_unsigned(7599, LUT_AMPL_WIDTH - 1),
		2442 => to_unsigned(7602, LUT_AMPL_WIDTH - 1),
		2443 => to_unsigned(7605, LUT_AMPL_WIDTH - 1),
		2444 => to_unsigned(7608, LUT_AMPL_WIDTH - 1),
		2445 => to_unsigned(7611, LUT_AMPL_WIDTH - 1),
		2446 => to_unsigned(7614, LUT_AMPL_WIDTH - 1),
		2447 => to_unsigned(7617, LUT_AMPL_WIDTH - 1),
		2448 => to_unsigned(7620, LUT_AMPL_WIDTH - 1),
		2449 => to_unsigned(7623, LUT_AMPL_WIDTH - 1),
		2450 => to_unsigned(7626, LUT_AMPL_WIDTH - 1),
		2451 => to_unsigned(7629, LUT_AMPL_WIDTH - 1),
		2452 => to_unsigned(7632, LUT_AMPL_WIDTH - 1),
		2453 => to_unsigned(7635, LUT_AMPL_WIDTH - 1),
		2454 => to_unsigned(7638, LUT_AMPL_WIDTH - 1),
		2455 => to_unsigned(7641, LUT_AMPL_WIDTH - 1),
		2456 => to_unsigned(7644, LUT_AMPL_WIDTH - 1),
		2457 => to_unsigned(7647, LUT_AMPL_WIDTH - 1),
		2458 => to_unsigned(7651, LUT_AMPL_WIDTH - 1),
		2459 => to_unsigned(7654, LUT_AMPL_WIDTH - 1),
		2460 => to_unsigned(7657, LUT_AMPL_WIDTH - 1),
		2461 => to_unsigned(7660, LUT_AMPL_WIDTH - 1),
		2462 => to_unsigned(7663, LUT_AMPL_WIDTH - 1),
		2463 => to_unsigned(7666, LUT_AMPL_WIDTH - 1),
		2464 => to_unsigned(7669, LUT_AMPL_WIDTH - 1),
		2465 => to_unsigned(7672, LUT_AMPL_WIDTH - 1),
		2466 => to_unsigned(7675, LUT_AMPL_WIDTH - 1),
		2467 => to_unsigned(7678, LUT_AMPL_WIDTH - 1),
		2468 => to_unsigned(7681, LUT_AMPL_WIDTH - 1),
		2469 => to_unsigned(7684, LUT_AMPL_WIDTH - 1),
		2470 => to_unsigned(7687, LUT_AMPL_WIDTH - 1),
		2471 => to_unsigned(7690, LUT_AMPL_WIDTH - 1),
		2472 => to_unsigned(7693, LUT_AMPL_WIDTH - 1),
		2473 => to_unsigned(7696, LUT_AMPL_WIDTH - 1),
		2474 => to_unsigned(7699, LUT_AMPL_WIDTH - 1),
		2475 => to_unsigned(7702, LUT_AMPL_WIDTH - 1),
		2476 => to_unsigned(7705, LUT_AMPL_WIDTH - 1),
		2477 => to_unsigned(7709, LUT_AMPL_WIDTH - 1),
		2478 => to_unsigned(7712, LUT_AMPL_WIDTH - 1),
		2479 => to_unsigned(7715, LUT_AMPL_WIDTH - 1),
		2480 => to_unsigned(7718, LUT_AMPL_WIDTH - 1),
		2481 => to_unsigned(7721, LUT_AMPL_WIDTH - 1),
		2482 => to_unsigned(7724, LUT_AMPL_WIDTH - 1),
		2483 => to_unsigned(7727, LUT_AMPL_WIDTH - 1),
		2484 => to_unsigned(7730, LUT_AMPL_WIDTH - 1),
		2485 => to_unsigned(7733, LUT_AMPL_WIDTH - 1),
		2486 => to_unsigned(7736, LUT_AMPL_WIDTH - 1),
		2487 => to_unsigned(7739, LUT_AMPL_WIDTH - 1),
		2488 => to_unsigned(7742, LUT_AMPL_WIDTH - 1),
		2489 => to_unsigned(7745, LUT_AMPL_WIDTH - 1),
		2490 => to_unsigned(7748, LUT_AMPL_WIDTH - 1),
		2491 => to_unsigned(7751, LUT_AMPL_WIDTH - 1),
		2492 => to_unsigned(7754, LUT_AMPL_WIDTH - 1),
		2493 => to_unsigned(7757, LUT_AMPL_WIDTH - 1),
		2494 => to_unsigned(7760, LUT_AMPL_WIDTH - 1),
		2495 => to_unsigned(7764, LUT_AMPL_WIDTH - 1),
		2496 => to_unsigned(7767, LUT_AMPL_WIDTH - 1),
		2497 => to_unsigned(7770, LUT_AMPL_WIDTH - 1),
		2498 => to_unsigned(7773, LUT_AMPL_WIDTH - 1),
		2499 => to_unsigned(7776, LUT_AMPL_WIDTH - 1),
		2500 => to_unsigned(7779, LUT_AMPL_WIDTH - 1),
		2501 => to_unsigned(7782, LUT_AMPL_WIDTH - 1),
		2502 => to_unsigned(7785, LUT_AMPL_WIDTH - 1),
		2503 => to_unsigned(7788, LUT_AMPL_WIDTH - 1),
		2504 => to_unsigned(7791, LUT_AMPL_WIDTH - 1),
		2505 => to_unsigned(7794, LUT_AMPL_WIDTH - 1),
		2506 => to_unsigned(7797, LUT_AMPL_WIDTH - 1),
		2507 => to_unsigned(7800, LUT_AMPL_WIDTH - 1),
		2508 => to_unsigned(7803, LUT_AMPL_WIDTH - 1),
		2509 => to_unsigned(7806, LUT_AMPL_WIDTH - 1),
		2510 => to_unsigned(7809, LUT_AMPL_WIDTH - 1),
		2511 => to_unsigned(7812, LUT_AMPL_WIDTH - 1),
		2512 => to_unsigned(7815, LUT_AMPL_WIDTH - 1),
		2513 => to_unsigned(7818, LUT_AMPL_WIDTH - 1),
		2514 => to_unsigned(7821, LUT_AMPL_WIDTH - 1),
		2515 => to_unsigned(7825, LUT_AMPL_WIDTH - 1),
		2516 => to_unsigned(7828, LUT_AMPL_WIDTH - 1),
		2517 => to_unsigned(7831, LUT_AMPL_WIDTH - 1),
		2518 => to_unsigned(7834, LUT_AMPL_WIDTH - 1),
		2519 => to_unsigned(7837, LUT_AMPL_WIDTH - 1),
		2520 => to_unsigned(7840, LUT_AMPL_WIDTH - 1),
		2521 => to_unsigned(7843, LUT_AMPL_WIDTH - 1),
		2522 => to_unsigned(7846, LUT_AMPL_WIDTH - 1),
		2523 => to_unsigned(7849, LUT_AMPL_WIDTH - 1),
		2524 => to_unsigned(7852, LUT_AMPL_WIDTH - 1),
		2525 => to_unsigned(7855, LUT_AMPL_WIDTH - 1),
		2526 => to_unsigned(7858, LUT_AMPL_WIDTH - 1),
		2527 => to_unsigned(7861, LUT_AMPL_WIDTH - 1),
		2528 => to_unsigned(7864, LUT_AMPL_WIDTH - 1),
		2529 => to_unsigned(7867, LUT_AMPL_WIDTH - 1),
		2530 => to_unsigned(7870, LUT_AMPL_WIDTH - 1),
		2531 => to_unsigned(7873, LUT_AMPL_WIDTH - 1),
		2532 => to_unsigned(7876, LUT_AMPL_WIDTH - 1),
		2533 => to_unsigned(7879, LUT_AMPL_WIDTH - 1),
		2534 => to_unsigned(7882, LUT_AMPL_WIDTH - 1),
		2535 => to_unsigned(7886, LUT_AMPL_WIDTH - 1),
		2536 => to_unsigned(7889, LUT_AMPL_WIDTH - 1),
		2537 => to_unsigned(7892, LUT_AMPL_WIDTH - 1),
		2538 => to_unsigned(7895, LUT_AMPL_WIDTH - 1),
		2539 => to_unsigned(7898, LUT_AMPL_WIDTH - 1),
		2540 => to_unsigned(7901, LUT_AMPL_WIDTH - 1),
		2541 => to_unsigned(7904, LUT_AMPL_WIDTH - 1),
		2542 => to_unsigned(7907, LUT_AMPL_WIDTH - 1),
		2543 => to_unsigned(7910, LUT_AMPL_WIDTH - 1),
		2544 => to_unsigned(7913, LUT_AMPL_WIDTH - 1),
		2545 => to_unsigned(7916, LUT_AMPL_WIDTH - 1),
		2546 => to_unsigned(7919, LUT_AMPL_WIDTH - 1),
		2547 => to_unsigned(7922, LUT_AMPL_WIDTH - 1),
		2548 => to_unsigned(7925, LUT_AMPL_WIDTH - 1),
		2549 => to_unsigned(7928, LUT_AMPL_WIDTH - 1),
		2550 => to_unsigned(7931, LUT_AMPL_WIDTH - 1),
		2551 => to_unsigned(7934, LUT_AMPL_WIDTH - 1),
		2552 => to_unsigned(7937, LUT_AMPL_WIDTH - 1),
		2553 => to_unsigned(7940, LUT_AMPL_WIDTH - 1),
		2554 => to_unsigned(7943, LUT_AMPL_WIDTH - 1),
		2555 => to_unsigned(7946, LUT_AMPL_WIDTH - 1),
		2556 => to_unsigned(7950, LUT_AMPL_WIDTH - 1),
		2557 => to_unsigned(7953, LUT_AMPL_WIDTH - 1),
		2558 => to_unsigned(7956, LUT_AMPL_WIDTH - 1),
		2559 => to_unsigned(7959, LUT_AMPL_WIDTH - 1),
		2560 => to_unsigned(7962, LUT_AMPL_WIDTH - 1),
		2561 => to_unsigned(7965, LUT_AMPL_WIDTH - 1),
		2562 => to_unsigned(7968, LUT_AMPL_WIDTH - 1),
		2563 => to_unsigned(7971, LUT_AMPL_WIDTH - 1),
		2564 => to_unsigned(7974, LUT_AMPL_WIDTH - 1),
		2565 => to_unsigned(7977, LUT_AMPL_WIDTH - 1),
		2566 => to_unsigned(7980, LUT_AMPL_WIDTH - 1),
		2567 => to_unsigned(7983, LUT_AMPL_WIDTH - 1),
		2568 => to_unsigned(7986, LUT_AMPL_WIDTH - 1),
		2569 => to_unsigned(7989, LUT_AMPL_WIDTH - 1),
		2570 => to_unsigned(7992, LUT_AMPL_WIDTH - 1),
		2571 => to_unsigned(7995, LUT_AMPL_WIDTH - 1),
		2572 => to_unsigned(7998, LUT_AMPL_WIDTH - 1),
		2573 => to_unsigned(8001, LUT_AMPL_WIDTH - 1),
		2574 => to_unsigned(8004, LUT_AMPL_WIDTH - 1),
		2575 => to_unsigned(8007, LUT_AMPL_WIDTH - 1),
		2576 => to_unsigned(8010, LUT_AMPL_WIDTH - 1),
		2577 => to_unsigned(8014, LUT_AMPL_WIDTH - 1),
		2578 => to_unsigned(8017, LUT_AMPL_WIDTH - 1),
		2579 => to_unsigned(8020, LUT_AMPL_WIDTH - 1),
		2580 => to_unsigned(8023, LUT_AMPL_WIDTH - 1),
		2581 => to_unsigned(8026, LUT_AMPL_WIDTH - 1),
		2582 => to_unsigned(8029, LUT_AMPL_WIDTH - 1),
		2583 => to_unsigned(8032, LUT_AMPL_WIDTH - 1),
		2584 => to_unsigned(8035, LUT_AMPL_WIDTH - 1),
		2585 => to_unsigned(8038, LUT_AMPL_WIDTH - 1),
		2586 => to_unsigned(8041, LUT_AMPL_WIDTH - 1),
		2587 => to_unsigned(8044, LUT_AMPL_WIDTH - 1),
		2588 => to_unsigned(8047, LUT_AMPL_WIDTH - 1),
		2589 => to_unsigned(8050, LUT_AMPL_WIDTH - 1),
		2590 => to_unsigned(8053, LUT_AMPL_WIDTH - 1),
		2591 => to_unsigned(8056, LUT_AMPL_WIDTH - 1),
		2592 => to_unsigned(8059, LUT_AMPL_WIDTH - 1),
		2593 => to_unsigned(8062, LUT_AMPL_WIDTH - 1),
		2594 => to_unsigned(8065, LUT_AMPL_WIDTH - 1),
		2595 => to_unsigned(8068, LUT_AMPL_WIDTH - 1),
		2596 => to_unsigned(8071, LUT_AMPL_WIDTH - 1),
		2597 => to_unsigned(8074, LUT_AMPL_WIDTH - 1),
		2598 => to_unsigned(8077, LUT_AMPL_WIDTH - 1),
		2599 => to_unsigned(8081, LUT_AMPL_WIDTH - 1),
		2600 => to_unsigned(8084, LUT_AMPL_WIDTH - 1),
		2601 => to_unsigned(8087, LUT_AMPL_WIDTH - 1),
		2602 => to_unsigned(8090, LUT_AMPL_WIDTH - 1),
		2603 => to_unsigned(8093, LUT_AMPL_WIDTH - 1),
		2604 => to_unsigned(8096, LUT_AMPL_WIDTH - 1),
		2605 => to_unsigned(8099, LUT_AMPL_WIDTH - 1),
		2606 => to_unsigned(8102, LUT_AMPL_WIDTH - 1),
		2607 => to_unsigned(8105, LUT_AMPL_WIDTH - 1),
		2608 => to_unsigned(8108, LUT_AMPL_WIDTH - 1),
		2609 => to_unsigned(8111, LUT_AMPL_WIDTH - 1),
		2610 => to_unsigned(8114, LUT_AMPL_WIDTH - 1),
		2611 => to_unsigned(8117, LUT_AMPL_WIDTH - 1),
		2612 => to_unsigned(8120, LUT_AMPL_WIDTH - 1),
		2613 => to_unsigned(8123, LUT_AMPL_WIDTH - 1),
		2614 => to_unsigned(8126, LUT_AMPL_WIDTH - 1),
		2615 => to_unsigned(8129, LUT_AMPL_WIDTH - 1),
		2616 => to_unsigned(8132, LUT_AMPL_WIDTH - 1),
		2617 => to_unsigned(8135, LUT_AMPL_WIDTH - 1),
		2618 => to_unsigned(8138, LUT_AMPL_WIDTH - 1),
		2619 => to_unsigned(8141, LUT_AMPL_WIDTH - 1),
		2620 => to_unsigned(8144, LUT_AMPL_WIDTH - 1),
		2621 => to_unsigned(8147, LUT_AMPL_WIDTH - 1),
		2622 => to_unsigned(8151, LUT_AMPL_WIDTH - 1),
		2623 => to_unsigned(8154, LUT_AMPL_WIDTH - 1),
		2624 => to_unsigned(8157, LUT_AMPL_WIDTH - 1),
		2625 => to_unsigned(8160, LUT_AMPL_WIDTH - 1),
		2626 => to_unsigned(8163, LUT_AMPL_WIDTH - 1),
		2627 => to_unsigned(8166, LUT_AMPL_WIDTH - 1),
		2628 => to_unsigned(8169, LUT_AMPL_WIDTH - 1),
		2629 => to_unsigned(8172, LUT_AMPL_WIDTH - 1),
		2630 => to_unsigned(8175, LUT_AMPL_WIDTH - 1),
		2631 => to_unsigned(8178, LUT_AMPL_WIDTH - 1),
		2632 => to_unsigned(8181, LUT_AMPL_WIDTH - 1),
		2633 => to_unsigned(8184, LUT_AMPL_WIDTH - 1),
		2634 => to_unsigned(8187, LUT_AMPL_WIDTH - 1),
		2635 => to_unsigned(8190, LUT_AMPL_WIDTH - 1),
		2636 => to_unsigned(8193, LUT_AMPL_WIDTH - 1),
		2637 => to_unsigned(8196, LUT_AMPL_WIDTH - 1),
		2638 => to_unsigned(8199, LUT_AMPL_WIDTH - 1),
		2639 => to_unsigned(8202, LUT_AMPL_WIDTH - 1),
		2640 => to_unsigned(8205, LUT_AMPL_WIDTH - 1),
		2641 => to_unsigned(8208, LUT_AMPL_WIDTH - 1),
		2642 => to_unsigned(8211, LUT_AMPL_WIDTH - 1),
		2643 => to_unsigned(8214, LUT_AMPL_WIDTH - 1),
		2644 => to_unsigned(8217, LUT_AMPL_WIDTH - 1),
		2645 => to_unsigned(8220, LUT_AMPL_WIDTH - 1),
		2646 => to_unsigned(8224, LUT_AMPL_WIDTH - 1),
		2647 => to_unsigned(8227, LUT_AMPL_WIDTH - 1),
		2648 => to_unsigned(8230, LUT_AMPL_WIDTH - 1),
		2649 => to_unsigned(8233, LUT_AMPL_WIDTH - 1),
		2650 => to_unsigned(8236, LUT_AMPL_WIDTH - 1),
		2651 => to_unsigned(8239, LUT_AMPL_WIDTH - 1),
		2652 => to_unsigned(8242, LUT_AMPL_WIDTH - 1),
		2653 => to_unsigned(8245, LUT_AMPL_WIDTH - 1),
		2654 => to_unsigned(8248, LUT_AMPL_WIDTH - 1),
		2655 => to_unsigned(8251, LUT_AMPL_WIDTH - 1),
		2656 => to_unsigned(8254, LUT_AMPL_WIDTH - 1),
		2657 => to_unsigned(8257, LUT_AMPL_WIDTH - 1),
		2658 => to_unsigned(8260, LUT_AMPL_WIDTH - 1),
		2659 => to_unsigned(8263, LUT_AMPL_WIDTH - 1),
		2660 => to_unsigned(8266, LUT_AMPL_WIDTH - 1),
		2661 => to_unsigned(8269, LUT_AMPL_WIDTH - 1),
		2662 => to_unsigned(8272, LUT_AMPL_WIDTH - 1),
		2663 => to_unsigned(8275, LUT_AMPL_WIDTH - 1),
		2664 => to_unsigned(8278, LUT_AMPL_WIDTH - 1),
		2665 => to_unsigned(8281, LUT_AMPL_WIDTH - 1),
		2666 => to_unsigned(8284, LUT_AMPL_WIDTH - 1),
		2667 => to_unsigned(8287, LUT_AMPL_WIDTH - 1),
		2668 => to_unsigned(8290, LUT_AMPL_WIDTH - 1),
		2669 => to_unsigned(8293, LUT_AMPL_WIDTH - 1),
		2670 => to_unsigned(8296, LUT_AMPL_WIDTH - 1),
		2671 => to_unsigned(8300, LUT_AMPL_WIDTH - 1),
		2672 => to_unsigned(8303, LUT_AMPL_WIDTH - 1),
		2673 => to_unsigned(8306, LUT_AMPL_WIDTH - 1),
		2674 => to_unsigned(8309, LUT_AMPL_WIDTH - 1),
		2675 => to_unsigned(8312, LUT_AMPL_WIDTH - 1),
		2676 => to_unsigned(8315, LUT_AMPL_WIDTH - 1),
		2677 => to_unsigned(8318, LUT_AMPL_WIDTH - 1),
		2678 => to_unsigned(8321, LUT_AMPL_WIDTH - 1),
		2679 => to_unsigned(8324, LUT_AMPL_WIDTH - 1),
		2680 => to_unsigned(8327, LUT_AMPL_WIDTH - 1),
		2681 => to_unsigned(8330, LUT_AMPL_WIDTH - 1),
		2682 => to_unsigned(8333, LUT_AMPL_WIDTH - 1),
		2683 => to_unsigned(8336, LUT_AMPL_WIDTH - 1),
		2684 => to_unsigned(8339, LUT_AMPL_WIDTH - 1),
		2685 => to_unsigned(8342, LUT_AMPL_WIDTH - 1),
		2686 => to_unsigned(8345, LUT_AMPL_WIDTH - 1),
		2687 => to_unsigned(8348, LUT_AMPL_WIDTH - 1),
		2688 => to_unsigned(8351, LUT_AMPL_WIDTH - 1),
		2689 => to_unsigned(8354, LUT_AMPL_WIDTH - 1),
		2690 => to_unsigned(8357, LUT_AMPL_WIDTH - 1),
		2691 => to_unsigned(8360, LUT_AMPL_WIDTH - 1),
		2692 => to_unsigned(8363, LUT_AMPL_WIDTH - 1),
		2693 => to_unsigned(8366, LUT_AMPL_WIDTH - 1),
		2694 => to_unsigned(8369, LUT_AMPL_WIDTH - 1),
		2695 => to_unsigned(8372, LUT_AMPL_WIDTH - 1),
		2696 => to_unsigned(8375, LUT_AMPL_WIDTH - 1),
		2697 => to_unsigned(8379, LUT_AMPL_WIDTH - 1),
		2698 => to_unsigned(8382, LUT_AMPL_WIDTH - 1),
		2699 => to_unsigned(8385, LUT_AMPL_WIDTH - 1),
		2700 => to_unsigned(8388, LUT_AMPL_WIDTH - 1),
		2701 => to_unsigned(8391, LUT_AMPL_WIDTH - 1),
		2702 => to_unsigned(8394, LUT_AMPL_WIDTH - 1),
		2703 => to_unsigned(8397, LUT_AMPL_WIDTH - 1),
		2704 => to_unsigned(8400, LUT_AMPL_WIDTH - 1),
		2705 => to_unsigned(8403, LUT_AMPL_WIDTH - 1),
		2706 => to_unsigned(8406, LUT_AMPL_WIDTH - 1),
		2707 => to_unsigned(8409, LUT_AMPL_WIDTH - 1),
		2708 => to_unsigned(8412, LUT_AMPL_WIDTH - 1),
		2709 => to_unsigned(8415, LUT_AMPL_WIDTH - 1),
		2710 => to_unsigned(8418, LUT_AMPL_WIDTH - 1),
		2711 => to_unsigned(8421, LUT_AMPL_WIDTH - 1),
		2712 => to_unsigned(8424, LUT_AMPL_WIDTH - 1),
		2713 => to_unsigned(8427, LUT_AMPL_WIDTH - 1),
		2714 => to_unsigned(8430, LUT_AMPL_WIDTH - 1),
		2715 => to_unsigned(8433, LUT_AMPL_WIDTH - 1),
		2716 => to_unsigned(8436, LUT_AMPL_WIDTH - 1),
		2717 => to_unsigned(8439, LUT_AMPL_WIDTH - 1),
		2718 => to_unsigned(8442, LUT_AMPL_WIDTH - 1),
		2719 => to_unsigned(8445, LUT_AMPL_WIDTH - 1),
		2720 => to_unsigned(8448, LUT_AMPL_WIDTH - 1),
		2721 => to_unsigned(8451, LUT_AMPL_WIDTH - 1),
		2722 => to_unsigned(8454, LUT_AMPL_WIDTH - 1),
		2723 => to_unsigned(8457, LUT_AMPL_WIDTH - 1),
		2724 => to_unsigned(8460, LUT_AMPL_WIDTH - 1),
		2725 => to_unsigned(8464, LUT_AMPL_WIDTH - 1),
		2726 => to_unsigned(8467, LUT_AMPL_WIDTH - 1),
		2727 => to_unsigned(8470, LUT_AMPL_WIDTH - 1),
		2728 => to_unsigned(8473, LUT_AMPL_WIDTH - 1),
		2729 => to_unsigned(8476, LUT_AMPL_WIDTH - 1),
		2730 => to_unsigned(8479, LUT_AMPL_WIDTH - 1),
		2731 => to_unsigned(8482, LUT_AMPL_WIDTH - 1),
		2732 => to_unsigned(8485, LUT_AMPL_WIDTH - 1),
		2733 => to_unsigned(8488, LUT_AMPL_WIDTH - 1),
		2734 => to_unsigned(8491, LUT_AMPL_WIDTH - 1),
		2735 => to_unsigned(8494, LUT_AMPL_WIDTH - 1),
		2736 => to_unsigned(8497, LUT_AMPL_WIDTH - 1),
		2737 => to_unsigned(8500, LUT_AMPL_WIDTH - 1),
		2738 => to_unsigned(8503, LUT_AMPL_WIDTH - 1),
		2739 => to_unsigned(8506, LUT_AMPL_WIDTH - 1),
		2740 => to_unsigned(8509, LUT_AMPL_WIDTH - 1),
		2741 => to_unsigned(8512, LUT_AMPL_WIDTH - 1),
		2742 => to_unsigned(8515, LUT_AMPL_WIDTH - 1),
		2743 => to_unsigned(8518, LUT_AMPL_WIDTH - 1),
		2744 => to_unsigned(8521, LUT_AMPL_WIDTH - 1),
		2745 => to_unsigned(8524, LUT_AMPL_WIDTH - 1),
		2746 => to_unsigned(8527, LUT_AMPL_WIDTH - 1),
		2747 => to_unsigned(8530, LUT_AMPL_WIDTH - 1),
		2748 => to_unsigned(8533, LUT_AMPL_WIDTH - 1),
		2749 => to_unsigned(8536, LUT_AMPL_WIDTH - 1),
		2750 => to_unsigned(8539, LUT_AMPL_WIDTH - 1),
		2751 => to_unsigned(8542, LUT_AMPL_WIDTH - 1),
		2752 => to_unsigned(8545, LUT_AMPL_WIDTH - 1),
		2753 => to_unsigned(8548, LUT_AMPL_WIDTH - 1),
		2754 => to_unsigned(8552, LUT_AMPL_WIDTH - 1),
		2755 => to_unsigned(8555, LUT_AMPL_WIDTH - 1),
		2756 => to_unsigned(8558, LUT_AMPL_WIDTH - 1),
		2757 => to_unsigned(8561, LUT_AMPL_WIDTH - 1),
		2758 => to_unsigned(8564, LUT_AMPL_WIDTH - 1),
		2759 => to_unsigned(8567, LUT_AMPL_WIDTH - 1),
		2760 => to_unsigned(8570, LUT_AMPL_WIDTH - 1),
		2761 => to_unsigned(8573, LUT_AMPL_WIDTH - 1),
		2762 => to_unsigned(8576, LUT_AMPL_WIDTH - 1),
		2763 => to_unsigned(8579, LUT_AMPL_WIDTH - 1),
		2764 => to_unsigned(8582, LUT_AMPL_WIDTH - 1),
		2765 => to_unsigned(8585, LUT_AMPL_WIDTH - 1),
		2766 => to_unsigned(8588, LUT_AMPL_WIDTH - 1),
		2767 => to_unsigned(8591, LUT_AMPL_WIDTH - 1),
		2768 => to_unsigned(8594, LUT_AMPL_WIDTH - 1),
		2769 => to_unsigned(8597, LUT_AMPL_WIDTH - 1),
		2770 => to_unsigned(8600, LUT_AMPL_WIDTH - 1),
		2771 => to_unsigned(8603, LUT_AMPL_WIDTH - 1),
		2772 => to_unsigned(8606, LUT_AMPL_WIDTH - 1),
		2773 => to_unsigned(8609, LUT_AMPL_WIDTH - 1),
		2774 => to_unsigned(8612, LUT_AMPL_WIDTH - 1),
		2775 => to_unsigned(8615, LUT_AMPL_WIDTH - 1),
		2776 => to_unsigned(8618, LUT_AMPL_WIDTH - 1),
		2777 => to_unsigned(8621, LUT_AMPL_WIDTH - 1),
		2778 => to_unsigned(8624, LUT_AMPL_WIDTH - 1),
		2779 => to_unsigned(8627, LUT_AMPL_WIDTH - 1),
		2780 => to_unsigned(8630, LUT_AMPL_WIDTH - 1),
		2781 => to_unsigned(8633, LUT_AMPL_WIDTH - 1),
		2782 => to_unsigned(8636, LUT_AMPL_WIDTH - 1),
		2783 => to_unsigned(8639, LUT_AMPL_WIDTH - 1),
		2784 => to_unsigned(8642, LUT_AMPL_WIDTH - 1),
		2785 => to_unsigned(8645, LUT_AMPL_WIDTH - 1),
		2786 => to_unsigned(8649, LUT_AMPL_WIDTH - 1),
		2787 => to_unsigned(8652, LUT_AMPL_WIDTH - 1),
		2788 => to_unsigned(8655, LUT_AMPL_WIDTH - 1),
		2789 => to_unsigned(8658, LUT_AMPL_WIDTH - 1),
		2790 => to_unsigned(8661, LUT_AMPL_WIDTH - 1),
		2791 => to_unsigned(8664, LUT_AMPL_WIDTH - 1),
		2792 => to_unsigned(8667, LUT_AMPL_WIDTH - 1),
		2793 => to_unsigned(8670, LUT_AMPL_WIDTH - 1),
		2794 => to_unsigned(8673, LUT_AMPL_WIDTH - 1),
		2795 => to_unsigned(8676, LUT_AMPL_WIDTH - 1),
		2796 => to_unsigned(8679, LUT_AMPL_WIDTH - 1),
		2797 => to_unsigned(8682, LUT_AMPL_WIDTH - 1),
		2798 => to_unsigned(8685, LUT_AMPL_WIDTH - 1),
		2799 => to_unsigned(8688, LUT_AMPL_WIDTH - 1),
		2800 => to_unsigned(8691, LUT_AMPL_WIDTH - 1),
		2801 => to_unsigned(8694, LUT_AMPL_WIDTH - 1),
		2802 => to_unsigned(8697, LUT_AMPL_WIDTH - 1),
		2803 => to_unsigned(8700, LUT_AMPL_WIDTH - 1),
		2804 => to_unsigned(8703, LUT_AMPL_WIDTH - 1),
		2805 => to_unsigned(8706, LUT_AMPL_WIDTH - 1),
		2806 => to_unsigned(8709, LUT_AMPL_WIDTH - 1),
		2807 => to_unsigned(8712, LUT_AMPL_WIDTH - 1),
		2808 => to_unsigned(8715, LUT_AMPL_WIDTH - 1),
		2809 => to_unsigned(8718, LUT_AMPL_WIDTH - 1),
		2810 => to_unsigned(8721, LUT_AMPL_WIDTH - 1),
		2811 => to_unsigned(8724, LUT_AMPL_WIDTH - 1),
		2812 => to_unsigned(8727, LUT_AMPL_WIDTH - 1),
		2813 => to_unsigned(8730, LUT_AMPL_WIDTH - 1),
		2814 => to_unsigned(8733, LUT_AMPL_WIDTH - 1),
		2815 => to_unsigned(8736, LUT_AMPL_WIDTH - 1),
		2816 => to_unsigned(8739, LUT_AMPL_WIDTH - 1),
		2817 => to_unsigned(8742, LUT_AMPL_WIDTH - 1),
		2818 => to_unsigned(8745, LUT_AMPL_WIDTH - 1),
		2819 => to_unsigned(8748, LUT_AMPL_WIDTH - 1),
		2820 => to_unsigned(8751, LUT_AMPL_WIDTH - 1),
		2821 => to_unsigned(8755, LUT_AMPL_WIDTH - 1),
		2822 => to_unsigned(8758, LUT_AMPL_WIDTH - 1),
		2823 => to_unsigned(8761, LUT_AMPL_WIDTH - 1),
		2824 => to_unsigned(8764, LUT_AMPL_WIDTH - 1),
		2825 => to_unsigned(8767, LUT_AMPL_WIDTH - 1),
		2826 => to_unsigned(8770, LUT_AMPL_WIDTH - 1),
		2827 => to_unsigned(8773, LUT_AMPL_WIDTH - 1),
		2828 => to_unsigned(8776, LUT_AMPL_WIDTH - 1),
		2829 => to_unsigned(8779, LUT_AMPL_WIDTH - 1),
		2830 => to_unsigned(8782, LUT_AMPL_WIDTH - 1),
		2831 => to_unsigned(8785, LUT_AMPL_WIDTH - 1),
		2832 => to_unsigned(8788, LUT_AMPL_WIDTH - 1),
		2833 => to_unsigned(8791, LUT_AMPL_WIDTH - 1),
		2834 => to_unsigned(8794, LUT_AMPL_WIDTH - 1),
		2835 => to_unsigned(8797, LUT_AMPL_WIDTH - 1),
		2836 => to_unsigned(8800, LUT_AMPL_WIDTH - 1),
		2837 => to_unsigned(8803, LUT_AMPL_WIDTH - 1),
		2838 => to_unsigned(8806, LUT_AMPL_WIDTH - 1),
		2839 => to_unsigned(8809, LUT_AMPL_WIDTH - 1),
		2840 => to_unsigned(8812, LUT_AMPL_WIDTH - 1),
		2841 => to_unsigned(8815, LUT_AMPL_WIDTH - 1),
		2842 => to_unsigned(8818, LUT_AMPL_WIDTH - 1),
		2843 => to_unsigned(8821, LUT_AMPL_WIDTH - 1),
		2844 => to_unsigned(8824, LUT_AMPL_WIDTH - 1),
		2845 => to_unsigned(8827, LUT_AMPL_WIDTH - 1),
		2846 => to_unsigned(8830, LUT_AMPL_WIDTH - 1),
		2847 => to_unsigned(8833, LUT_AMPL_WIDTH - 1),
		2848 => to_unsigned(8836, LUT_AMPL_WIDTH - 1),
		2849 => to_unsigned(8839, LUT_AMPL_WIDTH - 1),
		2850 => to_unsigned(8842, LUT_AMPL_WIDTH - 1),
		2851 => to_unsigned(8845, LUT_AMPL_WIDTH - 1),
		2852 => to_unsigned(8848, LUT_AMPL_WIDTH - 1),
		2853 => to_unsigned(8851, LUT_AMPL_WIDTH - 1),
		2854 => to_unsigned(8854, LUT_AMPL_WIDTH - 1),
		2855 => to_unsigned(8857, LUT_AMPL_WIDTH - 1),
		2856 => to_unsigned(8860, LUT_AMPL_WIDTH - 1),
		2857 => to_unsigned(8863, LUT_AMPL_WIDTH - 1),
		2858 => to_unsigned(8866, LUT_AMPL_WIDTH - 1),
		2859 => to_unsigned(8869, LUT_AMPL_WIDTH - 1),
		2860 => to_unsigned(8873, LUT_AMPL_WIDTH - 1),
		2861 => to_unsigned(8876, LUT_AMPL_WIDTH - 1),
		2862 => to_unsigned(8879, LUT_AMPL_WIDTH - 1),
		2863 => to_unsigned(8882, LUT_AMPL_WIDTH - 1),
		2864 => to_unsigned(8885, LUT_AMPL_WIDTH - 1),
		2865 => to_unsigned(8888, LUT_AMPL_WIDTH - 1),
		2866 => to_unsigned(8891, LUT_AMPL_WIDTH - 1),
		2867 => to_unsigned(8894, LUT_AMPL_WIDTH - 1),
		2868 => to_unsigned(8897, LUT_AMPL_WIDTH - 1),
		2869 => to_unsigned(8900, LUT_AMPL_WIDTH - 1),
		2870 => to_unsigned(8903, LUT_AMPL_WIDTH - 1),
		2871 => to_unsigned(8906, LUT_AMPL_WIDTH - 1),
		2872 => to_unsigned(8909, LUT_AMPL_WIDTH - 1),
		2873 => to_unsigned(8912, LUT_AMPL_WIDTH - 1),
		2874 => to_unsigned(8915, LUT_AMPL_WIDTH - 1),
		2875 => to_unsigned(8918, LUT_AMPL_WIDTH - 1),
		2876 => to_unsigned(8921, LUT_AMPL_WIDTH - 1),
		2877 => to_unsigned(8924, LUT_AMPL_WIDTH - 1),
		2878 => to_unsigned(8927, LUT_AMPL_WIDTH - 1),
		2879 => to_unsigned(8930, LUT_AMPL_WIDTH - 1),
		2880 => to_unsigned(8933, LUT_AMPL_WIDTH - 1),
		2881 => to_unsigned(8936, LUT_AMPL_WIDTH - 1),
		2882 => to_unsigned(8939, LUT_AMPL_WIDTH - 1),
		2883 => to_unsigned(8942, LUT_AMPL_WIDTH - 1),
		2884 => to_unsigned(8945, LUT_AMPL_WIDTH - 1),
		2885 => to_unsigned(8948, LUT_AMPL_WIDTH - 1),
		2886 => to_unsigned(8951, LUT_AMPL_WIDTH - 1),
		2887 => to_unsigned(8954, LUT_AMPL_WIDTH - 1),
		2888 => to_unsigned(8957, LUT_AMPL_WIDTH - 1),
		2889 => to_unsigned(8960, LUT_AMPL_WIDTH - 1),
		2890 => to_unsigned(8963, LUT_AMPL_WIDTH - 1),
		2891 => to_unsigned(8966, LUT_AMPL_WIDTH - 1),
		2892 => to_unsigned(8969, LUT_AMPL_WIDTH - 1),
		2893 => to_unsigned(8972, LUT_AMPL_WIDTH - 1),
		2894 => to_unsigned(8975, LUT_AMPL_WIDTH - 1),
		2895 => to_unsigned(8978, LUT_AMPL_WIDTH - 1),
		2896 => to_unsigned(8981, LUT_AMPL_WIDTH - 1),
		2897 => to_unsigned(8984, LUT_AMPL_WIDTH - 1),
		2898 => to_unsigned(8987, LUT_AMPL_WIDTH - 1),
		2899 => to_unsigned(8990, LUT_AMPL_WIDTH - 1),
		2900 => to_unsigned(8993, LUT_AMPL_WIDTH - 1),
		2901 => to_unsigned(8996, LUT_AMPL_WIDTH - 1),
		2902 => to_unsigned(8999, LUT_AMPL_WIDTH - 1),
		2903 => to_unsigned(9002, LUT_AMPL_WIDTH - 1),
		2904 => to_unsigned(9006, LUT_AMPL_WIDTH - 1),
		2905 => to_unsigned(9009, LUT_AMPL_WIDTH - 1),
		2906 => to_unsigned(9012, LUT_AMPL_WIDTH - 1),
		2907 => to_unsigned(9015, LUT_AMPL_WIDTH - 1),
		2908 => to_unsigned(9018, LUT_AMPL_WIDTH - 1),
		2909 => to_unsigned(9021, LUT_AMPL_WIDTH - 1),
		2910 => to_unsigned(9024, LUT_AMPL_WIDTH - 1),
		2911 => to_unsigned(9027, LUT_AMPL_WIDTH - 1),
		2912 => to_unsigned(9030, LUT_AMPL_WIDTH - 1),
		2913 => to_unsigned(9033, LUT_AMPL_WIDTH - 1),
		2914 => to_unsigned(9036, LUT_AMPL_WIDTH - 1),
		2915 => to_unsigned(9039, LUT_AMPL_WIDTH - 1),
		2916 => to_unsigned(9042, LUT_AMPL_WIDTH - 1),
		2917 => to_unsigned(9045, LUT_AMPL_WIDTH - 1),
		2918 => to_unsigned(9048, LUT_AMPL_WIDTH - 1),
		2919 => to_unsigned(9051, LUT_AMPL_WIDTH - 1),
		2920 => to_unsigned(9054, LUT_AMPL_WIDTH - 1),
		2921 => to_unsigned(9057, LUT_AMPL_WIDTH - 1),
		2922 => to_unsigned(9060, LUT_AMPL_WIDTH - 1),
		2923 => to_unsigned(9063, LUT_AMPL_WIDTH - 1),
		2924 => to_unsigned(9066, LUT_AMPL_WIDTH - 1),
		2925 => to_unsigned(9069, LUT_AMPL_WIDTH - 1),
		2926 => to_unsigned(9072, LUT_AMPL_WIDTH - 1),
		2927 => to_unsigned(9075, LUT_AMPL_WIDTH - 1),
		2928 => to_unsigned(9078, LUT_AMPL_WIDTH - 1),
		2929 => to_unsigned(9081, LUT_AMPL_WIDTH - 1),
		2930 => to_unsigned(9084, LUT_AMPL_WIDTH - 1),
		2931 => to_unsigned(9087, LUT_AMPL_WIDTH - 1),
		2932 => to_unsigned(9090, LUT_AMPL_WIDTH - 1),
		2933 => to_unsigned(9093, LUT_AMPL_WIDTH - 1),
		2934 => to_unsigned(9096, LUT_AMPL_WIDTH - 1),
		2935 => to_unsigned(9099, LUT_AMPL_WIDTH - 1),
		2936 => to_unsigned(9102, LUT_AMPL_WIDTH - 1),
		2937 => to_unsigned(9105, LUT_AMPL_WIDTH - 1),
		2938 => to_unsigned(9108, LUT_AMPL_WIDTH - 1),
		2939 => to_unsigned(9111, LUT_AMPL_WIDTH - 1),
		2940 => to_unsigned(9114, LUT_AMPL_WIDTH - 1),
		2941 => to_unsigned(9117, LUT_AMPL_WIDTH - 1),
		2942 => to_unsigned(9120, LUT_AMPL_WIDTH - 1),
		2943 => to_unsigned(9123, LUT_AMPL_WIDTH - 1),
		2944 => to_unsigned(9126, LUT_AMPL_WIDTH - 1),
		2945 => to_unsigned(9129, LUT_AMPL_WIDTH - 1),
		2946 => to_unsigned(9132, LUT_AMPL_WIDTH - 1),
		2947 => to_unsigned(9135, LUT_AMPL_WIDTH - 1),
		2948 => to_unsigned(9138, LUT_AMPL_WIDTH - 1),
		2949 => to_unsigned(9141, LUT_AMPL_WIDTH - 1),
		2950 => to_unsigned(9144, LUT_AMPL_WIDTH - 1),
		2951 => to_unsigned(9147, LUT_AMPL_WIDTH - 1),
		2952 => to_unsigned(9150, LUT_AMPL_WIDTH - 1),
		2953 => to_unsigned(9153, LUT_AMPL_WIDTH - 1),
		2954 => to_unsigned(9156, LUT_AMPL_WIDTH - 1),
		2955 => to_unsigned(9159, LUT_AMPL_WIDTH - 1),
		2956 => to_unsigned(9162, LUT_AMPL_WIDTH - 1),
		2957 => to_unsigned(9165, LUT_AMPL_WIDTH - 1),
		2958 => to_unsigned(9168, LUT_AMPL_WIDTH - 1),
		2959 => to_unsigned(9172, LUT_AMPL_WIDTH - 1),
		2960 => to_unsigned(9175, LUT_AMPL_WIDTH - 1),
		2961 => to_unsigned(9178, LUT_AMPL_WIDTH - 1),
		2962 => to_unsigned(9181, LUT_AMPL_WIDTH - 1),
		2963 => to_unsigned(9184, LUT_AMPL_WIDTH - 1),
		2964 => to_unsigned(9187, LUT_AMPL_WIDTH - 1),
		2965 => to_unsigned(9190, LUT_AMPL_WIDTH - 1),
		2966 => to_unsigned(9193, LUT_AMPL_WIDTH - 1),
		2967 => to_unsigned(9196, LUT_AMPL_WIDTH - 1),
		2968 => to_unsigned(9199, LUT_AMPL_WIDTH - 1),
		2969 => to_unsigned(9202, LUT_AMPL_WIDTH - 1),
		2970 => to_unsigned(9205, LUT_AMPL_WIDTH - 1),
		2971 => to_unsigned(9208, LUT_AMPL_WIDTH - 1),
		2972 => to_unsigned(9211, LUT_AMPL_WIDTH - 1),
		2973 => to_unsigned(9214, LUT_AMPL_WIDTH - 1),
		2974 => to_unsigned(9217, LUT_AMPL_WIDTH - 1),
		2975 => to_unsigned(9220, LUT_AMPL_WIDTH - 1),
		2976 => to_unsigned(9223, LUT_AMPL_WIDTH - 1),
		2977 => to_unsigned(9226, LUT_AMPL_WIDTH - 1),
		2978 => to_unsigned(9229, LUT_AMPL_WIDTH - 1),
		2979 => to_unsigned(9232, LUT_AMPL_WIDTH - 1),
		2980 => to_unsigned(9235, LUT_AMPL_WIDTH - 1),
		2981 => to_unsigned(9238, LUT_AMPL_WIDTH - 1),
		2982 => to_unsigned(9241, LUT_AMPL_WIDTH - 1),
		2983 => to_unsigned(9244, LUT_AMPL_WIDTH - 1),
		2984 => to_unsigned(9247, LUT_AMPL_WIDTH - 1),
		2985 => to_unsigned(9250, LUT_AMPL_WIDTH - 1),
		2986 => to_unsigned(9253, LUT_AMPL_WIDTH - 1),
		2987 => to_unsigned(9256, LUT_AMPL_WIDTH - 1),
		2988 => to_unsigned(9259, LUT_AMPL_WIDTH - 1),
		2989 => to_unsigned(9262, LUT_AMPL_WIDTH - 1),
		2990 => to_unsigned(9265, LUT_AMPL_WIDTH - 1),
		2991 => to_unsigned(9268, LUT_AMPL_WIDTH - 1),
		2992 => to_unsigned(9271, LUT_AMPL_WIDTH - 1),
		2993 => to_unsigned(9274, LUT_AMPL_WIDTH - 1),
		2994 => to_unsigned(9277, LUT_AMPL_WIDTH - 1),
		2995 => to_unsigned(9280, LUT_AMPL_WIDTH - 1),
		2996 => to_unsigned(9283, LUT_AMPL_WIDTH - 1),
		2997 => to_unsigned(9286, LUT_AMPL_WIDTH - 1),
		2998 => to_unsigned(9289, LUT_AMPL_WIDTH - 1),
		2999 => to_unsigned(9292, LUT_AMPL_WIDTH - 1),
		3000 => to_unsigned(9295, LUT_AMPL_WIDTH - 1),
		3001 => to_unsigned(9298, LUT_AMPL_WIDTH - 1),
		3002 => to_unsigned(9301, LUT_AMPL_WIDTH - 1),
		3003 => to_unsigned(9304, LUT_AMPL_WIDTH - 1),
		3004 => to_unsigned(9307, LUT_AMPL_WIDTH - 1),
		3005 => to_unsigned(9310, LUT_AMPL_WIDTH - 1),
		3006 => to_unsigned(9313, LUT_AMPL_WIDTH - 1),
		3007 => to_unsigned(9316, LUT_AMPL_WIDTH - 1),
		3008 => to_unsigned(9319, LUT_AMPL_WIDTH - 1),
		3009 => to_unsigned(9322, LUT_AMPL_WIDTH - 1),
		3010 => to_unsigned(9325, LUT_AMPL_WIDTH - 1),
		3011 => to_unsigned(9328, LUT_AMPL_WIDTH - 1),
		3012 => to_unsigned(9331, LUT_AMPL_WIDTH - 1),
		3013 => to_unsigned(9334, LUT_AMPL_WIDTH - 1),
		3014 => to_unsigned(9337, LUT_AMPL_WIDTH - 1),
		3015 => to_unsigned(9340, LUT_AMPL_WIDTH - 1),
		3016 => to_unsigned(9343, LUT_AMPL_WIDTH - 1),
		3017 => to_unsigned(9346, LUT_AMPL_WIDTH - 1),
		3018 => to_unsigned(9349, LUT_AMPL_WIDTH - 1),
		3019 => to_unsigned(9352, LUT_AMPL_WIDTH - 1),
		3020 => to_unsigned(9355, LUT_AMPL_WIDTH - 1),
		3021 => to_unsigned(9358, LUT_AMPL_WIDTH - 1),
		3022 => to_unsigned(9361, LUT_AMPL_WIDTH - 1),
		3023 => to_unsigned(9364, LUT_AMPL_WIDTH - 1),
		3024 => to_unsigned(9367, LUT_AMPL_WIDTH - 1),
		3025 => to_unsigned(9370, LUT_AMPL_WIDTH - 1),
		3026 => to_unsigned(9373, LUT_AMPL_WIDTH - 1),
		3027 => to_unsigned(9376, LUT_AMPL_WIDTH - 1),
		3028 => to_unsigned(9379, LUT_AMPL_WIDTH - 1),
		3029 => to_unsigned(9382, LUT_AMPL_WIDTH - 1),
		3030 => to_unsigned(9385, LUT_AMPL_WIDTH - 1),
		3031 => to_unsigned(9388, LUT_AMPL_WIDTH - 1),
		3032 => to_unsigned(9391, LUT_AMPL_WIDTH - 1),
		3033 => to_unsigned(9394, LUT_AMPL_WIDTH - 1),
		3034 => to_unsigned(9397, LUT_AMPL_WIDTH - 1),
		3035 => to_unsigned(9400, LUT_AMPL_WIDTH - 1),
		3036 => to_unsigned(9403, LUT_AMPL_WIDTH - 1),
		3037 => to_unsigned(9406, LUT_AMPL_WIDTH - 1),
		3038 => to_unsigned(9409, LUT_AMPL_WIDTH - 1),
		3039 => to_unsigned(9413, LUT_AMPL_WIDTH - 1),
		3040 => to_unsigned(9416, LUT_AMPL_WIDTH - 1),
		3041 => to_unsigned(9419, LUT_AMPL_WIDTH - 1),
		3042 => to_unsigned(9422, LUT_AMPL_WIDTH - 1),
		3043 => to_unsigned(9425, LUT_AMPL_WIDTH - 1),
		3044 => to_unsigned(9428, LUT_AMPL_WIDTH - 1),
		3045 => to_unsigned(9431, LUT_AMPL_WIDTH - 1),
		3046 => to_unsigned(9434, LUT_AMPL_WIDTH - 1),
		3047 => to_unsigned(9437, LUT_AMPL_WIDTH - 1),
		3048 => to_unsigned(9440, LUT_AMPL_WIDTH - 1),
		3049 => to_unsigned(9443, LUT_AMPL_WIDTH - 1),
		3050 => to_unsigned(9446, LUT_AMPL_WIDTH - 1),
		3051 => to_unsigned(9449, LUT_AMPL_WIDTH - 1),
		3052 => to_unsigned(9452, LUT_AMPL_WIDTH - 1),
		3053 => to_unsigned(9455, LUT_AMPL_WIDTH - 1),
		3054 => to_unsigned(9458, LUT_AMPL_WIDTH - 1),
		3055 => to_unsigned(9461, LUT_AMPL_WIDTH - 1),
		3056 => to_unsigned(9464, LUT_AMPL_WIDTH - 1),
		3057 => to_unsigned(9467, LUT_AMPL_WIDTH - 1),
		3058 => to_unsigned(9470, LUT_AMPL_WIDTH - 1),
		3059 => to_unsigned(9473, LUT_AMPL_WIDTH - 1),
		3060 => to_unsigned(9476, LUT_AMPL_WIDTH - 1),
		3061 => to_unsigned(9479, LUT_AMPL_WIDTH - 1),
		3062 => to_unsigned(9482, LUT_AMPL_WIDTH - 1),
		3063 => to_unsigned(9485, LUT_AMPL_WIDTH - 1),
		3064 => to_unsigned(9488, LUT_AMPL_WIDTH - 1),
		3065 => to_unsigned(9491, LUT_AMPL_WIDTH - 1),
		3066 => to_unsigned(9494, LUT_AMPL_WIDTH - 1),
		3067 => to_unsigned(9497, LUT_AMPL_WIDTH - 1),
		3068 => to_unsigned(9500, LUT_AMPL_WIDTH - 1),
		3069 => to_unsigned(9503, LUT_AMPL_WIDTH - 1),
		3070 => to_unsigned(9506, LUT_AMPL_WIDTH - 1),
		3071 => to_unsigned(9509, LUT_AMPL_WIDTH - 1),
		3072 => to_unsigned(9512, LUT_AMPL_WIDTH - 1),
		3073 => to_unsigned(9515, LUT_AMPL_WIDTH - 1),
		3074 => to_unsigned(9518, LUT_AMPL_WIDTH - 1),
		3075 => to_unsigned(9521, LUT_AMPL_WIDTH - 1),
		3076 => to_unsigned(9524, LUT_AMPL_WIDTH - 1),
		3077 => to_unsigned(9527, LUT_AMPL_WIDTH - 1),
		3078 => to_unsigned(9530, LUT_AMPL_WIDTH - 1),
		3079 => to_unsigned(9533, LUT_AMPL_WIDTH - 1),
		3080 => to_unsigned(9536, LUT_AMPL_WIDTH - 1),
		3081 => to_unsigned(9539, LUT_AMPL_WIDTH - 1),
		3082 => to_unsigned(9542, LUT_AMPL_WIDTH - 1),
		3083 => to_unsigned(9545, LUT_AMPL_WIDTH - 1),
		3084 => to_unsigned(9548, LUT_AMPL_WIDTH - 1),
		3085 => to_unsigned(9551, LUT_AMPL_WIDTH - 1),
		3086 => to_unsigned(9554, LUT_AMPL_WIDTH - 1),
		3087 => to_unsigned(9557, LUT_AMPL_WIDTH - 1),
		3088 => to_unsigned(9560, LUT_AMPL_WIDTH - 1),
		3089 => to_unsigned(9563, LUT_AMPL_WIDTH - 1),
		3090 => to_unsigned(9566, LUT_AMPL_WIDTH - 1),
		3091 => to_unsigned(9569, LUT_AMPL_WIDTH - 1),
		3092 => to_unsigned(9572, LUT_AMPL_WIDTH - 1),
		3093 => to_unsigned(9575, LUT_AMPL_WIDTH - 1),
		3094 => to_unsigned(9578, LUT_AMPL_WIDTH - 1),
		3095 => to_unsigned(9581, LUT_AMPL_WIDTH - 1),
		3096 => to_unsigned(9584, LUT_AMPL_WIDTH - 1),
		3097 => to_unsigned(9587, LUT_AMPL_WIDTH - 1),
		3098 => to_unsigned(9590, LUT_AMPL_WIDTH - 1),
		3099 => to_unsigned(9593, LUT_AMPL_WIDTH - 1),
		3100 => to_unsigned(9596, LUT_AMPL_WIDTH - 1),
		3101 => to_unsigned(9599, LUT_AMPL_WIDTH - 1),
		3102 => to_unsigned(9602, LUT_AMPL_WIDTH - 1),
		3103 => to_unsigned(9605, LUT_AMPL_WIDTH - 1),
		3104 => to_unsigned(9608, LUT_AMPL_WIDTH - 1),
		3105 => to_unsigned(9611, LUT_AMPL_WIDTH - 1),
		3106 => to_unsigned(9614, LUT_AMPL_WIDTH - 1),
		3107 => to_unsigned(9617, LUT_AMPL_WIDTH - 1),
		3108 => to_unsigned(9620, LUT_AMPL_WIDTH - 1),
		3109 => to_unsigned(9623, LUT_AMPL_WIDTH - 1),
		3110 => to_unsigned(9626, LUT_AMPL_WIDTH - 1),
		3111 => to_unsigned(9629, LUT_AMPL_WIDTH - 1),
		3112 => to_unsigned(9632, LUT_AMPL_WIDTH - 1),
		3113 => to_unsigned(9635, LUT_AMPL_WIDTH - 1),
		3114 => to_unsigned(9638, LUT_AMPL_WIDTH - 1),
		3115 => to_unsigned(9641, LUT_AMPL_WIDTH - 1),
		3116 => to_unsigned(9644, LUT_AMPL_WIDTH - 1),
		3117 => to_unsigned(9647, LUT_AMPL_WIDTH - 1),
		3118 => to_unsigned(9650, LUT_AMPL_WIDTH - 1),
		3119 => to_unsigned(9653, LUT_AMPL_WIDTH - 1),
		3120 => to_unsigned(9656, LUT_AMPL_WIDTH - 1),
		3121 => to_unsigned(9659, LUT_AMPL_WIDTH - 1),
		3122 => to_unsigned(9662, LUT_AMPL_WIDTH - 1),
		3123 => to_unsigned(9665, LUT_AMPL_WIDTH - 1),
		3124 => to_unsigned(9668, LUT_AMPL_WIDTH - 1),
		3125 => to_unsigned(9671, LUT_AMPL_WIDTH - 1),
		3126 => to_unsigned(9674, LUT_AMPL_WIDTH - 1),
		3127 => to_unsigned(9677, LUT_AMPL_WIDTH - 1),
		3128 => to_unsigned(9680, LUT_AMPL_WIDTH - 1),
		3129 => to_unsigned(9683, LUT_AMPL_WIDTH - 1),
		3130 => to_unsigned(9686, LUT_AMPL_WIDTH - 1),
		3131 => to_unsigned(9689, LUT_AMPL_WIDTH - 1),
		3132 => to_unsigned(9692, LUT_AMPL_WIDTH - 1),
		3133 => to_unsigned(9695, LUT_AMPL_WIDTH - 1),
		3134 => to_unsigned(9698, LUT_AMPL_WIDTH - 1),
		3135 => to_unsigned(9701, LUT_AMPL_WIDTH - 1),
		3136 => to_unsigned(9704, LUT_AMPL_WIDTH - 1),
		3137 => to_unsigned(9707, LUT_AMPL_WIDTH - 1),
		3138 => to_unsigned(9710, LUT_AMPL_WIDTH - 1),
		3139 => to_unsigned(9713, LUT_AMPL_WIDTH - 1),
		3140 => to_unsigned(9716, LUT_AMPL_WIDTH - 1),
		3141 => to_unsigned(9719, LUT_AMPL_WIDTH - 1),
		3142 => to_unsigned(9722, LUT_AMPL_WIDTH - 1),
		3143 => to_unsigned(9725, LUT_AMPL_WIDTH - 1),
		3144 => to_unsigned(9728, LUT_AMPL_WIDTH - 1),
		3145 => to_unsigned(9731, LUT_AMPL_WIDTH - 1),
		3146 => to_unsigned(9734, LUT_AMPL_WIDTH - 1),
		3147 => to_unsigned(9737, LUT_AMPL_WIDTH - 1),
		3148 => to_unsigned(9740, LUT_AMPL_WIDTH - 1),
		3149 => to_unsigned(9743, LUT_AMPL_WIDTH - 1),
		3150 => to_unsigned(9746, LUT_AMPL_WIDTH - 1),
		3151 => to_unsigned(9749, LUT_AMPL_WIDTH - 1),
		3152 => to_unsigned(9752, LUT_AMPL_WIDTH - 1),
		3153 => to_unsigned(9755, LUT_AMPL_WIDTH - 1),
		3154 => to_unsigned(9758, LUT_AMPL_WIDTH - 1),
		3155 => to_unsigned(9761, LUT_AMPL_WIDTH - 1),
		3156 => to_unsigned(9764, LUT_AMPL_WIDTH - 1),
		3157 => to_unsigned(9767, LUT_AMPL_WIDTH - 1),
		3158 => to_unsigned(9770, LUT_AMPL_WIDTH - 1),
		3159 => to_unsigned(9773, LUT_AMPL_WIDTH - 1),
		3160 => to_unsigned(9776, LUT_AMPL_WIDTH - 1),
		3161 => to_unsigned(9779, LUT_AMPL_WIDTH - 1),
		3162 => to_unsigned(9782, LUT_AMPL_WIDTH - 1),
		3163 => to_unsigned(9785, LUT_AMPL_WIDTH - 1),
		3164 => to_unsigned(9788, LUT_AMPL_WIDTH - 1),
		3165 => to_unsigned(9791, LUT_AMPL_WIDTH - 1),
		3166 => to_unsigned(9794, LUT_AMPL_WIDTH - 1),
		3167 => to_unsigned(9797, LUT_AMPL_WIDTH - 1),
		3168 => to_unsigned(9800, LUT_AMPL_WIDTH - 1),
		3169 => to_unsigned(9803, LUT_AMPL_WIDTH - 1),
		3170 => to_unsigned(9806, LUT_AMPL_WIDTH - 1),
		3171 => to_unsigned(9809, LUT_AMPL_WIDTH - 1),
		3172 => to_unsigned(9812, LUT_AMPL_WIDTH - 1),
		3173 => to_unsigned(9815, LUT_AMPL_WIDTH - 1),
		3174 => to_unsigned(9818, LUT_AMPL_WIDTH - 1),
		3175 => to_unsigned(9821, LUT_AMPL_WIDTH - 1),
		3176 => to_unsigned(9824, LUT_AMPL_WIDTH - 1),
		3177 => to_unsigned(9827, LUT_AMPL_WIDTH - 1),
		3178 => to_unsigned(9830, LUT_AMPL_WIDTH - 1),
		3179 => to_unsigned(9833, LUT_AMPL_WIDTH - 1),
		3180 => to_unsigned(9836, LUT_AMPL_WIDTH - 1),
		3181 => to_unsigned(9839, LUT_AMPL_WIDTH - 1),
		3182 => to_unsigned(9842, LUT_AMPL_WIDTH - 1),
		3183 => to_unsigned(9845, LUT_AMPL_WIDTH - 1),
		3184 => to_unsigned(9848, LUT_AMPL_WIDTH - 1),
		3185 => to_unsigned(9851, LUT_AMPL_WIDTH - 1),
		3186 => to_unsigned(9854, LUT_AMPL_WIDTH - 1),
		3187 => to_unsigned(9857, LUT_AMPL_WIDTH - 1),
		3188 => to_unsigned(9860, LUT_AMPL_WIDTH - 1),
		3189 => to_unsigned(9863, LUT_AMPL_WIDTH - 1),
		3190 => to_unsigned(9866, LUT_AMPL_WIDTH - 1),
		3191 => to_unsigned(9869, LUT_AMPL_WIDTH - 1),
		3192 => to_unsigned(9872, LUT_AMPL_WIDTH - 1),
		3193 => to_unsigned(9875, LUT_AMPL_WIDTH - 1),
		3194 => to_unsigned(9878, LUT_AMPL_WIDTH - 1),
		3195 => to_unsigned(9881, LUT_AMPL_WIDTH - 1),
		3196 => to_unsigned(9884, LUT_AMPL_WIDTH - 1),
		3197 => to_unsigned(9887, LUT_AMPL_WIDTH - 1),
		3198 => to_unsigned(9890, LUT_AMPL_WIDTH - 1),
		3199 => to_unsigned(9893, LUT_AMPL_WIDTH - 1),
		3200 => to_unsigned(9896, LUT_AMPL_WIDTH - 1),
		3201 => to_unsigned(9899, LUT_AMPL_WIDTH - 1),
		3202 => to_unsigned(9902, LUT_AMPL_WIDTH - 1),
		3203 => to_unsigned(9905, LUT_AMPL_WIDTH - 1),
		3204 => to_unsigned(9908, LUT_AMPL_WIDTH - 1),
		3205 => to_unsigned(9911, LUT_AMPL_WIDTH - 1),
		3206 => to_unsigned(9914, LUT_AMPL_WIDTH - 1),
		3207 => to_unsigned(9917, LUT_AMPL_WIDTH - 1),
		3208 => to_unsigned(9920, LUT_AMPL_WIDTH - 1),
		3209 => to_unsigned(9923, LUT_AMPL_WIDTH - 1),
		3210 => to_unsigned(9926, LUT_AMPL_WIDTH - 1),
		3211 => to_unsigned(9929, LUT_AMPL_WIDTH - 1),
		3212 => to_unsigned(9932, LUT_AMPL_WIDTH - 1),
		3213 => to_unsigned(9935, LUT_AMPL_WIDTH - 1),
		3214 => to_unsigned(9938, LUT_AMPL_WIDTH - 1),
		3215 => to_unsigned(9941, LUT_AMPL_WIDTH - 1),
		3216 => to_unsigned(9944, LUT_AMPL_WIDTH - 1),
		3217 => to_unsigned(9947, LUT_AMPL_WIDTH - 1),
		3218 => to_unsigned(9950, LUT_AMPL_WIDTH - 1),
		3219 => to_unsigned(9953, LUT_AMPL_WIDTH - 1),
		3220 => to_unsigned(9956, LUT_AMPL_WIDTH - 1),
		3221 => to_unsigned(9959, LUT_AMPL_WIDTH - 1),
		3222 => to_unsigned(9962, LUT_AMPL_WIDTH - 1),
		3223 => to_unsigned(9965, LUT_AMPL_WIDTH - 1),
		3224 => to_unsigned(9968, LUT_AMPL_WIDTH - 1),
		3225 => to_unsigned(9971, LUT_AMPL_WIDTH - 1),
		3226 => to_unsigned(9974, LUT_AMPL_WIDTH - 1),
		3227 => to_unsigned(9977, LUT_AMPL_WIDTH - 1),
		3228 => to_unsigned(9980, LUT_AMPL_WIDTH - 1),
		3229 => to_unsigned(9983, LUT_AMPL_WIDTH - 1),
		3230 => to_unsigned(9986, LUT_AMPL_WIDTH - 1),
		3231 => to_unsigned(9989, LUT_AMPL_WIDTH - 1),
		3232 => to_unsigned(9992, LUT_AMPL_WIDTH - 1),
		3233 => to_unsigned(9995, LUT_AMPL_WIDTH - 1),
		3234 => to_unsigned(9998, LUT_AMPL_WIDTH - 1),
		3235 => to_unsigned(10001, LUT_AMPL_WIDTH - 1),
		3236 => to_unsigned(10004, LUT_AMPL_WIDTH - 1),
		3237 => to_unsigned(10007, LUT_AMPL_WIDTH - 1),
		3238 => to_unsigned(10010, LUT_AMPL_WIDTH - 1),
		3239 => to_unsigned(10013, LUT_AMPL_WIDTH - 1),
		3240 => to_unsigned(10016, LUT_AMPL_WIDTH - 1),
		3241 => to_unsigned(10019, LUT_AMPL_WIDTH - 1),
		3242 => to_unsigned(10022, LUT_AMPL_WIDTH - 1),
		3243 => to_unsigned(10025, LUT_AMPL_WIDTH - 1),
		3244 => to_unsigned(10028, LUT_AMPL_WIDTH - 1),
		3245 => to_unsigned(10031, LUT_AMPL_WIDTH - 1),
		3246 => to_unsigned(10033, LUT_AMPL_WIDTH - 1),
		3247 => to_unsigned(10036, LUT_AMPL_WIDTH - 1),
		3248 => to_unsigned(10039, LUT_AMPL_WIDTH - 1),
		3249 => to_unsigned(10042, LUT_AMPL_WIDTH - 1),
		3250 => to_unsigned(10045, LUT_AMPL_WIDTH - 1),
		3251 => to_unsigned(10048, LUT_AMPL_WIDTH - 1),
		3252 => to_unsigned(10051, LUT_AMPL_WIDTH - 1),
		3253 => to_unsigned(10054, LUT_AMPL_WIDTH - 1),
		3254 => to_unsigned(10057, LUT_AMPL_WIDTH - 1),
		3255 => to_unsigned(10060, LUT_AMPL_WIDTH - 1),
		3256 => to_unsigned(10063, LUT_AMPL_WIDTH - 1),
		3257 => to_unsigned(10066, LUT_AMPL_WIDTH - 1),
		3258 => to_unsigned(10069, LUT_AMPL_WIDTH - 1),
		3259 => to_unsigned(10072, LUT_AMPL_WIDTH - 1),
		3260 => to_unsigned(10075, LUT_AMPL_WIDTH - 1),
		3261 => to_unsigned(10078, LUT_AMPL_WIDTH - 1),
		3262 => to_unsigned(10081, LUT_AMPL_WIDTH - 1),
		3263 => to_unsigned(10084, LUT_AMPL_WIDTH - 1),
		3264 => to_unsigned(10087, LUT_AMPL_WIDTH - 1),
		3265 => to_unsigned(10090, LUT_AMPL_WIDTH - 1),
		3266 => to_unsigned(10093, LUT_AMPL_WIDTH - 1),
		3267 => to_unsigned(10096, LUT_AMPL_WIDTH - 1),
		3268 => to_unsigned(10099, LUT_AMPL_WIDTH - 1),
		3269 => to_unsigned(10102, LUT_AMPL_WIDTH - 1),
		3270 => to_unsigned(10105, LUT_AMPL_WIDTH - 1),
		3271 => to_unsigned(10108, LUT_AMPL_WIDTH - 1),
		3272 => to_unsigned(10111, LUT_AMPL_WIDTH - 1),
		3273 => to_unsigned(10114, LUT_AMPL_WIDTH - 1),
		3274 => to_unsigned(10117, LUT_AMPL_WIDTH - 1),
		3275 => to_unsigned(10120, LUT_AMPL_WIDTH - 1),
		3276 => to_unsigned(10123, LUT_AMPL_WIDTH - 1),
		3277 => to_unsigned(10126, LUT_AMPL_WIDTH - 1),
		3278 => to_unsigned(10129, LUT_AMPL_WIDTH - 1),
		3279 => to_unsigned(10132, LUT_AMPL_WIDTH - 1),
		3280 => to_unsigned(10135, LUT_AMPL_WIDTH - 1),
		3281 => to_unsigned(10138, LUT_AMPL_WIDTH - 1),
		3282 => to_unsigned(10141, LUT_AMPL_WIDTH - 1),
		3283 => to_unsigned(10144, LUT_AMPL_WIDTH - 1),
		3284 => to_unsigned(10147, LUT_AMPL_WIDTH - 1),
		3285 => to_unsigned(10150, LUT_AMPL_WIDTH - 1),
		3286 => to_unsigned(10153, LUT_AMPL_WIDTH - 1),
		3287 => to_unsigned(10156, LUT_AMPL_WIDTH - 1),
		3288 => to_unsigned(10159, LUT_AMPL_WIDTH - 1),
		3289 => to_unsigned(10162, LUT_AMPL_WIDTH - 1),
		3290 => to_unsigned(10165, LUT_AMPL_WIDTH - 1),
		3291 => to_unsigned(10168, LUT_AMPL_WIDTH - 1),
		3292 => to_unsigned(10171, LUT_AMPL_WIDTH - 1),
		3293 => to_unsigned(10174, LUT_AMPL_WIDTH - 1),
		3294 => to_unsigned(10177, LUT_AMPL_WIDTH - 1),
		3295 => to_unsigned(10180, LUT_AMPL_WIDTH - 1),
		3296 => to_unsigned(10183, LUT_AMPL_WIDTH - 1),
		3297 => to_unsigned(10186, LUT_AMPL_WIDTH - 1),
		3298 => to_unsigned(10189, LUT_AMPL_WIDTH - 1),
		3299 => to_unsigned(10192, LUT_AMPL_WIDTH - 1),
		3300 => to_unsigned(10195, LUT_AMPL_WIDTH - 1),
		3301 => to_unsigned(10198, LUT_AMPL_WIDTH - 1),
		3302 => to_unsigned(10201, LUT_AMPL_WIDTH - 1),
		3303 => to_unsigned(10204, LUT_AMPL_WIDTH - 1),
		3304 => to_unsigned(10207, LUT_AMPL_WIDTH - 1),
		3305 => to_unsigned(10210, LUT_AMPL_WIDTH - 1),
		3306 => to_unsigned(10213, LUT_AMPL_WIDTH - 1),
		3307 => to_unsigned(10216, LUT_AMPL_WIDTH - 1),
		3308 => to_unsigned(10219, LUT_AMPL_WIDTH - 1),
		3309 => to_unsigned(10222, LUT_AMPL_WIDTH - 1),
		3310 => to_unsigned(10225, LUT_AMPL_WIDTH - 1),
		3311 => to_unsigned(10228, LUT_AMPL_WIDTH - 1),
		3312 => to_unsigned(10231, LUT_AMPL_WIDTH - 1),
		3313 => to_unsigned(10234, LUT_AMPL_WIDTH - 1),
		3314 => to_unsigned(10237, LUT_AMPL_WIDTH - 1),
		3315 => to_unsigned(10240, LUT_AMPL_WIDTH - 1),
		3316 => to_unsigned(10243, LUT_AMPL_WIDTH - 1),
		3317 => to_unsigned(10246, LUT_AMPL_WIDTH - 1),
		3318 => to_unsigned(10249, LUT_AMPL_WIDTH - 1),
		3319 => to_unsigned(10252, LUT_AMPL_WIDTH - 1),
		3320 => to_unsigned(10255, LUT_AMPL_WIDTH - 1),
		3321 => to_unsigned(10258, LUT_AMPL_WIDTH - 1),
		3322 => to_unsigned(10261, LUT_AMPL_WIDTH - 1),
		3323 => to_unsigned(10263, LUT_AMPL_WIDTH - 1),
		3324 => to_unsigned(10266, LUT_AMPL_WIDTH - 1),
		3325 => to_unsigned(10269, LUT_AMPL_WIDTH - 1),
		3326 => to_unsigned(10272, LUT_AMPL_WIDTH - 1),
		3327 => to_unsigned(10275, LUT_AMPL_WIDTH - 1),
		3328 => to_unsigned(10278, LUT_AMPL_WIDTH - 1),
		3329 => to_unsigned(10281, LUT_AMPL_WIDTH - 1),
		3330 => to_unsigned(10284, LUT_AMPL_WIDTH - 1),
		3331 => to_unsigned(10287, LUT_AMPL_WIDTH - 1),
		3332 => to_unsigned(10290, LUT_AMPL_WIDTH - 1),
		3333 => to_unsigned(10293, LUT_AMPL_WIDTH - 1),
		3334 => to_unsigned(10296, LUT_AMPL_WIDTH - 1),
		3335 => to_unsigned(10299, LUT_AMPL_WIDTH - 1),
		3336 => to_unsigned(10302, LUT_AMPL_WIDTH - 1),
		3337 => to_unsigned(10305, LUT_AMPL_WIDTH - 1),
		3338 => to_unsigned(10308, LUT_AMPL_WIDTH - 1),
		3339 => to_unsigned(10311, LUT_AMPL_WIDTH - 1),
		3340 => to_unsigned(10314, LUT_AMPL_WIDTH - 1),
		3341 => to_unsigned(10317, LUT_AMPL_WIDTH - 1),
		3342 => to_unsigned(10320, LUT_AMPL_WIDTH - 1),
		3343 => to_unsigned(10323, LUT_AMPL_WIDTH - 1),
		3344 => to_unsigned(10326, LUT_AMPL_WIDTH - 1),
		3345 => to_unsigned(10329, LUT_AMPL_WIDTH - 1),
		3346 => to_unsigned(10332, LUT_AMPL_WIDTH - 1),
		3347 => to_unsigned(10335, LUT_AMPL_WIDTH - 1),
		3348 => to_unsigned(10338, LUT_AMPL_WIDTH - 1),
		3349 => to_unsigned(10341, LUT_AMPL_WIDTH - 1),
		3350 => to_unsigned(10344, LUT_AMPL_WIDTH - 1),
		3351 => to_unsigned(10347, LUT_AMPL_WIDTH - 1),
		3352 => to_unsigned(10350, LUT_AMPL_WIDTH - 1),
		3353 => to_unsigned(10353, LUT_AMPL_WIDTH - 1),
		3354 => to_unsigned(10356, LUT_AMPL_WIDTH - 1),
		3355 => to_unsigned(10359, LUT_AMPL_WIDTH - 1),
		3356 => to_unsigned(10362, LUT_AMPL_WIDTH - 1),
		3357 => to_unsigned(10365, LUT_AMPL_WIDTH - 1),
		3358 => to_unsigned(10368, LUT_AMPL_WIDTH - 1),
		3359 => to_unsigned(10371, LUT_AMPL_WIDTH - 1),
		3360 => to_unsigned(10374, LUT_AMPL_WIDTH - 1),
		3361 => to_unsigned(10377, LUT_AMPL_WIDTH - 1),
		3362 => to_unsigned(10380, LUT_AMPL_WIDTH - 1),
		3363 => to_unsigned(10383, LUT_AMPL_WIDTH - 1),
		3364 => to_unsigned(10386, LUT_AMPL_WIDTH - 1),
		3365 => to_unsigned(10389, LUT_AMPL_WIDTH - 1),
		3366 => to_unsigned(10392, LUT_AMPL_WIDTH - 1),
		3367 => to_unsigned(10395, LUT_AMPL_WIDTH - 1),
		3368 => to_unsigned(10398, LUT_AMPL_WIDTH - 1),
		3369 => to_unsigned(10401, LUT_AMPL_WIDTH - 1),
		3370 => to_unsigned(10404, LUT_AMPL_WIDTH - 1),
		3371 => to_unsigned(10407, LUT_AMPL_WIDTH - 1),
		3372 => to_unsigned(10410, LUT_AMPL_WIDTH - 1),
		3373 => to_unsigned(10413, LUT_AMPL_WIDTH - 1),
		3374 => to_unsigned(10416, LUT_AMPL_WIDTH - 1),
		3375 => to_unsigned(10419, LUT_AMPL_WIDTH - 1),
		3376 => to_unsigned(10421, LUT_AMPL_WIDTH - 1),
		3377 => to_unsigned(10424, LUT_AMPL_WIDTH - 1),
		3378 => to_unsigned(10427, LUT_AMPL_WIDTH - 1),
		3379 => to_unsigned(10430, LUT_AMPL_WIDTH - 1),
		3380 => to_unsigned(10433, LUT_AMPL_WIDTH - 1),
		3381 => to_unsigned(10436, LUT_AMPL_WIDTH - 1),
		3382 => to_unsigned(10439, LUT_AMPL_WIDTH - 1),
		3383 => to_unsigned(10442, LUT_AMPL_WIDTH - 1),
		3384 => to_unsigned(10445, LUT_AMPL_WIDTH - 1),
		3385 => to_unsigned(10448, LUT_AMPL_WIDTH - 1),
		3386 => to_unsigned(10451, LUT_AMPL_WIDTH - 1),
		3387 => to_unsigned(10454, LUT_AMPL_WIDTH - 1),
		3388 => to_unsigned(10457, LUT_AMPL_WIDTH - 1),
		3389 => to_unsigned(10460, LUT_AMPL_WIDTH - 1),
		3390 => to_unsigned(10463, LUT_AMPL_WIDTH - 1),
		3391 => to_unsigned(10466, LUT_AMPL_WIDTH - 1),
		3392 => to_unsigned(10469, LUT_AMPL_WIDTH - 1),
		3393 => to_unsigned(10472, LUT_AMPL_WIDTH - 1),
		3394 => to_unsigned(10475, LUT_AMPL_WIDTH - 1),
		3395 => to_unsigned(10478, LUT_AMPL_WIDTH - 1),
		3396 => to_unsigned(10481, LUT_AMPL_WIDTH - 1),
		3397 => to_unsigned(10484, LUT_AMPL_WIDTH - 1),
		3398 => to_unsigned(10487, LUT_AMPL_WIDTH - 1),
		3399 => to_unsigned(10490, LUT_AMPL_WIDTH - 1),
		3400 => to_unsigned(10493, LUT_AMPL_WIDTH - 1),
		3401 => to_unsigned(10496, LUT_AMPL_WIDTH - 1),
		3402 => to_unsigned(10499, LUT_AMPL_WIDTH - 1),
		3403 => to_unsigned(10502, LUT_AMPL_WIDTH - 1),
		3404 => to_unsigned(10505, LUT_AMPL_WIDTH - 1),
		3405 => to_unsigned(10508, LUT_AMPL_WIDTH - 1),
		3406 => to_unsigned(10511, LUT_AMPL_WIDTH - 1),
		3407 => to_unsigned(10514, LUT_AMPL_WIDTH - 1),
		3408 => to_unsigned(10517, LUT_AMPL_WIDTH - 1),
		3409 => to_unsigned(10520, LUT_AMPL_WIDTH - 1),
		3410 => to_unsigned(10523, LUT_AMPL_WIDTH - 1),
		3411 => to_unsigned(10526, LUT_AMPL_WIDTH - 1),
		3412 => to_unsigned(10529, LUT_AMPL_WIDTH - 1),
		3413 => to_unsigned(10532, LUT_AMPL_WIDTH - 1),
		3414 => to_unsigned(10535, LUT_AMPL_WIDTH - 1),
		3415 => to_unsigned(10538, LUT_AMPL_WIDTH - 1),
		3416 => to_unsigned(10541, LUT_AMPL_WIDTH - 1),
		3417 => to_unsigned(10544, LUT_AMPL_WIDTH - 1),
		3418 => to_unsigned(10546, LUT_AMPL_WIDTH - 1),
		3419 => to_unsigned(10549, LUT_AMPL_WIDTH - 1),
		3420 => to_unsigned(10552, LUT_AMPL_WIDTH - 1),
		3421 => to_unsigned(10555, LUT_AMPL_WIDTH - 1),
		3422 => to_unsigned(10558, LUT_AMPL_WIDTH - 1),
		3423 => to_unsigned(10561, LUT_AMPL_WIDTH - 1),
		3424 => to_unsigned(10564, LUT_AMPL_WIDTH - 1),
		3425 => to_unsigned(10567, LUT_AMPL_WIDTH - 1),
		3426 => to_unsigned(10570, LUT_AMPL_WIDTH - 1),
		3427 => to_unsigned(10573, LUT_AMPL_WIDTH - 1),
		3428 => to_unsigned(10576, LUT_AMPL_WIDTH - 1),
		3429 => to_unsigned(10579, LUT_AMPL_WIDTH - 1),
		3430 => to_unsigned(10582, LUT_AMPL_WIDTH - 1),
		3431 => to_unsigned(10585, LUT_AMPL_WIDTH - 1),
		3432 => to_unsigned(10588, LUT_AMPL_WIDTH - 1),
		3433 => to_unsigned(10591, LUT_AMPL_WIDTH - 1),
		3434 => to_unsigned(10594, LUT_AMPL_WIDTH - 1),
		3435 => to_unsigned(10597, LUT_AMPL_WIDTH - 1),
		3436 => to_unsigned(10600, LUT_AMPL_WIDTH - 1),
		3437 => to_unsigned(10603, LUT_AMPL_WIDTH - 1),
		3438 => to_unsigned(10606, LUT_AMPL_WIDTH - 1),
		3439 => to_unsigned(10609, LUT_AMPL_WIDTH - 1),
		3440 => to_unsigned(10612, LUT_AMPL_WIDTH - 1),
		3441 => to_unsigned(10615, LUT_AMPL_WIDTH - 1),
		3442 => to_unsigned(10618, LUT_AMPL_WIDTH - 1),
		3443 => to_unsigned(10621, LUT_AMPL_WIDTH - 1),
		3444 => to_unsigned(10624, LUT_AMPL_WIDTH - 1),
		3445 => to_unsigned(10627, LUT_AMPL_WIDTH - 1),
		3446 => to_unsigned(10630, LUT_AMPL_WIDTH - 1),
		3447 => to_unsigned(10633, LUT_AMPL_WIDTH - 1),
		3448 => to_unsigned(10636, LUT_AMPL_WIDTH - 1),
		3449 => to_unsigned(10639, LUT_AMPL_WIDTH - 1),
		3450 => to_unsigned(10642, LUT_AMPL_WIDTH - 1),
		3451 => to_unsigned(10645, LUT_AMPL_WIDTH - 1),
		3452 => to_unsigned(10648, LUT_AMPL_WIDTH - 1),
		3453 => to_unsigned(10651, LUT_AMPL_WIDTH - 1),
		3454 => to_unsigned(10654, LUT_AMPL_WIDTH - 1),
		3455 => to_unsigned(10656, LUT_AMPL_WIDTH - 1),
		3456 => to_unsigned(10659, LUT_AMPL_WIDTH - 1),
		3457 => to_unsigned(10662, LUT_AMPL_WIDTH - 1),
		3458 => to_unsigned(10665, LUT_AMPL_WIDTH - 1),
		3459 => to_unsigned(10668, LUT_AMPL_WIDTH - 1),
		3460 => to_unsigned(10671, LUT_AMPL_WIDTH - 1),
		3461 => to_unsigned(10674, LUT_AMPL_WIDTH - 1),
		3462 => to_unsigned(10677, LUT_AMPL_WIDTH - 1),
		3463 => to_unsigned(10680, LUT_AMPL_WIDTH - 1),
		3464 => to_unsigned(10683, LUT_AMPL_WIDTH - 1),
		3465 => to_unsigned(10686, LUT_AMPL_WIDTH - 1),
		3466 => to_unsigned(10689, LUT_AMPL_WIDTH - 1),
		3467 => to_unsigned(10692, LUT_AMPL_WIDTH - 1),
		3468 => to_unsigned(10695, LUT_AMPL_WIDTH - 1),
		3469 => to_unsigned(10698, LUT_AMPL_WIDTH - 1),
		3470 => to_unsigned(10701, LUT_AMPL_WIDTH - 1),
		3471 => to_unsigned(10704, LUT_AMPL_WIDTH - 1),
		3472 => to_unsigned(10707, LUT_AMPL_WIDTH - 1),
		3473 => to_unsigned(10710, LUT_AMPL_WIDTH - 1),
		3474 => to_unsigned(10713, LUT_AMPL_WIDTH - 1),
		3475 => to_unsigned(10716, LUT_AMPL_WIDTH - 1),
		3476 => to_unsigned(10719, LUT_AMPL_WIDTH - 1),
		3477 => to_unsigned(10722, LUT_AMPL_WIDTH - 1),
		3478 => to_unsigned(10725, LUT_AMPL_WIDTH - 1),
		3479 => to_unsigned(10728, LUT_AMPL_WIDTH - 1),
		3480 => to_unsigned(10731, LUT_AMPL_WIDTH - 1),
		3481 => to_unsigned(10734, LUT_AMPL_WIDTH - 1),
		3482 => to_unsigned(10737, LUT_AMPL_WIDTH - 1),
		3483 => to_unsigned(10740, LUT_AMPL_WIDTH - 1),
		3484 => to_unsigned(10743, LUT_AMPL_WIDTH - 1),
		3485 => to_unsigned(10746, LUT_AMPL_WIDTH - 1),
		3486 => to_unsigned(10749, LUT_AMPL_WIDTH - 1),
		3487 => to_unsigned(10751, LUT_AMPL_WIDTH - 1),
		3488 => to_unsigned(10754, LUT_AMPL_WIDTH - 1),
		3489 => to_unsigned(10757, LUT_AMPL_WIDTH - 1),
		3490 => to_unsigned(10760, LUT_AMPL_WIDTH - 1),
		3491 => to_unsigned(10763, LUT_AMPL_WIDTH - 1),
		3492 => to_unsigned(10766, LUT_AMPL_WIDTH - 1),
		3493 => to_unsigned(10769, LUT_AMPL_WIDTH - 1),
		3494 => to_unsigned(10772, LUT_AMPL_WIDTH - 1),
		3495 => to_unsigned(10775, LUT_AMPL_WIDTH - 1),
		3496 => to_unsigned(10778, LUT_AMPL_WIDTH - 1),
		3497 => to_unsigned(10781, LUT_AMPL_WIDTH - 1),
		3498 => to_unsigned(10784, LUT_AMPL_WIDTH - 1),
		3499 => to_unsigned(10787, LUT_AMPL_WIDTH - 1),
		3500 => to_unsigned(10790, LUT_AMPL_WIDTH - 1),
		3501 => to_unsigned(10793, LUT_AMPL_WIDTH - 1),
		3502 => to_unsigned(10796, LUT_AMPL_WIDTH - 1),
		3503 => to_unsigned(10799, LUT_AMPL_WIDTH - 1),
		3504 => to_unsigned(10802, LUT_AMPL_WIDTH - 1),
		3505 => to_unsigned(10805, LUT_AMPL_WIDTH - 1),
		3506 => to_unsigned(10808, LUT_AMPL_WIDTH - 1),
		3507 => to_unsigned(10811, LUT_AMPL_WIDTH - 1),
		3508 => to_unsigned(10814, LUT_AMPL_WIDTH - 1),
		3509 => to_unsigned(10817, LUT_AMPL_WIDTH - 1),
		3510 => to_unsigned(10820, LUT_AMPL_WIDTH - 1),
		3511 => to_unsigned(10823, LUT_AMPL_WIDTH - 1),
		3512 => to_unsigned(10826, LUT_AMPL_WIDTH - 1),
		3513 => to_unsigned(10829, LUT_AMPL_WIDTH - 1),
		3514 => to_unsigned(10832, LUT_AMPL_WIDTH - 1),
		3515 => to_unsigned(10835, LUT_AMPL_WIDTH - 1),
		3516 => to_unsigned(10838, LUT_AMPL_WIDTH - 1),
		3517 => to_unsigned(10840, LUT_AMPL_WIDTH - 1),
		3518 => to_unsigned(10843, LUT_AMPL_WIDTH - 1),
		3519 => to_unsigned(10846, LUT_AMPL_WIDTH - 1),
		3520 => to_unsigned(10849, LUT_AMPL_WIDTH - 1),
		3521 => to_unsigned(10852, LUT_AMPL_WIDTH - 1),
		3522 => to_unsigned(10855, LUT_AMPL_WIDTH - 1),
		3523 => to_unsigned(10858, LUT_AMPL_WIDTH - 1),
		3524 => to_unsigned(10861, LUT_AMPL_WIDTH - 1),
		3525 => to_unsigned(10864, LUT_AMPL_WIDTH - 1),
		3526 => to_unsigned(10867, LUT_AMPL_WIDTH - 1),
		3527 => to_unsigned(10870, LUT_AMPL_WIDTH - 1),
		3528 => to_unsigned(10873, LUT_AMPL_WIDTH - 1),
		3529 => to_unsigned(10876, LUT_AMPL_WIDTH - 1),
		3530 => to_unsigned(10879, LUT_AMPL_WIDTH - 1),
		3531 => to_unsigned(10882, LUT_AMPL_WIDTH - 1),
		3532 => to_unsigned(10885, LUT_AMPL_WIDTH - 1),
		3533 => to_unsigned(10888, LUT_AMPL_WIDTH - 1),
		3534 => to_unsigned(10891, LUT_AMPL_WIDTH - 1),
		3535 => to_unsigned(10894, LUT_AMPL_WIDTH - 1),
		3536 => to_unsigned(10897, LUT_AMPL_WIDTH - 1),
		3537 => to_unsigned(10900, LUT_AMPL_WIDTH - 1),
		3538 => to_unsigned(10903, LUT_AMPL_WIDTH - 1),
		3539 => to_unsigned(10906, LUT_AMPL_WIDTH - 1),
		3540 => to_unsigned(10909, LUT_AMPL_WIDTH - 1),
		3541 => to_unsigned(10912, LUT_AMPL_WIDTH - 1),
		3542 => to_unsigned(10915, LUT_AMPL_WIDTH - 1),
		3543 => to_unsigned(10918, LUT_AMPL_WIDTH - 1),
		3544 => to_unsigned(10920, LUT_AMPL_WIDTH - 1),
		3545 => to_unsigned(10923, LUT_AMPL_WIDTH - 1),
		3546 => to_unsigned(10926, LUT_AMPL_WIDTH - 1),
		3547 => to_unsigned(10929, LUT_AMPL_WIDTH - 1),
		3548 => to_unsigned(10932, LUT_AMPL_WIDTH - 1),
		3549 => to_unsigned(10935, LUT_AMPL_WIDTH - 1),
		3550 => to_unsigned(10938, LUT_AMPL_WIDTH - 1),
		3551 => to_unsigned(10941, LUT_AMPL_WIDTH - 1),
		3552 => to_unsigned(10944, LUT_AMPL_WIDTH - 1),
		3553 => to_unsigned(10947, LUT_AMPL_WIDTH - 1),
		3554 => to_unsigned(10950, LUT_AMPL_WIDTH - 1),
		3555 => to_unsigned(10953, LUT_AMPL_WIDTH - 1),
		3556 => to_unsigned(10956, LUT_AMPL_WIDTH - 1),
		3557 => to_unsigned(10959, LUT_AMPL_WIDTH - 1),
		3558 => to_unsigned(10962, LUT_AMPL_WIDTH - 1),
		3559 => to_unsigned(10965, LUT_AMPL_WIDTH - 1),
		3560 => to_unsigned(10968, LUT_AMPL_WIDTH - 1),
		3561 => to_unsigned(10971, LUT_AMPL_WIDTH - 1),
		3562 => to_unsigned(10974, LUT_AMPL_WIDTH - 1),
		3563 => to_unsigned(10977, LUT_AMPL_WIDTH - 1),
		3564 => to_unsigned(10980, LUT_AMPL_WIDTH - 1),
		3565 => to_unsigned(10983, LUT_AMPL_WIDTH - 1),
		3566 => to_unsigned(10986, LUT_AMPL_WIDTH - 1),
		3567 => to_unsigned(10989, LUT_AMPL_WIDTH - 1),
		3568 => to_unsigned(10992, LUT_AMPL_WIDTH - 1),
		3569 => to_unsigned(10994, LUT_AMPL_WIDTH - 1),
		3570 => to_unsigned(10997, LUT_AMPL_WIDTH - 1),
		3571 => to_unsigned(11000, LUT_AMPL_WIDTH - 1),
		3572 => to_unsigned(11003, LUT_AMPL_WIDTH - 1),
		3573 => to_unsigned(11006, LUT_AMPL_WIDTH - 1),
		3574 => to_unsigned(11009, LUT_AMPL_WIDTH - 1),
		3575 => to_unsigned(11012, LUT_AMPL_WIDTH - 1),
		3576 => to_unsigned(11015, LUT_AMPL_WIDTH - 1),
		3577 => to_unsigned(11018, LUT_AMPL_WIDTH - 1),
		3578 => to_unsigned(11021, LUT_AMPL_WIDTH - 1),
		3579 => to_unsigned(11024, LUT_AMPL_WIDTH - 1),
		3580 => to_unsigned(11027, LUT_AMPL_WIDTH - 1),
		3581 => to_unsigned(11030, LUT_AMPL_WIDTH - 1),
		3582 => to_unsigned(11033, LUT_AMPL_WIDTH - 1),
		3583 => to_unsigned(11036, LUT_AMPL_WIDTH - 1),
		3584 => to_unsigned(11039, LUT_AMPL_WIDTH - 1),
		3585 => to_unsigned(11042, LUT_AMPL_WIDTH - 1),
		3586 => to_unsigned(11045, LUT_AMPL_WIDTH - 1),
		3587 => to_unsigned(11048, LUT_AMPL_WIDTH - 1),
		3588 => to_unsigned(11051, LUT_AMPL_WIDTH - 1),
		3589 => to_unsigned(11054, LUT_AMPL_WIDTH - 1),
		3590 => to_unsigned(11057, LUT_AMPL_WIDTH - 1),
		3591 => to_unsigned(11060, LUT_AMPL_WIDTH - 1),
		3592 => to_unsigned(11063, LUT_AMPL_WIDTH - 1),
		3593 => to_unsigned(11065, LUT_AMPL_WIDTH - 1),
		3594 => to_unsigned(11068, LUT_AMPL_WIDTH - 1),
		3595 => to_unsigned(11071, LUT_AMPL_WIDTH - 1),
		3596 => to_unsigned(11074, LUT_AMPL_WIDTH - 1),
		3597 => to_unsigned(11077, LUT_AMPL_WIDTH - 1),
		3598 => to_unsigned(11080, LUT_AMPL_WIDTH - 1),
		3599 => to_unsigned(11083, LUT_AMPL_WIDTH - 1),
		3600 => to_unsigned(11086, LUT_AMPL_WIDTH - 1),
		3601 => to_unsigned(11089, LUT_AMPL_WIDTH - 1),
		3602 => to_unsigned(11092, LUT_AMPL_WIDTH - 1),
		3603 => to_unsigned(11095, LUT_AMPL_WIDTH - 1),
		3604 => to_unsigned(11098, LUT_AMPL_WIDTH - 1),
		3605 => to_unsigned(11101, LUT_AMPL_WIDTH - 1),
		3606 => to_unsigned(11104, LUT_AMPL_WIDTH - 1),
		3607 => to_unsigned(11107, LUT_AMPL_WIDTH - 1),
		3608 => to_unsigned(11110, LUT_AMPL_WIDTH - 1),
		3609 => to_unsigned(11113, LUT_AMPL_WIDTH - 1),
		3610 => to_unsigned(11116, LUT_AMPL_WIDTH - 1),
		3611 => to_unsigned(11119, LUT_AMPL_WIDTH - 1),
		3612 => to_unsigned(11122, LUT_AMPL_WIDTH - 1),
		3613 => to_unsigned(11125, LUT_AMPL_WIDTH - 1),
		3614 => to_unsigned(11128, LUT_AMPL_WIDTH - 1),
		3615 => to_unsigned(11131, LUT_AMPL_WIDTH - 1),
		3616 => to_unsigned(11133, LUT_AMPL_WIDTH - 1),
		3617 => to_unsigned(11136, LUT_AMPL_WIDTH - 1),
		3618 => to_unsigned(11139, LUT_AMPL_WIDTH - 1),
		3619 => to_unsigned(11142, LUT_AMPL_WIDTH - 1),
		3620 => to_unsigned(11145, LUT_AMPL_WIDTH - 1),
		3621 => to_unsigned(11148, LUT_AMPL_WIDTH - 1),
		3622 => to_unsigned(11151, LUT_AMPL_WIDTH - 1),
		3623 => to_unsigned(11154, LUT_AMPL_WIDTH - 1),
		3624 => to_unsigned(11157, LUT_AMPL_WIDTH - 1),
		3625 => to_unsigned(11160, LUT_AMPL_WIDTH - 1),
		3626 => to_unsigned(11163, LUT_AMPL_WIDTH - 1),
		3627 => to_unsigned(11166, LUT_AMPL_WIDTH - 1),
		3628 => to_unsigned(11169, LUT_AMPL_WIDTH - 1),
		3629 => to_unsigned(11172, LUT_AMPL_WIDTH - 1),
		3630 => to_unsigned(11175, LUT_AMPL_WIDTH - 1),
		3631 => to_unsigned(11178, LUT_AMPL_WIDTH - 1),
		3632 => to_unsigned(11181, LUT_AMPL_WIDTH - 1),
		3633 => to_unsigned(11184, LUT_AMPL_WIDTH - 1),
		3634 => to_unsigned(11187, LUT_AMPL_WIDTH - 1),
		3635 => to_unsigned(11190, LUT_AMPL_WIDTH - 1),
		3636 => to_unsigned(11193, LUT_AMPL_WIDTH - 1),
		3637 => to_unsigned(11195, LUT_AMPL_WIDTH - 1),
		3638 => to_unsigned(11198, LUT_AMPL_WIDTH - 1),
		3639 => to_unsigned(11201, LUT_AMPL_WIDTH - 1),
		3640 => to_unsigned(11204, LUT_AMPL_WIDTH - 1),
		3641 => to_unsigned(11207, LUT_AMPL_WIDTH - 1),
		3642 => to_unsigned(11210, LUT_AMPL_WIDTH - 1),
		3643 => to_unsigned(11213, LUT_AMPL_WIDTH - 1),
		3644 => to_unsigned(11216, LUT_AMPL_WIDTH - 1),
		3645 => to_unsigned(11219, LUT_AMPL_WIDTH - 1),
		3646 => to_unsigned(11222, LUT_AMPL_WIDTH - 1),
		3647 => to_unsigned(11225, LUT_AMPL_WIDTH - 1),
		3648 => to_unsigned(11228, LUT_AMPL_WIDTH - 1),
		3649 => to_unsigned(11231, LUT_AMPL_WIDTH - 1),
		3650 => to_unsigned(11234, LUT_AMPL_WIDTH - 1),
		3651 => to_unsigned(11237, LUT_AMPL_WIDTH - 1),
		3652 => to_unsigned(11240, LUT_AMPL_WIDTH - 1),
		3653 => to_unsigned(11243, LUT_AMPL_WIDTH - 1),
		3654 => to_unsigned(11246, LUT_AMPL_WIDTH - 1),
		3655 => to_unsigned(11249, LUT_AMPL_WIDTH - 1),
		3656 => to_unsigned(11252, LUT_AMPL_WIDTH - 1),
		3657 => to_unsigned(11255, LUT_AMPL_WIDTH - 1),
		3658 => to_unsigned(11257, LUT_AMPL_WIDTH - 1),
		3659 => to_unsigned(11260, LUT_AMPL_WIDTH - 1),
		3660 => to_unsigned(11263, LUT_AMPL_WIDTH - 1),
		3661 => to_unsigned(11266, LUT_AMPL_WIDTH - 1),
		3662 => to_unsigned(11269, LUT_AMPL_WIDTH - 1),
		3663 => to_unsigned(11272, LUT_AMPL_WIDTH - 1),
		3664 => to_unsigned(11275, LUT_AMPL_WIDTH - 1),
		3665 => to_unsigned(11278, LUT_AMPL_WIDTH - 1),
		3666 => to_unsigned(11281, LUT_AMPL_WIDTH - 1),
		3667 => to_unsigned(11284, LUT_AMPL_WIDTH - 1),
		3668 => to_unsigned(11287, LUT_AMPL_WIDTH - 1),
		3669 => to_unsigned(11290, LUT_AMPL_WIDTH - 1),
		3670 => to_unsigned(11293, LUT_AMPL_WIDTH - 1),
		3671 => to_unsigned(11296, LUT_AMPL_WIDTH - 1),
		3672 => to_unsigned(11299, LUT_AMPL_WIDTH - 1),
		3673 => to_unsigned(11302, LUT_AMPL_WIDTH - 1),
		3674 => to_unsigned(11305, LUT_AMPL_WIDTH - 1),
		3675 => to_unsigned(11308, LUT_AMPL_WIDTH - 1),
		3676 => to_unsigned(11311, LUT_AMPL_WIDTH - 1),
		3677 => to_unsigned(11314, LUT_AMPL_WIDTH - 1),
		3678 => to_unsigned(11316, LUT_AMPL_WIDTH - 1),
		3679 => to_unsigned(11319, LUT_AMPL_WIDTH - 1),
		3680 => to_unsigned(11322, LUT_AMPL_WIDTH - 1),
		3681 => to_unsigned(11325, LUT_AMPL_WIDTH - 1),
		3682 => to_unsigned(11328, LUT_AMPL_WIDTH - 1),
		3683 => to_unsigned(11331, LUT_AMPL_WIDTH - 1),
		3684 => to_unsigned(11334, LUT_AMPL_WIDTH - 1),
		3685 => to_unsigned(11337, LUT_AMPL_WIDTH - 1),
		3686 => to_unsigned(11340, LUT_AMPL_WIDTH - 1),
		3687 => to_unsigned(11343, LUT_AMPL_WIDTH - 1),
		3688 => to_unsigned(11346, LUT_AMPL_WIDTH - 1),
		3689 => to_unsigned(11349, LUT_AMPL_WIDTH - 1),
		3690 => to_unsigned(11352, LUT_AMPL_WIDTH - 1),
		3691 => to_unsigned(11355, LUT_AMPL_WIDTH - 1),
		3692 => to_unsigned(11358, LUT_AMPL_WIDTH - 1),
		3693 => to_unsigned(11361, LUT_AMPL_WIDTH - 1),
		3694 => to_unsigned(11364, LUT_AMPL_WIDTH - 1),
		3695 => to_unsigned(11367, LUT_AMPL_WIDTH - 1),
		3696 => to_unsigned(11370, LUT_AMPL_WIDTH - 1),
		3697 => to_unsigned(11372, LUT_AMPL_WIDTH - 1),
		3698 => to_unsigned(11375, LUT_AMPL_WIDTH - 1),
		3699 => to_unsigned(11378, LUT_AMPL_WIDTH - 1),
		3700 => to_unsigned(11381, LUT_AMPL_WIDTH - 1),
		3701 => to_unsigned(11384, LUT_AMPL_WIDTH - 1),
		3702 => to_unsigned(11387, LUT_AMPL_WIDTH - 1),
		3703 => to_unsigned(11390, LUT_AMPL_WIDTH - 1),
		3704 => to_unsigned(11393, LUT_AMPL_WIDTH - 1),
		3705 => to_unsigned(11396, LUT_AMPL_WIDTH - 1),
		3706 => to_unsigned(11399, LUT_AMPL_WIDTH - 1),
		3707 => to_unsigned(11402, LUT_AMPL_WIDTH - 1),
		3708 => to_unsigned(11405, LUT_AMPL_WIDTH - 1),
		3709 => to_unsigned(11408, LUT_AMPL_WIDTH - 1),
		3710 => to_unsigned(11411, LUT_AMPL_WIDTH - 1),
		3711 => to_unsigned(11414, LUT_AMPL_WIDTH - 1),
		3712 => to_unsigned(11417, LUT_AMPL_WIDTH - 1),
		3713 => to_unsigned(11420, LUT_AMPL_WIDTH - 1),
		3714 => to_unsigned(11423, LUT_AMPL_WIDTH - 1),
		3715 => to_unsigned(11425, LUT_AMPL_WIDTH - 1),
		3716 => to_unsigned(11428, LUT_AMPL_WIDTH - 1),
		3717 => to_unsigned(11431, LUT_AMPL_WIDTH - 1),
		3718 => to_unsigned(11434, LUT_AMPL_WIDTH - 1),
		3719 => to_unsigned(11437, LUT_AMPL_WIDTH - 1),
		3720 => to_unsigned(11440, LUT_AMPL_WIDTH - 1),
		3721 => to_unsigned(11443, LUT_AMPL_WIDTH - 1),
		3722 => to_unsigned(11446, LUT_AMPL_WIDTH - 1),
		3723 => to_unsigned(11449, LUT_AMPL_WIDTH - 1),
		3724 => to_unsigned(11452, LUT_AMPL_WIDTH - 1),
		3725 => to_unsigned(11455, LUT_AMPL_WIDTH - 1),
		3726 => to_unsigned(11458, LUT_AMPL_WIDTH - 1),
		3727 => to_unsigned(11461, LUT_AMPL_WIDTH - 1),
		3728 => to_unsigned(11464, LUT_AMPL_WIDTH - 1),
		3729 => to_unsigned(11467, LUT_AMPL_WIDTH - 1),
		3730 => to_unsigned(11470, LUT_AMPL_WIDTH - 1),
		3731 => to_unsigned(11473, LUT_AMPL_WIDTH - 1),
		3732 => to_unsigned(11476, LUT_AMPL_WIDTH - 1),
		3733 => to_unsigned(11478, LUT_AMPL_WIDTH - 1),
		3734 => to_unsigned(11481, LUT_AMPL_WIDTH - 1),
		3735 => to_unsigned(11484, LUT_AMPL_WIDTH - 1),
		3736 => to_unsigned(11487, LUT_AMPL_WIDTH - 1),
		3737 => to_unsigned(11490, LUT_AMPL_WIDTH - 1),
		3738 => to_unsigned(11493, LUT_AMPL_WIDTH - 1),
		3739 => to_unsigned(11496, LUT_AMPL_WIDTH - 1),
		3740 => to_unsigned(11499, LUT_AMPL_WIDTH - 1),
		3741 => to_unsigned(11502, LUT_AMPL_WIDTH - 1),
		3742 => to_unsigned(11505, LUT_AMPL_WIDTH - 1),
		3743 => to_unsigned(11508, LUT_AMPL_WIDTH - 1),
		3744 => to_unsigned(11511, LUT_AMPL_WIDTH - 1),
		3745 => to_unsigned(11514, LUT_AMPL_WIDTH - 1),
		3746 => to_unsigned(11517, LUT_AMPL_WIDTH - 1),
		3747 => to_unsigned(11520, LUT_AMPL_WIDTH - 1),
		3748 => to_unsigned(11523, LUT_AMPL_WIDTH - 1),
		3749 => to_unsigned(11526, LUT_AMPL_WIDTH - 1),
		3750 => to_unsigned(11528, LUT_AMPL_WIDTH - 1),
		3751 => to_unsigned(11531, LUT_AMPL_WIDTH - 1),
		3752 => to_unsigned(11534, LUT_AMPL_WIDTH - 1),
		3753 => to_unsigned(11537, LUT_AMPL_WIDTH - 1),
		3754 => to_unsigned(11540, LUT_AMPL_WIDTH - 1),
		3755 => to_unsigned(11543, LUT_AMPL_WIDTH - 1),
		3756 => to_unsigned(11546, LUT_AMPL_WIDTH - 1),
		3757 => to_unsigned(11549, LUT_AMPL_WIDTH - 1),
		3758 => to_unsigned(11552, LUT_AMPL_WIDTH - 1),
		3759 => to_unsigned(11555, LUT_AMPL_WIDTH - 1),
		3760 => to_unsigned(11558, LUT_AMPL_WIDTH - 1),
		3761 => to_unsigned(11561, LUT_AMPL_WIDTH - 1),
		3762 => to_unsigned(11564, LUT_AMPL_WIDTH - 1),
		3763 => to_unsigned(11567, LUT_AMPL_WIDTH - 1),
		3764 => to_unsigned(11570, LUT_AMPL_WIDTH - 1),
		3765 => to_unsigned(11573, LUT_AMPL_WIDTH - 1),
		3766 => to_unsigned(11575, LUT_AMPL_WIDTH - 1),
		3767 => to_unsigned(11578, LUT_AMPL_WIDTH - 1),
		3768 => to_unsigned(11581, LUT_AMPL_WIDTH - 1),
		3769 => to_unsigned(11584, LUT_AMPL_WIDTH - 1),
		3770 => to_unsigned(11587, LUT_AMPL_WIDTH - 1),
		3771 => to_unsigned(11590, LUT_AMPL_WIDTH - 1),
		3772 => to_unsigned(11593, LUT_AMPL_WIDTH - 1),
		3773 => to_unsigned(11596, LUT_AMPL_WIDTH - 1),
		3774 => to_unsigned(11599, LUT_AMPL_WIDTH - 1),
		3775 => to_unsigned(11602, LUT_AMPL_WIDTH - 1),
		3776 => to_unsigned(11605, LUT_AMPL_WIDTH - 1),
		3777 => to_unsigned(11608, LUT_AMPL_WIDTH - 1),
		3778 => to_unsigned(11611, LUT_AMPL_WIDTH - 1),
		3779 => to_unsigned(11614, LUT_AMPL_WIDTH - 1),
		3780 => to_unsigned(11617, LUT_AMPL_WIDTH - 1),
		3781 => to_unsigned(11620, LUT_AMPL_WIDTH - 1),
		3782 => to_unsigned(11623, LUT_AMPL_WIDTH - 1),
		3783 => to_unsigned(11625, LUT_AMPL_WIDTH - 1),
		3784 => to_unsigned(11628, LUT_AMPL_WIDTH - 1),
		3785 => to_unsigned(11631, LUT_AMPL_WIDTH - 1),
		3786 => to_unsigned(11634, LUT_AMPL_WIDTH - 1),
		3787 => to_unsigned(11637, LUT_AMPL_WIDTH - 1),
		3788 => to_unsigned(11640, LUT_AMPL_WIDTH - 1),
		3789 => to_unsigned(11643, LUT_AMPL_WIDTH - 1),
		3790 => to_unsigned(11646, LUT_AMPL_WIDTH - 1),
		3791 => to_unsigned(11649, LUT_AMPL_WIDTH - 1),
		3792 => to_unsigned(11652, LUT_AMPL_WIDTH - 1),
		3793 => to_unsigned(11655, LUT_AMPL_WIDTH - 1),
		3794 => to_unsigned(11658, LUT_AMPL_WIDTH - 1),
		3795 => to_unsigned(11661, LUT_AMPL_WIDTH - 1),
		3796 => to_unsigned(11664, LUT_AMPL_WIDTH - 1),
		3797 => to_unsigned(11667, LUT_AMPL_WIDTH - 1),
		3798 => to_unsigned(11669, LUT_AMPL_WIDTH - 1),
		3799 => to_unsigned(11672, LUT_AMPL_WIDTH - 1),
		3800 => to_unsigned(11675, LUT_AMPL_WIDTH - 1),
		3801 => to_unsigned(11678, LUT_AMPL_WIDTH - 1),
		3802 => to_unsigned(11681, LUT_AMPL_WIDTH - 1),
		3803 => to_unsigned(11684, LUT_AMPL_WIDTH - 1),
		3804 => to_unsigned(11687, LUT_AMPL_WIDTH - 1),
		3805 => to_unsigned(11690, LUT_AMPL_WIDTH - 1),
		3806 => to_unsigned(11693, LUT_AMPL_WIDTH - 1),
		3807 => to_unsigned(11696, LUT_AMPL_WIDTH - 1),
		3808 => to_unsigned(11699, LUT_AMPL_WIDTH - 1),
		3809 => to_unsigned(11702, LUT_AMPL_WIDTH - 1),
		3810 => to_unsigned(11705, LUT_AMPL_WIDTH - 1),
		3811 => to_unsigned(11708, LUT_AMPL_WIDTH - 1),
		3812 => to_unsigned(11711, LUT_AMPL_WIDTH - 1),
		3813 => to_unsigned(11714, LUT_AMPL_WIDTH - 1),
		3814 => to_unsigned(11716, LUT_AMPL_WIDTH - 1),
		3815 => to_unsigned(11719, LUT_AMPL_WIDTH - 1),
		3816 => to_unsigned(11722, LUT_AMPL_WIDTH - 1),
		3817 => to_unsigned(11725, LUT_AMPL_WIDTH - 1),
		3818 => to_unsigned(11728, LUT_AMPL_WIDTH - 1),
		3819 => to_unsigned(11731, LUT_AMPL_WIDTH - 1),
		3820 => to_unsigned(11734, LUT_AMPL_WIDTH - 1),
		3821 => to_unsigned(11737, LUT_AMPL_WIDTH - 1),
		3822 => to_unsigned(11740, LUT_AMPL_WIDTH - 1),
		3823 => to_unsigned(11743, LUT_AMPL_WIDTH - 1),
		3824 => to_unsigned(11746, LUT_AMPL_WIDTH - 1),
		3825 => to_unsigned(11749, LUT_AMPL_WIDTH - 1),
		3826 => to_unsigned(11752, LUT_AMPL_WIDTH - 1),
		3827 => to_unsigned(11755, LUT_AMPL_WIDTH - 1),
		3828 => to_unsigned(11758, LUT_AMPL_WIDTH - 1),
		3829 => to_unsigned(11760, LUT_AMPL_WIDTH - 1),
		3830 => to_unsigned(11763, LUT_AMPL_WIDTH - 1),
		3831 => to_unsigned(11766, LUT_AMPL_WIDTH - 1),
		3832 => to_unsigned(11769, LUT_AMPL_WIDTH - 1),
		3833 => to_unsigned(11772, LUT_AMPL_WIDTH - 1),
		3834 => to_unsigned(11775, LUT_AMPL_WIDTH - 1),
		3835 => to_unsigned(11778, LUT_AMPL_WIDTH - 1),
		3836 => to_unsigned(11781, LUT_AMPL_WIDTH - 1),
		3837 => to_unsigned(11784, LUT_AMPL_WIDTH - 1),
		3838 => to_unsigned(11787, LUT_AMPL_WIDTH - 1),
		3839 => to_unsigned(11790, LUT_AMPL_WIDTH - 1),
		3840 => to_unsigned(11793, LUT_AMPL_WIDTH - 1),
		3841 => to_unsigned(11796, LUT_AMPL_WIDTH - 1),
		3842 => to_unsigned(11799, LUT_AMPL_WIDTH - 1),
		3843 => to_unsigned(11801, LUT_AMPL_WIDTH - 1),
		3844 => to_unsigned(11804, LUT_AMPL_WIDTH - 1),
		3845 => to_unsigned(11807, LUT_AMPL_WIDTH - 1),
		3846 => to_unsigned(11810, LUT_AMPL_WIDTH - 1),
		3847 => to_unsigned(11813, LUT_AMPL_WIDTH - 1),
		3848 => to_unsigned(11816, LUT_AMPL_WIDTH - 1),
		3849 => to_unsigned(11819, LUT_AMPL_WIDTH - 1),
		3850 => to_unsigned(11822, LUT_AMPL_WIDTH - 1),
		3851 => to_unsigned(11825, LUT_AMPL_WIDTH - 1),
		3852 => to_unsigned(11828, LUT_AMPL_WIDTH - 1),
		3853 => to_unsigned(11831, LUT_AMPL_WIDTH - 1),
		3854 => to_unsigned(11834, LUT_AMPL_WIDTH - 1),
		3855 => to_unsigned(11837, LUT_AMPL_WIDTH - 1),
		3856 => to_unsigned(11840, LUT_AMPL_WIDTH - 1),
		3857 => to_unsigned(11842, LUT_AMPL_WIDTH - 1),
		3858 => to_unsigned(11845, LUT_AMPL_WIDTH - 1),
		3859 => to_unsigned(11848, LUT_AMPL_WIDTH - 1),
		3860 => to_unsigned(11851, LUT_AMPL_WIDTH - 1),
		3861 => to_unsigned(11854, LUT_AMPL_WIDTH - 1),
		3862 => to_unsigned(11857, LUT_AMPL_WIDTH - 1),
		3863 => to_unsigned(11860, LUT_AMPL_WIDTH - 1),
		3864 => to_unsigned(11863, LUT_AMPL_WIDTH - 1),
		3865 => to_unsigned(11866, LUT_AMPL_WIDTH - 1),
		3866 => to_unsigned(11869, LUT_AMPL_WIDTH - 1),
		3867 => to_unsigned(11872, LUT_AMPL_WIDTH - 1),
		3868 => to_unsigned(11875, LUT_AMPL_WIDTH - 1),
		3869 => to_unsigned(11878, LUT_AMPL_WIDTH - 1),
		3870 => to_unsigned(11881, LUT_AMPL_WIDTH - 1),
		3871 => to_unsigned(11883, LUT_AMPL_WIDTH - 1),
		3872 => to_unsigned(11886, LUT_AMPL_WIDTH - 1),
		3873 => to_unsigned(11889, LUT_AMPL_WIDTH - 1),
		3874 => to_unsigned(11892, LUT_AMPL_WIDTH - 1),
		3875 => to_unsigned(11895, LUT_AMPL_WIDTH - 1),
		3876 => to_unsigned(11898, LUT_AMPL_WIDTH - 1),
		3877 => to_unsigned(11901, LUT_AMPL_WIDTH - 1),
		3878 => to_unsigned(11904, LUT_AMPL_WIDTH - 1),
		3879 => to_unsigned(11907, LUT_AMPL_WIDTH - 1),
		3880 => to_unsigned(11910, LUT_AMPL_WIDTH - 1),
		3881 => to_unsigned(11913, LUT_AMPL_WIDTH - 1),
		3882 => to_unsigned(11916, LUT_AMPL_WIDTH - 1),
		3883 => to_unsigned(11919, LUT_AMPL_WIDTH - 1),
		3884 => to_unsigned(11922, LUT_AMPL_WIDTH - 1),
		3885 => to_unsigned(11924, LUT_AMPL_WIDTH - 1),
		3886 => to_unsigned(11927, LUT_AMPL_WIDTH - 1),
		3887 => to_unsigned(11930, LUT_AMPL_WIDTH - 1),
		3888 => to_unsigned(11933, LUT_AMPL_WIDTH - 1),
		3889 => to_unsigned(11936, LUT_AMPL_WIDTH - 1),
		3890 => to_unsigned(11939, LUT_AMPL_WIDTH - 1),
		3891 => to_unsigned(11942, LUT_AMPL_WIDTH - 1),
		3892 => to_unsigned(11945, LUT_AMPL_WIDTH - 1),
		3893 => to_unsigned(11948, LUT_AMPL_WIDTH - 1),
		3894 => to_unsigned(11951, LUT_AMPL_WIDTH - 1),
		3895 => to_unsigned(11954, LUT_AMPL_WIDTH - 1),
		3896 => to_unsigned(11957, LUT_AMPL_WIDTH - 1),
		3897 => to_unsigned(11960, LUT_AMPL_WIDTH - 1),
		3898 => to_unsigned(11962, LUT_AMPL_WIDTH - 1),
		3899 => to_unsigned(11965, LUT_AMPL_WIDTH - 1),
		3900 => to_unsigned(11968, LUT_AMPL_WIDTH - 1),
		3901 => to_unsigned(11971, LUT_AMPL_WIDTH - 1),
		3902 => to_unsigned(11974, LUT_AMPL_WIDTH - 1),
		3903 => to_unsigned(11977, LUT_AMPL_WIDTH - 1),
		3904 => to_unsigned(11980, LUT_AMPL_WIDTH - 1),
		3905 => to_unsigned(11983, LUT_AMPL_WIDTH - 1),
		3906 => to_unsigned(11986, LUT_AMPL_WIDTH - 1),
		3907 => to_unsigned(11989, LUT_AMPL_WIDTH - 1),
		3908 => to_unsigned(11992, LUT_AMPL_WIDTH - 1),
		3909 => to_unsigned(11995, LUT_AMPL_WIDTH - 1),
		3910 => to_unsigned(11998, LUT_AMPL_WIDTH - 1),
		3911 => to_unsigned(12001, LUT_AMPL_WIDTH - 1),
		3912 => to_unsigned(12003, LUT_AMPL_WIDTH - 1),
		3913 => to_unsigned(12006, LUT_AMPL_WIDTH - 1),
		3914 => to_unsigned(12009, LUT_AMPL_WIDTH - 1),
		3915 => to_unsigned(12012, LUT_AMPL_WIDTH - 1),
		3916 => to_unsigned(12015, LUT_AMPL_WIDTH - 1),
		3917 => to_unsigned(12018, LUT_AMPL_WIDTH - 1),
		3918 => to_unsigned(12021, LUT_AMPL_WIDTH - 1),
		3919 => to_unsigned(12024, LUT_AMPL_WIDTH - 1),
		3920 => to_unsigned(12027, LUT_AMPL_WIDTH - 1),
		3921 => to_unsigned(12030, LUT_AMPL_WIDTH - 1),
		3922 => to_unsigned(12033, LUT_AMPL_WIDTH - 1),
		3923 => to_unsigned(12036, LUT_AMPL_WIDTH - 1),
		3924 => to_unsigned(12038, LUT_AMPL_WIDTH - 1),
		3925 => to_unsigned(12041, LUT_AMPL_WIDTH - 1),
		3926 => to_unsigned(12044, LUT_AMPL_WIDTH - 1),
		3927 => to_unsigned(12047, LUT_AMPL_WIDTH - 1),
		3928 => to_unsigned(12050, LUT_AMPL_WIDTH - 1),
		3929 => to_unsigned(12053, LUT_AMPL_WIDTH - 1),
		3930 => to_unsigned(12056, LUT_AMPL_WIDTH - 1),
		3931 => to_unsigned(12059, LUT_AMPL_WIDTH - 1),
		3932 => to_unsigned(12062, LUT_AMPL_WIDTH - 1),
		3933 => to_unsigned(12065, LUT_AMPL_WIDTH - 1),
		3934 => to_unsigned(12068, LUT_AMPL_WIDTH - 1),
		3935 => to_unsigned(12071, LUT_AMPL_WIDTH - 1),
		3936 => to_unsigned(12074, LUT_AMPL_WIDTH - 1),
		3937 => to_unsigned(12076, LUT_AMPL_WIDTH - 1),
		3938 => to_unsigned(12079, LUT_AMPL_WIDTH - 1),
		3939 => to_unsigned(12082, LUT_AMPL_WIDTH - 1),
		3940 => to_unsigned(12085, LUT_AMPL_WIDTH - 1),
		3941 => to_unsigned(12088, LUT_AMPL_WIDTH - 1),
		3942 => to_unsigned(12091, LUT_AMPL_WIDTH - 1),
		3943 => to_unsigned(12094, LUT_AMPL_WIDTH - 1),
		3944 => to_unsigned(12097, LUT_AMPL_WIDTH - 1),
		3945 => to_unsigned(12100, LUT_AMPL_WIDTH - 1),
		3946 => to_unsigned(12103, LUT_AMPL_WIDTH - 1),
		3947 => to_unsigned(12106, LUT_AMPL_WIDTH - 1),
		3948 => to_unsigned(12109, LUT_AMPL_WIDTH - 1),
		3949 => to_unsigned(12112, LUT_AMPL_WIDTH - 1),
		3950 => to_unsigned(12114, LUT_AMPL_WIDTH - 1),
		3951 => to_unsigned(12117, LUT_AMPL_WIDTH - 1),
		3952 => to_unsigned(12120, LUT_AMPL_WIDTH - 1),
		3953 => to_unsigned(12123, LUT_AMPL_WIDTH - 1),
		3954 => to_unsigned(12126, LUT_AMPL_WIDTH - 1),
		3955 => to_unsigned(12129, LUT_AMPL_WIDTH - 1),
		3956 => to_unsigned(12132, LUT_AMPL_WIDTH - 1),
		3957 => to_unsigned(12135, LUT_AMPL_WIDTH - 1),
		3958 => to_unsigned(12138, LUT_AMPL_WIDTH - 1),
		3959 => to_unsigned(12141, LUT_AMPL_WIDTH - 1),
		3960 => to_unsigned(12144, LUT_AMPL_WIDTH - 1),
		3961 => to_unsigned(12147, LUT_AMPL_WIDTH - 1),
		3962 => to_unsigned(12149, LUT_AMPL_WIDTH - 1),
		3963 => to_unsigned(12152, LUT_AMPL_WIDTH - 1),
		3964 => to_unsigned(12155, LUT_AMPL_WIDTH - 1),
		3965 => to_unsigned(12158, LUT_AMPL_WIDTH - 1),
		3966 => to_unsigned(12161, LUT_AMPL_WIDTH - 1),
		3967 => to_unsigned(12164, LUT_AMPL_WIDTH - 1),
		3968 => to_unsigned(12167, LUT_AMPL_WIDTH - 1),
		3969 => to_unsigned(12170, LUT_AMPL_WIDTH - 1),
		3970 => to_unsigned(12173, LUT_AMPL_WIDTH - 1),
		3971 => to_unsigned(12176, LUT_AMPL_WIDTH - 1),
		3972 => to_unsigned(12179, LUT_AMPL_WIDTH - 1),
		3973 => to_unsigned(12182, LUT_AMPL_WIDTH - 1),
		3974 => to_unsigned(12184, LUT_AMPL_WIDTH - 1),
		3975 => to_unsigned(12187, LUT_AMPL_WIDTH - 1),
		3976 => to_unsigned(12190, LUT_AMPL_WIDTH - 1),
		3977 => to_unsigned(12193, LUT_AMPL_WIDTH - 1),
		3978 => to_unsigned(12196, LUT_AMPL_WIDTH - 1),
		3979 => to_unsigned(12199, LUT_AMPL_WIDTH - 1),
		3980 => to_unsigned(12202, LUT_AMPL_WIDTH - 1),
		3981 => to_unsigned(12205, LUT_AMPL_WIDTH - 1),
		3982 => to_unsigned(12208, LUT_AMPL_WIDTH - 1),
		3983 => to_unsigned(12211, LUT_AMPL_WIDTH - 1),
		3984 => to_unsigned(12214, LUT_AMPL_WIDTH - 1),
		3985 => to_unsigned(12217, LUT_AMPL_WIDTH - 1),
		3986 => to_unsigned(12219, LUT_AMPL_WIDTH - 1),
		3987 => to_unsigned(12222, LUT_AMPL_WIDTH - 1),
		3988 => to_unsigned(12225, LUT_AMPL_WIDTH - 1),
		3989 => to_unsigned(12228, LUT_AMPL_WIDTH - 1),
		3990 => to_unsigned(12231, LUT_AMPL_WIDTH - 1),
		3991 => to_unsigned(12234, LUT_AMPL_WIDTH - 1),
		3992 => to_unsigned(12237, LUT_AMPL_WIDTH - 1),
		3993 => to_unsigned(12240, LUT_AMPL_WIDTH - 1),
		3994 => to_unsigned(12243, LUT_AMPL_WIDTH - 1),
		3995 => to_unsigned(12246, LUT_AMPL_WIDTH - 1),
		3996 => to_unsigned(12249, LUT_AMPL_WIDTH - 1),
		3997 => to_unsigned(12251, LUT_AMPL_WIDTH - 1),
		3998 => to_unsigned(12254, LUT_AMPL_WIDTH - 1),
		3999 => to_unsigned(12257, LUT_AMPL_WIDTH - 1),
		4000 => to_unsigned(12260, LUT_AMPL_WIDTH - 1),
		4001 => to_unsigned(12263, LUT_AMPL_WIDTH - 1),
		4002 => to_unsigned(12266, LUT_AMPL_WIDTH - 1),
		4003 => to_unsigned(12269, LUT_AMPL_WIDTH - 1),
		4004 => to_unsigned(12272, LUT_AMPL_WIDTH - 1),
		4005 => to_unsigned(12275, LUT_AMPL_WIDTH - 1),
		4006 => to_unsigned(12278, LUT_AMPL_WIDTH - 1),
		4007 => to_unsigned(12281, LUT_AMPL_WIDTH - 1),
		4008 => to_unsigned(12284, LUT_AMPL_WIDTH - 1),
		4009 => to_unsigned(12286, LUT_AMPL_WIDTH - 1),
		4010 => to_unsigned(12289, LUT_AMPL_WIDTH - 1),
		4011 => to_unsigned(12292, LUT_AMPL_WIDTH - 1),
		4012 => to_unsigned(12295, LUT_AMPL_WIDTH - 1),
		4013 => to_unsigned(12298, LUT_AMPL_WIDTH - 1),
		4014 => to_unsigned(12301, LUT_AMPL_WIDTH - 1),
		4015 => to_unsigned(12304, LUT_AMPL_WIDTH - 1),
		4016 => to_unsigned(12307, LUT_AMPL_WIDTH - 1),
		4017 => to_unsigned(12310, LUT_AMPL_WIDTH - 1),
		4018 => to_unsigned(12313, LUT_AMPL_WIDTH - 1),
		4019 => to_unsigned(12316, LUT_AMPL_WIDTH - 1),
		4020 => to_unsigned(12318, LUT_AMPL_WIDTH - 1),
		4021 => to_unsigned(12321, LUT_AMPL_WIDTH - 1),
		4022 => to_unsigned(12324, LUT_AMPL_WIDTH - 1),
		4023 => to_unsigned(12327, LUT_AMPL_WIDTH - 1),
		4024 => to_unsigned(12330, LUT_AMPL_WIDTH - 1),
		4025 => to_unsigned(12333, LUT_AMPL_WIDTH - 1),
		4026 => to_unsigned(12336, LUT_AMPL_WIDTH - 1),
		4027 => to_unsigned(12339, LUT_AMPL_WIDTH - 1),
		4028 => to_unsigned(12342, LUT_AMPL_WIDTH - 1),
		4029 => to_unsigned(12345, LUT_AMPL_WIDTH - 1),
		4030 => to_unsigned(12348, LUT_AMPL_WIDTH - 1),
		4031 => to_unsigned(12350, LUT_AMPL_WIDTH - 1),
		4032 => to_unsigned(12353, LUT_AMPL_WIDTH - 1),
		4033 => to_unsigned(12356, LUT_AMPL_WIDTH - 1),
		4034 => to_unsigned(12359, LUT_AMPL_WIDTH - 1),
		4035 => to_unsigned(12362, LUT_AMPL_WIDTH - 1),
		4036 => to_unsigned(12365, LUT_AMPL_WIDTH - 1),
		4037 => to_unsigned(12368, LUT_AMPL_WIDTH - 1),
		4038 => to_unsigned(12371, LUT_AMPL_WIDTH - 1),
		4039 => to_unsigned(12374, LUT_AMPL_WIDTH - 1),
		4040 => to_unsigned(12377, LUT_AMPL_WIDTH - 1),
		4041 => to_unsigned(12380, LUT_AMPL_WIDTH - 1),
		4042 => to_unsigned(12382, LUT_AMPL_WIDTH - 1),
		4043 => to_unsigned(12385, LUT_AMPL_WIDTH - 1),
		4044 => to_unsigned(12388, LUT_AMPL_WIDTH - 1),
		4045 => to_unsigned(12391, LUT_AMPL_WIDTH - 1),
		4046 => to_unsigned(12394, LUT_AMPL_WIDTH - 1),
		4047 => to_unsigned(12397, LUT_AMPL_WIDTH - 1),
		4048 => to_unsigned(12400, LUT_AMPL_WIDTH - 1),
		4049 => to_unsigned(12403, LUT_AMPL_WIDTH - 1),
		4050 => to_unsigned(12406, LUT_AMPL_WIDTH - 1),
		4051 => to_unsigned(12409, LUT_AMPL_WIDTH - 1),
		4052 => to_unsigned(12412, LUT_AMPL_WIDTH - 1),
		4053 => to_unsigned(12414, LUT_AMPL_WIDTH - 1),
		4054 => to_unsigned(12417, LUT_AMPL_WIDTH - 1),
		4055 => to_unsigned(12420, LUT_AMPL_WIDTH - 1),
		4056 => to_unsigned(12423, LUT_AMPL_WIDTH - 1),
		4057 => to_unsigned(12426, LUT_AMPL_WIDTH - 1),
		4058 => to_unsigned(12429, LUT_AMPL_WIDTH - 1),
		4059 => to_unsigned(12432, LUT_AMPL_WIDTH - 1),
		4060 => to_unsigned(12435, LUT_AMPL_WIDTH - 1),
		4061 => to_unsigned(12438, LUT_AMPL_WIDTH - 1),
		4062 => to_unsigned(12441, LUT_AMPL_WIDTH - 1),
		4063 => to_unsigned(12444, LUT_AMPL_WIDTH - 1),
		4064 => to_unsigned(12446, LUT_AMPL_WIDTH - 1),
		4065 => to_unsigned(12449, LUT_AMPL_WIDTH - 1),
		4066 => to_unsigned(12452, LUT_AMPL_WIDTH - 1),
		4067 => to_unsigned(12455, LUT_AMPL_WIDTH - 1),
		4068 => to_unsigned(12458, LUT_AMPL_WIDTH - 1),
		4069 => to_unsigned(12461, LUT_AMPL_WIDTH - 1),
		4070 => to_unsigned(12464, LUT_AMPL_WIDTH - 1),
		4071 => to_unsigned(12467, LUT_AMPL_WIDTH - 1),
		4072 => to_unsigned(12470, LUT_AMPL_WIDTH - 1),
		4073 => to_unsigned(12473, LUT_AMPL_WIDTH - 1),
		4074 => to_unsigned(12476, LUT_AMPL_WIDTH - 1),
		4075 => to_unsigned(12478, LUT_AMPL_WIDTH - 1),
		4076 => to_unsigned(12481, LUT_AMPL_WIDTH - 1),
		4077 => to_unsigned(12484, LUT_AMPL_WIDTH - 1),
		4078 => to_unsigned(12487, LUT_AMPL_WIDTH - 1),
		4079 => to_unsigned(12490, LUT_AMPL_WIDTH - 1),
		4080 => to_unsigned(12493, LUT_AMPL_WIDTH - 1),
		4081 => to_unsigned(12496, LUT_AMPL_WIDTH - 1),
		4082 => to_unsigned(12499, LUT_AMPL_WIDTH - 1),
		4083 => to_unsigned(12502, LUT_AMPL_WIDTH - 1),
		4084 => to_unsigned(12505, LUT_AMPL_WIDTH - 1),
		4085 => to_unsigned(12507, LUT_AMPL_WIDTH - 1),
		4086 => to_unsigned(12510, LUT_AMPL_WIDTH - 1),
		4087 => to_unsigned(12513, LUT_AMPL_WIDTH - 1),
		4088 => to_unsigned(12516, LUT_AMPL_WIDTH - 1),
		4089 => to_unsigned(12519, LUT_AMPL_WIDTH - 1),
		4090 => to_unsigned(12522, LUT_AMPL_WIDTH - 1),
		4091 => to_unsigned(12525, LUT_AMPL_WIDTH - 1),
		4092 => to_unsigned(12528, LUT_AMPL_WIDTH - 1),
		4093 => to_unsigned(12531, LUT_AMPL_WIDTH - 1),
		4094 => to_unsigned(12534, LUT_AMPL_WIDTH - 1),
		4095 => to_unsigned(12536, LUT_AMPL_WIDTH - 1),
		4096 => to_unsigned(12539, LUT_AMPL_WIDTH - 1),
		4097 => to_unsigned(12542, LUT_AMPL_WIDTH - 1),
		4098 => to_unsigned(12545, LUT_AMPL_WIDTH - 1),
		4099 => to_unsigned(12548, LUT_AMPL_WIDTH - 1),
		4100 => to_unsigned(12551, LUT_AMPL_WIDTH - 1),
		4101 => to_unsigned(12554, LUT_AMPL_WIDTH - 1),
		4102 => to_unsigned(12557, LUT_AMPL_WIDTH - 1),
		4103 => to_unsigned(12560, LUT_AMPL_WIDTH - 1),
		4104 => to_unsigned(12563, LUT_AMPL_WIDTH - 1),
		4105 => to_unsigned(12566, LUT_AMPL_WIDTH - 1),
		4106 => to_unsigned(12568, LUT_AMPL_WIDTH - 1),
		4107 => to_unsigned(12571, LUT_AMPL_WIDTH - 1),
		4108 => to_unsigned(12574, LUT_AMPL_WIDTH - 1),
		4109 => to_unsigned(12577, LUT_AMPL_WIDTH - 1),
		4110 => to_unsigned(12580, LUT_AMPL_WIDTH - 1),
		4111 => to_unsigned(12583, LUT_AMPL_WIDTH - 1),
		4112 => to_unsigned(12586, LUT_AMPL_WIDTH - 1),
		4113 => to_unsigned(12589, LUT_AMPL_WIDTH - 1),
		4114 => to_unsigned(12592, LUT_AMPL_WIDTH - 1),
		4115 => to_unsigned(12595, LUT_AMPL_WIDTH - 1),
		4116 => to_unsigned(12597, LUT_AMPL_WIDTH - 1),
		4117 => to_unsigned(12600, LUT_AMPL_WIDTH - 1),
		4118 => to_unsigned(12603, LUT_AMPL_WIDTH - 1),
		4119 => to_unsigned(12606, LUT_AMPL_WIDTH - 1),
		4120 => to_unsigned(12609, LUT_AMPL_WIDTH - 1),
		4121 => to_unsigned(12612, LUT_AMPL_WIDTH - 1),
		4122 => to_unsigned(12615, LUT_AMPL_WIDTH - 1),
		4123 => to_unsigned(12618, LUT_AMPL_WIDTH - 1),
		4124 => to_unsigned(12621, LUT_AMPL_WIDTH - 1),
		4125 => to_unsigned(12624, LUT_AMPL_WIDTH - 1),
		4126 => to_unsigned(12626, LUT_AMPL_WIDTH - 1),
		4127 => to_unsigned(12629, LUT_AMPL_WIDTH - 1),
		4128 => to_unsigned(12632, LUT_AMPL_WIDTH - 1),
		4129 => to_unsigned(12635, LUT_AMPL_WIDTH - 1),
		4130 => to_unsigned(12638, LUT_AMPL_WIDTH - 1),
		4131 => to_unsigned(12641, LUT_AMPL_WIDTH - 1),
		4132 => to_unsigned(12644, LUT_AMPL_WIDTH - 1),
		4133 => to_unsigned(12647, LUT_AMPL_WIDTH - 1),
		4134 => to_unsigned(12650, LUT_AMPL_WIDTH - 1),
		4135 => to_unsigned(12652, LUT_AMPL_WIDTH - 1),
		4136 => to_unsigned(12655, LUT_AMPL_WIDTH - 1),
		4137 => to_unsigned(12658, LUT_AMPL_WIDTH - 1),
		4138 => to_unsigned(12661, LUT_AMPL_WIDTH - 1),
		4139 => to_unsigned(12664, LUT_AMPL_WIDTH - 1),
		4140 => to_unsigned(12667, LUT_AMPL_WIDTH - 1),
		4141 => to_unsigned(12670, LUT_AMPL_WIDTH - 1),
		4142 => to_unsigned(12673, LUT_AMPL_WIDTH - 1),
		4143 => to_unsigned(12676, LUT_AMPL_WIDTH - 1),
		4144 => to_unsigned(12679, LUT_AMPL_WIDTH - 1),
		4145 => to_unsigned(12681, LUT_AMPL_WIDTH - 1),
		4146 => to_unsigned(12684, LUT_AMPL_WIDTH - 1),
		4147 => to_unsigned(12687, LUT_AMPL_WIDTH - 1),
		4148 => to_unsigned(12690, LUT_AMPL_WIDTH - 1),
		4149 => to_unsigned(12693, LUT_AMPL_WIDTH - 1),
		4150 => to_unsigned(12696, LUT_AMPL_WIDTH - 1),
		4151 => to_unsigned(12699, LUT_AMPL_WIDTH - 1),
		4152 => to_unsigned(12702, LUT_AMPL_WIDTH - 1),
		4153 => to_unsigned(12705, LUT_AMPL_WIDTH - 1),
		4154 => to_unsigned(12708, LUT_AMPL_WIDTH - 1),
		4155 => to_unsigned(12710, LUT_AMPL_WIDTH - 1),
		4156 => to_unsigned(12713, LUT_AMPL_WIDTH - 1),
		4157 => to_unsigned(12716, LUT_AMPL_WIDTH - 1),
		4158 => to_unsigned(12719, LUT_AMPL_WIDTH - 1),
		4159 => to_unsigned(12722, LUT_AMPL_WIDTH - 1),
		4160 => to_unsigned(12725, LUT_AMPL_WIDTH - 1),
		4161 => to_unsigned(12728, LUT_AMPL_WIDTH - 1),
		4162 => to_unsigned(12731, LUT_AMPL_WIDTH - 1),
		4163 => to_unsigned(12734, LUT_AMPL_WIDTH - 1),
		4164 => to_unsigned(12736, LUT_AMPL_WIDTH - 1),
		4165 => to_unsigned(12739, LUT_AMPL_WIDTH - 1),
		4166 => to_unsigned(12742, LUT_AMPL_WIDTH - 1),
		4167 => to_unsigned(12745, LUT_AMPL_WIDTH - 1),
		4168 => to_unsigned(12748, LUT_AMPL_WIDTH - 1),
		4169 => to_unsigned(12751, LUT_AMPL_WIDTH - 1),
		4170 => to_unsigned(12754, LUT_AMPL_WIDTH - 1),
		4171 => to_unsigned(12757, LUT_AMPL_WIDTH - 1),
		4172 => to_unsigned(12760, LUT_AMPL_WIDTH - 1),
		4173 => to_unsigned(12763, LUT_AMPL_WIDTH - 1),
		4174 => to_unsigned(12765, LUT_AMPL_WIDTH - 1),
		4175 => to_unsigned(12768, LUT_AMPL_WIDTH - 1),
		4176 => to_unsigned(12771, LUT_AMPL_WIDTH - 1),
		4177 => to_unsigned(12774, LUT_AMPL_WIDTH - 1),
		4178 => to_unsigned(12777, LUT_AMPL_WIDTH - 1),
		4179 => to_unsigned(12780, LUT_AMPL_WIDTH - 1),
		4180 => to_unsigned(12783, LUT_AMPL_WIDTH - 1),
		4181 => to_unsigned(12786, LUT_AMPL_WIDTH - 1),
		4182 => to_unsigned(12789, LUT_AMPL_WIDTH - 1),
		4183 => to_unsigned(12791, LUT_AMPL_WIDTH - 1),
		4184 => to_unsigned(12794, LUT_AMPL_WIDTH - 1),
		4185 => to_unsigned(12797, LUT_AMPL_WIDTH - 1),
		4186 => to_unsigned(12800, LUT_AMPL_WIDTH - 1),
		4187 => to_unsigned(12803, LUT_AMPL_WIDTH - 1),
		4188 => to_unsigned(12806, LUT_AMPL_WIDTH - 1),
		4189 => to_unsigned(12809, LUT_AMPL_WIDTH - 1),
		4190 => to_unsigned(12812, LUT_AMPL_WIDTH - 1),
		4191 => to_unsigned(12815, LUT_AMPL_WIDTH - 1),
		4192 => to_unsigned(12817, LUT_AMPL_WIDTH - 1),
		4193 => to_unsigned(12820, LUT_AMPL_WIDTH - 1),
		4194 => to_unsigned(12823, LUT_AMPL_WIDTH - 1),
		4195 => to_unsigned(12826, LUT_AMPL_WIDTH - 1),
		4196 => to_unsigned(12829, LUT_AMPL_WIDTH - 1),
		4197 => to_unsigned(12832, LUT_AMPL_WIDTH - 1),
		4198 => to_unsigned(12835, LUT_AMPL_WIDTH - 1),
		4199 => to_unsigned(12838, LUT_AMPL_WIDTH - 1),
		4200 => to_unsigned(12841, LUT_AMPL_WIDTH - 1),
		4201 => to_unsigned(12843, LUT_AMPL_WIDTH - 1),
		4202 => to_unsigned(12846, LUT_AMPL_WIDTH - 1),
		4203 => to_unsigned(12849, LUT_AMPL_WIDTH - 1),
		4204 => to_unsigned(12852, LUT_AMPL_WIDTH - 1),
		4205 => to_unsigned(12855, LUT_AMPL_WIDTH - 1),
		4206 => to_unsigned(12858, LUT_AMPL_WIDTH - 1),
		4207 => to_unsigned(12861, LUT_AMPL_WIDTH - 1),
		4208 => to_unsigned(12864, LUT_AMPL_WIDTH - 1),
		4209 => to_unsigned(12867, LUT_AMPL_WIDTH - 1),
		4210 => to_unsigned(12870, LUT_AMPL_WIDTH - 1),
		4211 => to_unsigned(12872, LUT_AMPL_WIDTH - 1),
		4212 => to_unsigned(12875, LUT_AMPL_WIDTH - 1),
		4213 => to_unsigned(12878, LUT_AMPL_WIDTH - 1),
		4214 => to_unsigned(12881, LUT_AMPL_WIDTH - 1),
		4215 => to_unsigned(12884, LUT_AMPL_WIDTH - 1),
		4216 => to_unsigned(12887, LUT_AMPL_WIDTH - 1),
		4217 => to_unsigned(12890, LUT_AMPL_WIDTH - 1),
		4218 => to_unsigned(12893, LUT_AMPL_WIDTH - 1),
		4219 => to_unsigned(12895, LUT_AMPL_WIDTH - 1),
		4220 => to_unsigned(12898, LUT_AMPL_WIDTH - 1),
		4221 => to_unsigned(12901, LUT_AMPL_WIDTH - 1),
		4222 => to_unsigned(12904, LUT_AMPL_WIDTH - 1),
		4223 => to_unsigned(12907, LUT_AMPL_WIDTH - 1),
		4224 => to_unsigned(12910, LUT_AMPL_WIDTH - 1),
		4225 => to_unsigned(12913, LUT_AMPL_WIDTH - 1),
		4226 => to_unsigned(12916, LUT_AMPL_WIDTH - 1),
		4227 => to_unsigned(12919, LUT_AMPL_WIDTH - 1),
		4228 => to_unsigned(12921, LUT_AMPL_WIDTH - 1),
		4229 => to_unsigned(12924, LUT_AMPL_WIDTH - 1),
		4230 => to_unsigned(12927, LUT_AMPL_WIDTH - 1),
		4231 => to_unsigned(12930, LUT_AMPL_WIDTH - 1),
		4232 => to_unsigned(12933, LUT_AMPL_WIDTH - 1),
		4233 => to_unsigned(12936, LUT_AMPL_WIDTH - 1),
		4234 => to_unsigned(12939, LUT_AMPL_WIDTH - 1),
		4235 => to_unsigned(12942, LUT_AMPL_WIDTH - 1),
		4236 => to_unsigned(12945, LUT_AMPL_WIDTH - 1),
		4237 => to_unsigned(12947, LUT_AMPL_WIDTH - 1),
		4238 => to_unsigned(12950, LUT_AMPL_WIDTH - 1),
		4239 => to_unsigned(12953, LUT_AMPL_WIDTH - 1),
		4240 => to_unsigned(12956, LUT_AMPL_WIDTH - 1),
		4241 => to_unsigned(12959, LUT_AMPL_WIDTH - 1),
		4242 => to_unsigned(12962, LUT_AMPL_WIDTH - 1),
		4243 => to_unsigned(12965, LUT_AMPL_WIDTH - 1),
		4244 => to_unsigned(12968, LUT_AMPL_WIDTH - 1),
		4245 => to_unsigned(12971, LUT_AMPL_WIDTH - 1),
		4246 => to_unsigned(12973, LUT_AMPL_WIDTH - 1),
		4247 => to_unsigned(12976, LUT_AMPL_WIDTH - 1),
		4248 => to_unsigned(12979, LUT_AMPL_WIDTH - 1),
		4249 => to_unsigned(12982, LUT_AMPL_WIDTH - 1),
		4250 => to_unsigned(12985, LUT_AMPL_WIDTH - 1),
		4251 => to_unsigned(12988, LUT_AMPL_WIDTH - 1),
		4252 => to_unsigned(12991, LUT_AMPL_WIDTH - 1),
		4253 => to_unsigned(12994, LUT_AMPL_WIDTH - 1),
		4254 => to_unsigned(12997, LUT_AMPL_WIDTH - 1),
		4255 => to_unsigned(12999, LUT_AMPL_WIDTH - 1),
		4256 => to_unsigned(13002, LUT_AMPL_WIDTH - 1),
		4257 => to_unsigned(13005, LUT_AMPL_WIDTH - 1),
		4258 => to_unsigned(13008, LUT_AMPL_WIDTH - 1),
		4259 => to_unsigned(13011, LUT_AMPL_WIDTH - 1),
		4260 => to_unsigned(13014, LUT_AMPL_WIDTH - 1),
		4261 => to_unsigned(13017, LUT_AMPL_WIDTH - 1),
		4262 => to_unsigned(13020, LUT_AMPL_WIDTH - 1),
		4263 => to_unsigned(13022, LUT_AMPL_WIDTH - 1),
		4264 => to_unsigned(13025, LUT_AMPL_WIDTH - 1),
		4265 => to_unsigned(13028, LUT_AMPL_WIDTH - 1),
		4266 => to_unsigned(13031, LUT_AMPL_WIDTH - 1),
		4267 => to_unsigned(13034, LUT_AMPL_WIDTH - 1),
		4268 => to_unsigned(13037, LUT_AMPL_WIDTH - 1),
		4269 => to_unsigned(13040, LUT_AMPL_WIDTH - 1),
		4270 => to_unsigned(13043, LUT_AMPL_WIDTH - 1),
		4271 => to_unsigned(13046, LUT_AMPL_WIDTH - 1),
		4272 => to_unsigned(13048, LUT_AMPL_WIDTH - 1),
		4273 => to_unsigned(13051, LUT_AMPL_WIDTH - 1),
		4274 => to_unsigned(13054, LUT_AMPL_WIDTH - 1),
		4275 => to_unsigned(13057, LUT_AMPL_WIDTH - 1),
		4276 => to_unsigned(13060, LUT_AMPL_WIDTH - 1),
		4277 => to_unsigned(13063, LUT_AMPL_WIDTH - 1),
		4278 => to_unsigned(13066, LUT_AMPL_WIDTH - 1),
		4279 => to_unsigned(13069, LUT_AMPL_WIDTH - 1),
		4280 => to_unsigned(13071, LUT_AMPL_WIDTH - 1),
		4281 => to_unsigned(13074, LUT_AMPL_WIDTH - 1),
		4282 => to_unsigned(13077, LUT_AMPL_WIDTH - 1),
		4283 => to_unsigned(13080, LUT_AMPL_WIDTH - 1),
		4284 => to_unsigned(13083, LUT_AMPL_WIDTH - 1),
		4285 => to_unsigned(13086, LUT_AMPL_WIDTH - 1),
		4286 => to_unsigned(13089, LUT_AMPL_WIDTH - 1),
		4287 => to_unsigned(13092, LUT_AMPL_WIDTH - 1),
		4288 => to_unsigned(13094, LUT_AMPL_WIDTH - 1),
		4289 => to_unsigned(13097, LUT_AMPL_WIDTH - 1),
		4290 => to_unsigned(13100, LUT_AMPL_WIDTH - 1),
		4291 => to_unsigned(13103, LUT_AMPL_WIDTH - 1),
		4292 => to_unsigned(13106, LUT_AMPL_WIDTH - 1),
		4293 => to_unsigned(13109, LUT_AMPL_WIDTH - 1),
		4294 => to_unsigned(13112, LUT_AMPL_WIDTH - 1),
		4295 => to_unsigned(13115, LUT_AMPL_WIDTH - 1),
		4296 => to_unsigned(13118, LUT_AMPL_WIDTH - 1),
		4297 => to_unsigned(13120, LUT_AMPL_WIDTH - 1),
		4298 => to_unsigned(13123, LUT_AMPL_WIDTH - 1),
		4299 => to_unsigned(13126, LUT_AMPL_WIDTH - 1),
		4300 => to_unsigned(13129, LUT_AMPL_WIDTH - 1),
		4301 => to_unsigned(13132, LUT_AMPL_WIDTH - 1),
		4302 => to_unsigned(13135, LUT_AMPL_WIDTH - 1),
		4303 => to_unsigned(13138, LUT_AMPL_WIDTH - 1),
		4304 => to_unsigned(13141, LUT_AMPL_WIDTH - 1),
		4305 => to_unsigned(13143, LUT_AMPL_WIDTH - 1),
		4306 => to_unsigned(13146, LUT_AMPL_WIDTH - 1),
		4307 => to_unsigned(13149, LUT_AMPL_WIDTH - 1),
		4308 => to_unsigned(13152, LUT_AMPL_WIDTH - 1),
		4309 => to_unsigned(13155, LUT_AMPL_WIDTH - 1),
		4310 => to_unsigned(13158, LUT_AMPL_WIDTH - 1),
		4311 => to_unsigned(13161, LUT_AMPL_WIDTH - 1),
		4312 => to_unsigned(13164, LUT_AMPL_WIDTH - 1),
		4313 => to_unsigned(13166, LUT_AMPL_WIDTH - 1),
		4314 => to_unsigned(13169, LUT_AMPL_WIDTH - 1),
		4315 => to_unsigned(13172, LUT_AMPL_WIDTH - 1),
		4316 => to_unsigned(13175, LUT_AMPL_WIDTH - 1),
		4317 => to_unsigned(13178, LUT_AMPL_WIDTH - 1),
		4318 => to_unsigned(13181, LUT_AMPL_WIDTH - 1),
		4319 => to_unsigned(13184, LUT_AMPL_WIDTH - 1),
		4320 => to_unsigned(13187, LUT_AMPL_WIDTH - 1),
		4321 => to_unsigned(13189, LUT_AMPL_WIDTH - 1),
		4322 => to_unsigned(13192, LUT_AMPL_WIDTH - 1),
		4323 => to_unsigned(13195, LUT_AMPL_WIDTH - 1),
		4324 => to_unsigned(13198, LUT_AMPL_WIDTH - 1),
		4325 => to_unsigned(13201, LUT_AMPL_WIDTH - 1),
		4326 => to_unsigned(13204, LUT_AMPL_WIDTH - 1),
		4327 => to_unsigned(13207, LUT_AMPL_WIDTH - 1),
		4328 => to_unsigned(13210, LUT_AMPL_WIDTH - 1),
		4329 => to_unsigned(13212, LUT_AMPL_WIDTH - 1),
		4330 => to_unsigned(13215, LUT_AMPL_WIDTH - 1),
		4331 => to_unsigned(13218, LUT_AMPL_WIDTH - 1),
		4332 => to_unsigned(13221, LUT_AMPL_WIDTH - 1),
		4333 => to_unsigned(13224, LUT_AMPL_WIDTH - 1),
		4334 => to_unsigned(13227, LUT_AMPL_WIDTH - 1),
		4335 => to_unsigned(13230, LUT_AMPL_WIDTH - 1),
		4336 => to_unsigned(13233, LUT_AMPL_WIDTH - 1),
		4337 => to_unsigned(13235, LUT_AMPL_WIDTH - 1),
		4338 => to_unsigned(13238, LUT_AMPL_WIDTH - 1),
		4339 => to_unsigned(13241, LUT_AMPL_WIDTH - 1),
		4340 => to_unsigned(13244, LUT_AMPL_WIDTH - 1),
		4341 => to_unsigned(13247, LUT_AMPL_WIDTH - 1),
		4342 => to_unsigned(13250, LUT_AMPL_WIDTH - 1),
		4343 => to_unsigned(13253, LUT_AMPL_WIDTH - 1),
		4344 => to_unsigned(13256, LUT_AMPL_WIDTH - 1),
		4345 => to_unsigned(13258, LUT_AMPL_WIDTH - 1),
		4346 => to_unsigned(13261, LUT_AMPL_WIDTH - 1),
		4347 => to_unsigned(13264, LUT_AMPL_WIDTH - 1),
		4348 => to_unsigned(13267, LUT_AMPL_WIDTH - 1),
		4349 => to_unsigned(13270, LUT_AMPL_WIDTH - 1),
		4350 => to_unsigned(13273, LUT_AMPL_WIDTH - 1),
		4351 => to_unsigned(13276, LUT_AMPL_WIDTH - 1),
		4352 => to_unsigned(13279, LUT_AMPL_WIDTH - 1),
		4353 => to_unsigned(13281, LUT_AMPL_WIDTH - 1),
		4354 => to_unsigned(13284, LUT_AMPL_WIDTH - 1),
		4355 => to_unsigned(13287, LUT_AMPL_WIDTH - 1),
		4356 => to_unsigned(13290, LUT_AMPL_WIDTH - 1),
		4357 => to_unsigned(13293, LUT_AMPL_WIDTH - 1),
		4358 => to_unsigned(13296, LUT_AMPL_WIDTH - 1),
		4359 => to_unsigned(13299, LUT_AMPL_WIDTH - 1),
		4360 => to_unsigned(13302, LUT_AMPL_WIDTH - 1),
		4361 => to_unsigned(13304, LUT_AMPL_WIDTH - 1),
		4362 => to_unsigned(13307, LUT_AMPL_WIDTH - 1),
		4363 => to_unsigned(13310, LUT_AMPL_WIDTH - 1),
		4364 => to_unsigned(13313, LUT_AMPL_WIDTH - 1),
		4365 => to_unsigned(13316, LUT_AMPL_WIDTH - 1),
		4366 => to_unsigned(13319, LUT_AMPL_WIDTH - 1),
		4367 => to_unsigned(13322, LUT_AMPL_WIDTH - 1),
		4368 => to_unsigned(13324, LUT_AMPL_WIDTH - 1),
		4369 => to_unsigned(13327, LUT_AMPL_WIDTH - 1),
		4370 => to_unsigned(13330, LUT_AMPL_WIDTH - 1),
		4371 => to_unsigned(13333, LUT_AMPL_WIDTH - 1),
		4372 => to_unsigned(13336, LUT_AMPL_WIDTH - 1),
		4373 => to_unsigned(13339, LUT_AMPL_WIDTH - 1),
		4374 => to_unsigned(13342, LUT_AMPL_WIDTH - 1),
		4375 => to_unsigned(13345, LUT_AMPL_WIDTH - 1),
		4376 => to_unsigned(13347, LUT_AMPL_WIDTH - 1),
		4377 => to_unsigned(13350, LUT_AMPL_WIDTH - 1),
		4378 => to_unsigned(13353, LUT_AMPL_WIDTH - 1),
		4379 => to_unsigned(13356, LUT_AMPL_WIDTH - 1),
		4380 => to_unsigned(13359, LUT_AMPL_WIDTH - 1),
		4381 => to_unsigned(13362, LUT_AMPL_WIDTH - 1),
		4382 => to_unsigned(13365, LUT_AMPL_WIDTH - 1),
		4383 => to_unsigned(13368, LUT_AMPL_WIDTH - 1),
		4384 => to_unsigned(13370, LUT_AMPL_WIDTH - 1),
		4385 => to_unsigned(13373, LUT_AMPL_WIDTH - 1),
		4386 => to_unsigned(13376, LUT_AMPL_WIDTH - 1),
		4387 => to_unsigned(13379, LUT_AMPL_WIDTH - 1),
		4388 => to_unsigned(13382, LUT_AMPL_WIDTH - 1),
		4389 => to_unsigned(13385, LUT_AMPL_WIDTH - 1),
		4390 => to_unsigned(13388, LUT_AMPL_WIDTH - 1),
		4391 => to_unsigned(13390, LUT_AMPL_WIDTH - 1),
		4392 => to_unsigned(13393, LUT_AMPL_WIDTH - 1),
		4393 => to_unsigned(13396, LUT_AMPL_WIDTH - 1),
		4394 => to_unsigned(13399, LUT_AMPL_WIDTH - 1),
		4395 => to_unsigned(13402, LUT_AMPL_WIDTH - 1),
		4396 => to_unsigned(13405, LUT_AMPL_WIDTH - 1),
		4397 => to_unsigned(13408, LUT_AMPL_WIDTH - 1),
		4398 => to_unsigned(13411, LUT_AMPL_WIDTH - 1),
		4399 => to_unsigned(13413, LUT_AMPL_WIDTH - 1),
		4400 => to_unsigned(13416, LUT_AMPL_WIDTH - 1),
		4401 => to_unsigned(13419, LUT_AMPL_WIDTH - 1),
		4402 => to_unsigned(13422, LUT_AMPL_WIDTH - 1),
		4403 => to_unsigned(13425, LUT_AMPL_WIDTH - 1),
		4404 => to_unsigned(13428, LUT_AMPL_WIDTH - 1),
		4405 => to_unsigned(13431, LUT_AMPL_WIDTH - 1),
		4406 => to_unsigned(13433, LUT_AMPL_WIDTH - 1),
		4407 => to_unsigned(13436, LUT_AMPL_WIDTH - 1),
		4408 => to_unsigned(13439, LUT_AMPL_WIDTH - 1),
		4409 => to_unsigned(13442, LUT_AMPL_WIDTH - 1),
		4410 => to_unsigned(13445, LUT_AMPL_WIDTH - 1),
		4411 => to_unsigned(13448, LUT_AMPL_WIDTH - 1),
		4412 => to_unsigned(13451, LUT_AMPL_WIDTH - 1),
		4413 => to_unsigned(13454, LUT_AMPL_WIDTH - 1),
		4414 => to_unsigned(13456, LUT_AMPL_WIDTH - 1),
		4415 => to_unsigned(13459, LUT_AMPL_WIDTH - 1),
		4416 => to_unsigned(13462, LUT_AMPL_WIDTH - 1),
		4417 => to_unsigned(13465, LUT_AMPL_WIDTH - 1),
		4418 => to_unsigned(13468, LUT_AMPL_WIDTH - 1),
		4419 => to_unsigned(13471, LUT_AMPL_WIDTH - 1),
		4420 => to_unsigned(13474, LUT_AMPL_WIDTH - 1),
		4421 => to_unsigned(13476, LUT_AMPL_WIDTH - 1),
		4422 => to_unsigned(13479, LUT_AMPL_WIDTH - 1),
		4423 => to_unsigned(13482, LUT_AMPL_WIDTH - 1),
		4424 => to_unsigned(13485, LUT_AMPL_WIDTH - 1),
		4425 => to_unsigned(13488, LUT_AMPL_WIDTH - 1),
		4426 => to_unsigned(13491, LUT_AMPL_WIDTH - 1),
		4427 => to_unsigned(13494, LUT_AMPL_WIDTH - 1),
		4428 => to_unsigned(13496, LUT_AMPL_WIDTH - 1),
		4429 => to_unsigned(13499, LUT_AMPL_WIDTH - 1),
		4430 => to_unsigned(13502, LUT_AMPL_WIDTH - 1),
		4431 => to_unsigned(13505, LUT_AMPL_WIDTH - 1),
		4432 => to_unsigned(13508, LUT_AMPL_WIDTH - 1),
		4433 => to_unsigned(13511, LUT_AMPL_WIDTH - 1),
		4434 => to_unsigned(13514, LUT_AMPL_WIDTH - 1),
		4435 => to_unsigned(13516, LUT_AMPL_WIDTH - 1),
		4436 => to_unsigned(13519, LUT_AMPL_WIDTH - 1),
		4437 => to_unsigned(13522, LUT_AMPL_WIDTH - 1),
		4438 => to_unsigned(13525, LUT_AMPL_WIDTH - 1),
		4439 => to_unsigned(13528, LUT_AMPL_WIDTH - 1),
		4440 => to_unsigned(13531, LUT_AMPL_WIDTH - 1),
		4441 => to_unsigned(13534, LUT_AMPL_WIDTH - 1),
		4442 => to_unsigned(13537, LUT_AMPL_WIDTH - 1),
		4443 => to_unsigned(13539, LUT_AMPL_WIDTH - 1),
		4444 => to_unsigned(13542, LUT_AMPL_WIDTH - 1),
		4445 => to_unsigned(13545, LUT_AMPL_WIDTH - 1),
		4446 => to_unsigned(13548, LUT_AMPL_WIDTH - 1),
		4447 => to_unsigned(13551, LUT_AMPL_WIDTH - 1),
		4448 => to_unsigned(13554, LUT_AMPL_WIDTH - 1),
		4449 => to_unsigned(13557, LUT_AMPL_WIDTH - 1),
		4450 => to_unsigned(13559, LUT_AMPL_WIDTH - 1),
		4451 => to_unsigned(13562, LUT_AMPL_WIDTH - 1),
		4452 => to_unsigned(13565, LUT_AMPL_WIDTH - 1),
		4453 => to_unsigned(13568, LUT_AMPL_WIDTH - 1),
		4454 => to_unsigned(13571, LUT_AMPL_WIDTH - 1),
		4455 => to_unsigned(13574, LUT_AMPL_WIDTH - 1),
		4456 => to_unsigned(13577, LUT_AMPL_WIDTH - 1),
		4457 => to_unsigned(13579, LUT_AMPL_WIDTH - 1),
		4458 => to_unsigned(13582, LUT_AMPL_WIDTH - 1),
		4459 => to_unsigned(13585, LUT_AMPL_WIDTH - 1),
		4460 => to_unsigned(13588, LUT_AMPL_WIDTH - 1),
		4461 => to_unsigned(13591, LUT_AMPL_WIDTH - 1),
		4462 => to_unsigned(13594, LUT_AMPL_WIDTH - 1),
		4463 => to_unsigned(13597, LUT_AMPL_WIDTH - 1),
		4464 => to_unsigned(13599, LUT_AMPL_WIDTH - 1),
		4465 => to_unsigned(13602, LUT_AMPL_WIDTH - 1),
		4466 => to_unsigned(13605, LUT_AMPL_WIDTH - 1),
		4467 => to_unsigned(13608, LUT_AMPL_WIDTH - 1),
		4468 => to_unsigned(13611, LUT_AMPL_WIDTH - 1),
		4469 => to_unsigned(13614, LUT_AMPL_WIDTH - 1),
		4470 => to_unsigned(13617, LUT_AMPL_WIDTH - 1),
		4471 => to_unsigned(13619, LUT_AMPL_WIDTH - 1),
		4472 => to_unsigned(13622, LUT_AMPL_WIDTH - 1),
		4473 => to_unsigned(13625, LUT_AMPL_WIDTH - 1),
		4474 => to_unsigned(13628, LUT_AMPL_WIDTH - 1),
		4475 => to_unsigned(13631, LUT_AMPL_WIDTH - 1),
		4476 => to_unsigned(13634, LUT_AMPL_WIDTH - 1),
		4477 => to_unsigned(13637, LUT_AMPL_WIDTH - 1),
		4478 => to_unsigned(13639, LUT_AMPL_WIDTH - 1),
		4479 => to_unsigned(13642, LUT_AMPL_WIDTH - 1),
		4480 => to_unsigned(13645, LUT_AMPL_WIDTH - 1),
		4481 => to_unsigned(13648, LUT_AMPL_WIDTH - 1),
		4482 => to_unsigned(13651, LUT_AMPL_WIDTH - 1),
		4483 => to_unsigned(13654, LUT_AMPL_WIDTH - 1),
		4484 => to_unsigned(13657, LUT_AMPL_WIDTH - 1),
		4485 => to_unsigned(13659, LUT_AMPL_WIDTH - 1),
		4486 => to_unsigned(13662, LUT_AMPL_WIDTH - 1),
		4487 => to_unsigned(13665, LUT_AMPL_WIDTH - 1),
		4488 => to_unsigned(13668, LUT_AMPL_WIDTH - 1),
		4489 => to_unsigned(13671, LUT_AMPL_WIDTH - 1),
		4490 => to_unsigned(13674, LUT_AMPL_WIDTH - 1),
		4491 => to_unsigned(13677, LUT_AMPL_WIDTH - 1),
		4492 => to_unsigned(13679, LUT_AMPL_WIDTH - 1),
		4493 => to_unsigned(13682, LUT_AMPL_WIDTH - 1),
		4494 => to_unsigned(13685, LUT_AMPL_WIDTH - 1),
		4495 => to_unsigned(13688, LUT_AMPL_WIDTH - 1),
		4496 => to_unsigned(13691, LUT_AMPL_WIDTH - 1),
		4497 => to_unsigned(13694, LUT_AMPL_WIDTH - 1),
		4498 => to_unsigned(13697, LUT_AMPL_WIDTH - 1),
		4499 => to_unsigned(13699, LUT_AMPL_WIDTH - 1),
		4500 => to_unsigned(13702, LUT_AMPL_WIDTH - 1),
		4501 => to_unsigned(13705, LUT_AMPL_WIDTH - 1),
		4502 => to_unsigned(13708, LUT_AMPL_WIDTH - 1),
		4503 => to_unsigned(13711, LUT_AMPL_WIDTH - 1),
		4504 => to_unsigned(13714, LUT_AMPL_WIDTH - 1),
		4505 => to_unsigned(13717, LUT_AMPL_WIDTH - 1),
		4506 => to_unsigned(13719, LUT_AMPL_WIDTH - 1),
		4507 => to_unsigned(13722, LUT_AMPL_WIDTH - 1),
		4508 => to_unsigned(13725, LUT_AMPL_WIDTH - 1),
		4509 => to_unsigned(13728, LUT_AMPL_WIDTH - 1),
		4510 => to_unsigned(13731, LUT_AMPL_WIDTH - 1),
		4511 => to_unsigned(13734, LUT_AMPL_WIDTH - 1),
		4512 => to_unsigned(13736, LUT_AMPL_WIDTH - 1),
		4513 => to_unsigned(13739, LUT_AMPL_WIDTH - 1),
		4514 => to_unsigned(13742, LUT_AMPL_WIDTH - 1),
		4515 => to_unsigned(13745, LUT_AMPL_WIDTH - 1),
		4516 => to_unsigned(13748, LUT_AMPL_WIDTH - 1),
		4517 => to_unsigned(13751, LUT_AMPL_WIDTH - 1),
		4518 => to_unsigned(13754, LUT_AMPL_WIDTH - 1),
		4519 => to_unsigned(13756, LUT_AMPL_WIDTH - 1),
		4520 => to_unsigned(13759, LUT_AMPL_WIDTH - 1),
		4521 => to_unsigned(13762, LUT_AMPL_WIDTH - 1),
		4522 => to_unsigned(13765, LUT_AMPL_WIDTH - 1),
		4523 => to_unsigned(13768, LUT_AMPL_WIDTH - 1),
		4524 => to_unsigned(13771, LUT_AMPL_WIDTH - 1),
		4525 => to_unsigned(13774, LUT_AMPL_WIDTH - 1),
		4526 => to_unsigned(13776, LUT_AMPL_WIDTH - 1),
		4527 => to_unsigned(13779, LUT_AMPL_WIDTH - 1),
		4528 => to_unsigned(13782, LUT_AMPL_WIDTH - 1),
		4529 => to_unsigned(13785, LUT_AMPL_WIDTH - 1),
		4530 => to_unsigned(13788, LUT_AMPL_WIDTH - 1),
		4531 => to_unsigned(13791, LUT_AMPL_WIDTH - 1),
		4532 => to_unsigned(13793, LUT_AMPL_WIDTH - 1),
		4533 => to_unsigned(13796, LUT_AMPL_WIDTH - 1),
		4534 => to_unsigned(13799, LUT_AMPL_WIDTH - 1),
		4535 => to_unsigned(13802, LUT_AMPL_WIDTH - 1),
		4536 => to_unsigned(13805, LUT_AMPL_WIDTH - 1),
		4537 => to_unsigned(13808, LUT_AMPL_WIDTH - 1),
		4538 => to_unsigned(13811, LUT_AMPL_WIDTH - 1),
		4539 => to_unsigned(13813, LUT_AMPL_WIDTH - 1),
		4540 => to_unsigned(13816, LUT_AMPL_WIDTH - 1),
		4541 => to_unsigned(13819, LUT_AMPL_WIDTH - 1),
		4542 => to_unsigned(13822, LUT_AMPL_WIDTH - 1),
		4543 => to_unsigned(13825, LUT_AMPL_WIDTH - 1),
		4544 => to_unsigned(13828, LUT_AMPL_WIDTH - 1),
		4545 => to_unsigned(13831, LUT_AMPL_WIDTH - 1),
		4546 => to_unsigned(13833, LUT_AMPL_WIDTH - 1),
		4547 => to_unsigned(13836, LUT_AMPL_WIDTH - 1),
		4548 => to_unsigned(13839, LUT_AMPL_WIDTH - 1),
		4549 => to_unsigned(13842, LUT_AMPL_WIDTH - 1),
		4550 => to_unsigned(13845, LUT_AMPL_WIDTH - 1),
		4551 => to_unsigned(13848, LUT_AMPL_WIDTH - 1),
		4552 => to_unsigned(13850, LUT_AMPL_WIDTH - 1),
		4553 => to_unsigned(13853, LUT_AMPL_WIDTH - 1),
		4554 => to_unsigned(13856, LUT_AMPL_WIDTH - 1),
		4555 => to_unsigned(13859, LUT_AMPL_WIDTH - 1),
		4556 => to_unsigned(13862, LUT_AMPL_WIDTH - 1),
		4557 => to_unsigned(13865, LUT_AMPL_WIDTH - 1),
		4558 => to_unsigned(13868, LUT_AMPL_WIDTH - 1),
		4559 => to_unsigned(13870, LUT_AMPL_WIDTH - 1),
		4560 => to_unsigned(13873, LUT_AMPL_WIDTH - 1),
		4561 => to_unsigned(13876, LUT_AMPL_WIDTH - 1),
		4562 => to_unsigned(13879, LUT_AMPL_WIDTH - 1),
		4563 => to_unsigned(13882, LUT_AMPL_WIDTH - 1),
		4564 => to_unsigned(13885, LUT_AMPL_WIDTH - 1),
		4565 => to_unsigned(13887, LUT_AMPL_WIDTH - 1),
		4566 => to_unsigned(13890, LUT_AMPL_WIDTH - 1),
		4567 => to_unsigned(13893, LUT_AMPL_WIDTH - 1),
		4568 => to_unsigned(13896, LUT_AMPL_WIDTH - 1),
		4569 => to_unsigned(13899, LUT_AMPL_WIDTH - 1),
		4570 => to_unsigned(13902, LUT_AMPL_WIDTH - 1),
		4571 => to_unsigned(13905, LUT_AMPL_WIDTH - 1),
		4572 => to_unsigned(13907, LUT_AMPL_WIDTH - 1),
		4573 => to_unsigned(13910, LUT_AMPL_WIDTH - 1),
		4574 => to_unsigned(13913, LUT_AMPL_WIDTH - 1),
		4575 => to_unsigned(13916, LUT_AMPL_WIDTH - 1),
		4576 => to_unsigned(13919, LUT_AMPL_WIDTH - 1),
		4577 => to_unsigned(13922, LUT_AMPL_WIDTH - 1),
		4578 => to_unsigned(13924, LUT_AMPL_WIDTH - 1),
		4579 => to_unsigned(13927, LUT_AMPL_WIDTH - 1),
		4580 => to_unsigned(13930, LUT_AMPL_WIDTH - 1),
		4581 => to_unsigned(13933, LUT_AMPL_WIDTH - 1),
		4582 => to_unsigned(13936, LUT_AMPL_WIDTH - 1),
		4583 => to_unsigned(13939, LUT_AMPL_WIDTH - 1),
		4584 => to_unsigned(13942, LUT_AMPL_WIDTH - 1),
		4585 => to_unsigned(13944, LUT_AMPL_WIDTH - 1),
		4586 => to_unsigned(13947, LUT_AMPL_WIDTH - 1),
		4587 => to_unsigned(13950, LUT_AMPL_WIDTH - 1),
		4588 => to_unsigned(13953, LUT_AMPL_WIDTH - 1),
		4589 => to_unsigned(13956, LUT_AMPL_WIDTH - 1),
		4590 => to_unsigned(13959, LUT_AMPL_WIDTH - 1),
		4591 => to_unsigned(13961, LUT_AMPL_WIDTH - 1),
		4592 => to_unsigned(13964, LUT_AMPL_WIDTH - 1),
		4593 => to_unsigned(13967, LUT_AMPL_WIDTH - 1),
		4594 => to_unsigned(13970, LUT_AMPL_WIDTH - 1),
		4595 => to_unsigned(13973, LUT_AMPL_WIDTH - 1),
		4596 => to_unsigned(13976, LUT_AMPL_WIDTH - 1),
		4597 => to_unsigned(13978, LUT_AMPL_WIDTH - 1),
		4598 => to_unsigned(13981, LUT_AMPL_WIDTH - 1),
		4599 => to_unsigned(13984, LUT_AMPL_WIDTH - 1),
		4600 => to_unsigned(13987, LUT_AMPL_WIDTH - 1),
		4601 => to_unsigned(13990, LUT_AMPL_WIDTH - 1),
		4602 => to_unsigned(13993, LUT_AMPL_WIDTH - 1),
		4603 => to_unsigned(13995, LUT_AMPL_WIDTH - 1),
		4604 => to_unsigned(13998, LUT_AMPL_WIDTH - 1),
		4605 => to_unsigned(14001, LUT_AMPL_WIDTH - 1),
		4606 => to_unsigned(14004, LUT_AMPL_WIDTH - 1),
		4607 => to_unsigned(14007, LUT_AMPL_WIDTH - 1),
		4608 => to_unsigned(14010, LUT_AMPL_WIDTH - 1),
		4609 => to_unsigned(14013, LUT_AMPL_WIDTH - 1),
		4610 => to_unsigned(14015, LUT_AMPL_WIDTH - 1),
		4611 => to_unsigned(14018, LUT_AMPL_WIDTH - 1),
		4612 => to_unsigned(14021, LUT_AMPL_WIDTH - 1),
		4613 => to_unsigned(14024, LUT_AMPL_WIDTH - 1),
		4614 => to_unsigned(14027, LUT_AMPL_WIDTH - 1),
		4615 => to_unsigned(14030, LUT_AMPL_WIDTH - 1),
		4616 => to_unsigned(14032, LUT_AMPL_WIDTH - 1),
		4617 => to_unsigned(14035, LUT_AMPL_WIDTH - 1),
		4618 => to_unsigned(14038, LUT_AMPL_WIDTH - 1),
		4619 => to_unsigned(14041, LUT_AMPL_WIDTH - 1),
		4620 => to_unsigned(14044, LUT_AMPL_WIDTH - 1),
		4621 => to_unsigned(14047, LUT_AMPL_WIDTH - 1),
		4622 => to_unsigned(14049, LUT_AMPL_WIDTH - 1),
		4623 => to_unsigned(14052, LUT_AMPL_WIDTH - 1),
		4624 => to_unsigned(14055, LUT_AMPL_WIDTH - 1),
		4625 => to_unsigned(14058, LUT_AMPL_WIDTH - 1),
		4626 => to_unsigned(14061, LUT_AMPL_WIDTH - 1),
		4627 => to_unsigned(14064, LUT_AMPL_WIDTH - 1),
		4628 => to_unsigned(14066, LUT_AMPL_WIDTH - 1),
		4629 => to_unsigned(14069, LUT_AMPL_WIDTH - 1),
		4630 => to_unsigned(14072, LUT_AMPL_WIDTH - 1),
		4631 => to_unsigned(14075, LUT_AMPL_WIDTH - 1),
		4632 => to_unsigned(14078, LUT_AMPL_WIDTH - 1),
		4633 => to_unsigned(14081, LUT_AMPL_WIDTH - 1),
		4634 => to_unsigned(14083, LUT_AMPL_WIDTH - 1),
		4635 => to_unsigned(14086, LUT_AMPL_WIDTH - 1),
		4636 => to_unsigned(14089, LUT_AMPL_WIDTH - 1),
		4637 => to_unsigned(14092, LUT_AMPL_WIDTH - 1),
		4638 => to_unsigned(14095, LUT_AMPL_WIDTH - 1),
		4639 => to_unsigned(14098, LUT_AMPL_WIDTH - 1),
		4640 => to_unsigned(14101, LUT_AMPL_WIDTH - 1),
		4641 => to_unsigned(14103, LUT_AMPL_WIDTH - 1),
		4642 => to_unsigned(14106, LUT_AMPL_WIDTH - 1),
		4643 => to_unsigned(14109, LUT_AMPL_WIDTH - 1),
		4644 => to_unsigned(14112, LUT_AMPL_WIDTH - 1),
		4645 => to_unsigned(14115, LUT_AMPL_WIDTH - 1),
		4646 => to_unsigned(14118, LUT_AMPL_WIDTH - 1),
		4647 => to_unsigned(14120, LUT_AMPL_WIDTH - 1),
		4648 => to_unsigned(14123, LUT_AMPL_WIDTH - 1),
		4649 => to_unsigned(14126, LUT_AMPL_WIDTH - 1),
		4650 => to_unsigned(14129, LUT_AMPL_WIDTH - 1),
		4651 => to_unsigned(14132, LUT_AMPL_WIDTH - 1),
		4652 => to_unsigned(14135, LUT_AMPL_WIDTH - 1),
		4653 => to_unsigned(14137, LUT_AMPL_WIDTH - 1),
		4654 => to_unsigned(14140, LUT_AMPL_WIDTH - 1),
		4655 => to_unsigned(14143, LUT_AMPL_WIDTH - 1),
		4656 => to_unsigned(14146, LUT_AMPL_WIDTH - 1),
		4657 => to_unsigned(14149, LUT_AMPL_WIDTH - 1),
		4658 => to_unsigned(14152, LUT_AMPL_WIDTH - 1),
		4659 => to_unsigned(14154, LUT_AMPL_WIDTH - 1),
		4660 => to_unsigned(14157, LUT_AMPL_WIDTH - 1),
		4661 => to_unsigned(14160, LUT_AMPL_WIDTH - 1),
		4662 => to_unsigned(14163, LUT_AMPL_WIDTH - 1),
		4663 => to_unsigned(14166, LUT_AMPL_WIDTH - 1),
		4664 => to_unsigned(14169, LUT_AMPL_WIDTH - 1),
		4665 => to_unsigned(14171, LUT_AMPL_WIDTH - 1),
		4666 => to_unsigned(14174, LUT_AMPL_WIDTH - 1),
		4667 => to_unsigned(14177, LUT_AMPL_WIDTH - 1),
		4668 => to_unsigned(14180, LUT_AMPL_WIDTH - 1),
		4669 => to_unsigned(14183, LUT_AMPL_WIDTH - 1),
		4670 => to_unsigned(14186, LUT_AMPL_WIDTH - 1),
		4671 => to_unsigned(14188, LUT_AMPL_WIDTH - 1),
		4672 => to_unsigned(14191, LUT_AMPL_WIDTH - 1),
		4673 => to_unsigned(14194, LUT_AMPL_WIDTH - 1),
		4674 => to_unsigned(14197, LUT_AMPL_WIDTH - 1),
		4675 => to_unsigned(14200, LUT_AMPL_WIDTH - 1),
		4676 => to_unsigned(14203, LUT_AMPL_WIDTH - 1),
		4677 => to_unsigned(14205, LUT_AMPL_WIDTH - 1),
		4678 => to_unsigned(14208, LUT_AMPL_WIDTH - 1),
		4679 => to_unsigned(14211, LUT_AMPL_WIDTH - 1),
		4680 => to_unsigned(14214, LUT_AMPL_WIDTH - 1),
		4681 => to_unsigned(14217, LUT_AMPL_WIDTH - 1),
		4682 => to_unsigned(14219, LUT_AMPL_WIDTH - 1),
		4683 => to_unsigned(14222, LUT_AMPL_WIDTH - 1),
		4684 => to_unsigned(14225, LUT_AMPL_WIDTH - 1),
		4685 => to_unsigned(14228, LUT_AMPL_WIDTH - 1),
		4686 => to_unsigned(14231, LUT_AMPL_WIDTH - 1),
		4687 => to_unsigned(14234, LUT_AMPL_WIDTH - 1),
		4688 => to_unsigned(14236, LUT_AMPL_WIDTH - 1),
		4689 => to_unsigned(14239, LUT_AMPL_WIDTH - 1),
		4690 => to_unsigned(14242, LUT_AMPL_WIDTH - 1),
		4691 => to_unsigned(14245, LUT_AMPL_WIDTH - 1),
		4692 => to_unsigned(14248, LUT_AMPL_WIDTH - 1),
		4693 => to_unsigned(14251, LUT_AMPL_WIDTH - 1),
		4694 => to_unsigned(14253, LUT_AMPL_WIDTH - 1),
		4695 => to_unsigned(14256, LUT_AMPL_WIDTH - 1),
		4696 => to_unsigned(14259, LUT_AMPL_WIDTH - 1),
		4697 => to_unsigned(14262, LUT_AMPL_WIDTH - 1),
		4698 => to_unsigned(14265, LUT_AMPL_WIDTH - 1),
		4699 => to_unsigned(14268, LUT_AMPL_WIDTH - 1),
		4700 => to_unsigned(14270, LUT_AMPL_WIDTH - 1),
		4701 => to_unsigned(14273, LUT_AMPL_WIDTH - 1),
		4702 => to_unsigned(14276, LUT_AMPL_WIDTH - 1),
		4703 => to_unsigned(14279, LUT_AMPL_WIDTH - 1),
		4704 => to_unsigned(14282, LUT_AMPL_WIDTH - 1),
		4705 => to_unsigned(14285, LUT_AMPL_WIDTH - 1),
		4706 => to_unsigned(14287, LUT_AMPL_WIDTH - 1),
		4707 => to_unsigned(14290, LUT_AMPL_WIDTH - 1),
		4708 => to_unsigned(14293, LUT_AMPL_WIDTH - 1),
		4709 => to_unsigned(14296, LUT_AMPL_WIDTH - 1),
		4710 => to_unsigned(14299, LUT_AMPL_WIDTH - 1),
		4711 => to_unsigned(14302, LUT_AMPL_WIDTH - 1),
		4712 => to_unsigned(14304, LUT_AMPL_WIDTH - 1),
		4713 => to_unsigned(14307, LUT_AMPL_WIDTH - 1),
		4714 => to_unsigned(14310, LUT_AMPL_WIDTH - 1),
		4715 => to_unsigned(14313, LUT_AMPL_WIDTH - 1),
		4716 => to_unsigned(14316, LUT_AMPL_WIDTH - 1),
		4717 => to_unsigned(14318, LUT_AMPL_WIDTH - 1),
		4718 => to_unsigned(14321, LUT_AMPL_WIDTH - 1),
		4719 => to_unsigned(14324, LUT_AMPL_WIDTH - 1),
		4720 => to_unsigned(14327, LUT_AMPL_WIDTH - 1),
		4721 => to_unsigned(14330, LUT_AMPL_WIDTH - 1),
		4722 => to_unsigned(14333, LUT_AMPL_WIDTH - 1),
		4723 => to_unsigned(14335, LUT_AMPL_WIDTH - 1),
		4724 => to_unsigned(14338, LUT_AMPL_WIDTH - 1),
		4725 => to_unsigned(14341, LUT_AMPL_WIDTH - 1),
		4726 => to_unsigned(14344, LUT_AMPL_WIDTH - 1),
		4727 => to_unsigned(14347, LUT_AMPL_WIDTH - 1),
		4728 => to_unsigned(14350, LUT_AMPL_WIDTH - 1),
		4729 => to_unsigned(14352, LUT_AMPL_WIDTH - 1),
		4730 => to_unsigned(14355, LUT_AMPL_WIDTH - 1),
		4731 => to_unsigned(14358, LUT_AMPL_WIDTH - 1),
		4732 => to_unsigned(14361, LUT_AMPL_WIDTH - 1),
		4733 => to_unsigned(14364, LUT_AMPL_WIDTH - 1),
		4734 => to_unsigned(14366, LUT_AMPL_WIDTH - 1),
		4735 => to_unsigned(14369, LUT_AMPL_WIDTH - 1),
		4736 => to_unsigned(14372, LUT_AMPL_WIDTH - 1),
		4737 => to_unsigned(14375, LUT_AMPL_WIDTH - 1),
		4738 => to_unsigned(14378, LUT_AMPL_WIDTH - 1),
		4739 => to_unsigned(14381, LUT_AMPL_WIDTH - 1),
		4740 => to_unsigned(14383, LUT_AMPL_WIDTH - 1),
		4741 => to_unsigned(14386, LUT_AMPL_WIDTH - 1),
		4742 => to_unsigned(14389, LUT_AMPL_WIDTH - 1),
		4743 => to_unsigned(14392, LUT_AMPL_WIDTH - 1),
		4744 => to_unsigned(14395, LUT_AMPL_WIDTH - 1),
		4745 => to_unsigned(14398, LUT_AMPL_WIDTH - 1),
		4746 => to_unsigned(14400, LUT_AMPL_WIDTH - 1),
		4747 => to_unsigned(14403, LUT_AMPL_WIDTH - 1),
		4748 => to_unsigned(14406, LUT_AMPL_WIDTH - 1),
		4749 => to_unsigned(14409, LUT_AMPL_WIDTH - 1),
		4750 => to_unsigned(14412, LUT_AMPL_WIDTH - 1),
		4751 => to_unsigned(14414, LUT_AMPL_WIDTH - 1),
		4752 => to_unsigned(14417, LUT_AMPL_WIDTH - 1),
		4753 => to_unsigned(14420, LUT_AMPL_WIDTH - 1),
		4754 => to_unsigned(14423, LUT_AMPL_WIDTH - 1),
		4755 => to_unsigned(14426, LUT_AMPL_WIDTH - 1),
		4756 => to_unsigned(14429, LUT_AMPL_WIDTH - 1),
		4757 => to_unsigned(14431, LUT_AMPL_WIDTH - 1),
		4758 => to_unsigned(14434, LUT_AMPL_WIDTH - 1),
		4759 => to_unsigned(14437, LUT_AMPL_WIDTH - 1),
		4760 => to_unsigned(14440, LUT_AMPL_WIDTH - 1),
		4761 => to_unsigned(14443, LUT_AMPL_WIDTH - 1),
		4762 => to_unsigned(14445, LUT_AMPL_WIDTH - 1),
		4763 => to_unsigned(14448, LUT_AMPL_WIDTH - 1),
		4764 => to_unsigned(14451, LUT_AMPL_WIDTH - 1),
		4765 => to_unsigned(14454, LUT_AMPL_WIDTH - 1),
		4766 => to_unsigned(14457, LUT_AMPL_WIDTH - 1),
		4767 => to_unsigned(14460, LUT_AMPL_WIDTH - 1),
		4768 => to_unsigned(14462, LUT_AMPL_WIDTH - 1),
		4769 => to_unsigned(14465, LUT_AMPL_WIDTH - 1),
		4770 => to_unsigned(14468, LUT_AMPL_WIDTH - 1),
		4771 => to_unsigned(14471, LUT_AMPL_WIDTH - 1),
		4772 => to_unsigned(14474, LUT_AMPL_WIDTH - 1),
		4773 => to_unsigned(14477, LUT_AMPL_WIDTH - 1),
		4774 => to_unsigned(14479, LUT_AMPL_WIDTH - 1),
		4775 => to_unsigned(14482, LUT_AMPL_WIDTH - 1),
		4776 => to_unsigned(14485, LUT_AMPL_WIDTH - 1),
		4777 => to_unsigned(14488, LUT_AMPL_WIDTH - 1),
		4778 => to_unsigned(14491, LUT_AMPL_WIDTH - 1),
		4779 => to_unsigned(14493, LUT_AMPL_WIDTH - 1),
		4780 => to_unsigned(14496, LUT_AMPL_WIDTH - 1),
		4781 => to_unsigned(14499, LUT_AMPL_WIDTH - 1),
		4782 => to_unsigned(14502, LUT_AMPL_WIDTH - 1),
		4783 => to_unsigned(14505, LUT_AMPL_WIDTH - 1),
		4784 => to_unsigned(14507, LUT_AMPL_WIDTH - 1),
		4785 => to_unsigned(14510, LUT_AMPL_WIDTH - 1),
		4786 => to_unsigned(14513, LUT_AMPL_WIDTH - 1),
		4787 => to_unsigned(14516, LUT_AMPL_WIDTH - 1),
		4788 => to_unsigned(14519, LUT_AMPL_WIDTH - 1),
		4789 => to_unsigned(14522, LUT_AMPL_WIDTH - 1),
		4790 => to_unsigned(14524, LUT_AMPL_WIDTH - 1),
		4791 => to_unsigned(14527, LUT_AMPL_WIDTH - 1),
		4792 => to_unsigned(14530, LUT_AMPL_WIDTH - 1),
		4793 => to_unsigned(14533, LUT_AMPL_WIDTH - 1),
		4794 => to_unsigned(14536, LUT_AMPL_WIDTH - 1),
		4795 => to_unsigned(14538, LUT_AMPL_WIDTH - 1),
		4796 => to_unsigned(14541, LUT_AMPL_WIDTH - 1),
		4797 => to_unsigned(14544, LUT_AMPL_WIDTH - 1),
		4798 => to_unsigned(14547, LUT_AMPL_WIDTH - 1),
		4799 => to_unsigned(14550, LUT_AMPL_WIDTH - 1),
		4800 => to_unsigned(14553, LUT_AMPL_WIDTH - 1),
		4801 => to_unsigned(14555, LUT_AMPL_WIDTH - 1),
		4802 => to_unsigned(14558, LUT_AMPL_WIDTH - 1),
		4803 => to_unsigned(14561, LUT_AMPL_WIDTH - 1),
		4804 => to_unsigned(14564, LUT_AMPL_WIDTH - 1),
		4805 => to_unsigned(14567, LUT_AMPL_WIDTH - 1),
		4806 => to_unsigned(14569, LUT_AMPL_WIDTH - 1),
		4807 => to_unsigned(14572, LUT_AMPL_WIDTH - 1),
		4808 => to_unsigned(14575, LUT_AMPL_WIDTH - 1),
		4809 => to_unsigned(14578, LUT_AMPL_WIDTH - 1),
		4810 => to_unsigned(14581, LUT_AMPL_WIDTH - 1),
		4811 => to_unsigned(14584, LUT_AMPL_WIDTH - 1),
		4812 => to_unsigned(14586, LUT_AMPL_WIDTH - 1),
		4813 => to_unsigned(14589, LUT_AMPL_WIDTH - 1),
		4814 => to_unsigned(14592, LUT_AMPL_WIDTH - 1),
		4815 => to_unsigned(14595, LUT_AMPL_WIDTH - 1),
		4816 => to_unsigned(14598, LUT_AMPL_WIDTH - 1),
		4817 => to_unsigned(14600, LUT_AMPL_WIDTH - 1),
		4818 => to_unsigned(14603, LUT_AMPL_WIDTH - 1),
		4819 => to_unsigned(14606, LUT_AMPL_WIDTH - 1),
		4820 => to_unsigned(14609, LUT_AMPL_WIDTH - 1),
		4821 => to_unsigned(14612, LUT_AMPL_WIDTH - 1),
		4822 => to_unsigned(14614, LUT_AMPL_WIDTH - 1),
		4823 => to_unsigned(14617, LUT_AMPL_WIDTH - 1),
		4824 => to_unsigned(14620, LUT_AMPL_WIDTH - 1),
		4825 => to_unsigned(14623, LUT_AMPL_WIDTH - 1),
		4826 => to_unsigned(14626, LUT_AMPL_WIDTH - 1),
		4827 => to_unsigned(14628, LUT_AMPL_WIDTH - 1),
		4828 => to_unsigned(14631, LUT_AMPL_WIDTH - 1),
		4829 => to_unsigned(14634, LUT_AMPL_WIDTH - 1),
		4830 => to_unsigned(14637, LUT_AMPL_WIDTH - 1),
		4831 => to_unsigned(14640, LUT_AMPL_WIDTH - 1),
		4832 => to_unsigned(14643, LUT_AMPL_WIDTH - 1),
		4833 => to_unsigned(14645, LUT_AMPL_WIDTH - 1),
		4834 => to_unsigned(14648, LUT_AMPL_WIDTH - 1),
		4835 => to_unsigned(14651, LUT_AMPL_WIDTH - 1),
		4836 => to_unsigned(14654, LUT_AMPL_WIDTH - 1),
		4837 => to_unsigned(14657, LUT_AMPL_WIDTH - 1),
		4838 => to_unsigned(14659, LUT_AMPL_WIDTH - 1),
		4839 => to_unsigned(14662, LUT_AMPL_WIDTH - 1),
		4840 => to_unsigned(14665, LUT_AMPL_WIDTH - 1),
		4841 => to_unsigned(14668, LUT_AMPL_WIDTH - 1),
		4842 => to_unsigned(14671, LUT_AMPL_WIDTH - 1),
		4843 => to_unsigned(14673, LUT_AMPL_WIDTH - 1),
		4844 => to_unsigned(14676, LUT_AMPL_WIDTH - 1),
		4845 => to_unsigned(14679, LUT_AMPL_WIDTH - 1),
		4846 => to_unsigned(14682, LUT_AMPL_WIDTH - 1),
		4847 => to_unsigned(14685, LUT_AMPL_WIDTH - 1),
		4848 => to_unsigned(14688, LUT_AMPL_WIDTH - 1),
		4849 => to_unsigned(14690, LUT_AMPL_WIDTH - 1),
		4850 => to_unsigned(14693, LUT_AMPL_WIDTH - 1),
		4851 => to_unsigned(14696, LUT_AMPL_WIDTH - 1),
		4852 => to_unsigned(14699, LUT_AMPL_WIDTH - 1),
		4853 => to_unsigned(14702, LUT_AMPL_WIDTH - 1),
		4854 => to_unsigned(14704, LUT_AMPL_WIDTH - 1),
		4855 => to_unsigned(14707, LUT_AMPL_WIDTH - 1),
		4856 => to_unsigned(14710, LUT_AMPL_WIDTH - 1),
		4857 => to_unsigned(14713, LUT_AMPL_WIDTH - 1),
		4858 => to_unsigned(14716, LUT_AMPL_WIDTH - 1),
		4859 => to_unsigned(14718, LUT_AMPL_WIDTH - 1),
		4860 => to_unsigned(14721, LUT_AMPL_WIDTH - 1),
		4861 => to_unsigned(14724, LUT_AMPL_WIDTH - 1),
		4862 => to_unsigned(14727, LUT_AMPL_WIDTH - 1),
		4863 => to_unsigned(14730, LUT_AMPL_WIDTH - 1),
		4864 => to_unsigned(14732, LUT_AMPL_WIDTH - 1),
		4865 => to_unsigned(14735, LUT_AMPL_WIDTH - 1),
		4866 => to_unsigned(14738, LUT_AMPL_WIDTH - 1),
		4867 => to_unsigned(14741, LUT_AMPL_WIDTH - 1),
		4868 => to_unsigned(14744, LUT_AMPL_WIDTH - 1),
		4869 => to_unsigned(14746, LUT_AMPL_WIDTH - 1),
		4870 => to_unsigned(14749, LUT_AMPL_WIDTH - 1),
		4871 => to_unsigned(14752, LUT_AMPL_WIDTH - 1),
		4872 => to_unsigned(14755, LUT_AMPL_WIDTH - 1),
		4873 => to_unsigned(14758, LUT_AMPL_WIDTH - 1),
		4874 => to_unsigned(14760, LUT_AMPL_WIDTH - 1),
		4875 => to_unsigned(14763, LUT_AMPL_WIDTH - 1),
		4876 => to_unsigned(14766, LUT_AMPL_WIDTH - 1),
		4877 => to_unsigned(14769, LUT_AMPL_WIDTH - 1),
		4878 => to_unsigned(14772, LUT_AMPL_WIDTH - 1),
		4879 => to_unsigned(14774, LUT_AMPL_WIDTH - 1),
		4880 => to_unsigned(14777, LUT_AMPL_WIDTH - 1),
		4881 => to_unsigned(14780, LUT_AMPL_WIDTH - 1),
		4882 => to_unsigned(14783, LUT_AMPL_WIDTH - 1),
		4883 => to_unsigned(14786, LUT_AMPL_WIDTH - 1),
		4884 => to_unsigned(14789, LUT_AMPL_WIDTH - 1),
		4885 => to_unsigned(14791, LUT_AMPL_WIDTH - 1),
		4886 => to_unsigned(14794, LUT_AMPL_WIDTH - 1),
		4887 => to_unsigned(14797, LUT_AMPL_WIDTH - 1),
		4888 => to_unsigned(14800, LUT_AMPL_WIDTH - 1),
		4889 => to_unsigned(14803, LUT_AMPL_WIDTH - 1),
		4890 => to_unsigned(14805, LUT_AMPL_WIDTH - 1),
		4891 => to_unsigned(14808, LUT_AMPL_WIDTH - 1),
		4892 => to_unsigned(14811, LUT_AMPL_WIDTH - 1),
		4893 => to_unsigned(14814, LUT_AMPL_WIDTH - 1),
		4894 => to_unsigned(14817, LUT_AMPL_WIDTH - 1),
		4895 => to_unsigned(14819, LUT_AMPL_WIDTH - 1),
		4896 => to_unsigned(14822, LUT_AMPL_WIDTH - 1),
		4897 => to_unsigned(14825, LUT_AMPL_WIDTH - 1),
		4898 => to_unsigned(14828, LUT_AMPL_WIDTH - 1),
		4899 => to_unsigned(14831, LUT_AMPL_WIDTH - 1),
		4900 => to_unsigned(14833, LUT_AMPL_WIDTH - 1),
		4901 => to_unsigned(14836, LUT_AMPL_WIDTH - 1),
		4902 => to_unsigned(14839, LUT_AMPL_WIDTH - 1),
		4903 => to_unsigned(14842, LUT_AMPL_WIDTH - 1),
		4904 => to_unsigned(14845, LUT_AMPL_WIDTH - 1),
		4905 => to_unsigned(14847, LUT_AMPL_WIDTH - 1),
		4906 => to_unsigned(14850, LUT_AMPL_WIDTH - 1),
		4907 => to_unsigned(14853, LUT_AMPL_WIDTH - 1),
		4908 => to_unsigned(14856, LUT_AMPL_WIDTH - 1),
		4909 => to_unsigned(14859, LUT_AMPL_WIDTH - 1),
		4910 => to_unsigned(14861, LUT_AMPL_WIDTH - 1),
		4911 => to_unsigned(14864, LUT_AMPL_WIDTH - 1),
		4912 => to_unsigned(14867, LUT_AMPL_WIDTH - 1),
		4913 => to_unsigned(14870, LUT_AMPL_WIDTH - 1),
		4914 => to_unsigned(14873, LUT_AMPL_WIDTH - 1),
		4915 => to_unsigned(14875, LUT_AMPL_WIDTH - 1),
		4916 => to_unsigned(14878, LUT_AMPL_WIDTH - 1),
		4917 => to_unsigned(14881, LUT_AMPL_WIDTH - 1),
		4918 => to_unsigned(14884, LUT_AMPL_WIDTH - 1),
		4919 => to_unsigned(14887, LUT_AMPL_WIDTH - 1),
		4920 => to_unsigned(14889, LUT_AMPL_WIDTH - 1),
		4921 => to_unsigned(14892, LUT_AMPL_WIDTH - 1),
		4922 => to_unsigned(14895, LUT_AMPL_WIDTH - 1),
		4923 => to_unsigned(14898, LUT_AMPL_WIDTH - 1),
		4924 => to_unsigned(14901, LUT_AMPL_WIDTH - 1),
		4925 => to_unsigned(14903, LUT_AMPL_WIDTH - 1),
		4926 => to_unsigned(14906, LUT_AMPL_WIDTH - 1),
		4927 => to_unsigned(14909, LUT_AMPL_WIDTH - 1),
		4928 => to_unsigned(14912, LUT_AMPL_WIDTH - 1),
		4929 => to_unsigned(14915, LUT_AMPL_WIDTH - 1),
		4930 => to_unsigned(14917, LUT_AMPL_WIDTH - 1),
		4931 => to_unsigned(14920, LUT_AMPL_WIDTH - 1),
		4932 => to_unsigned(14923, LUT_AMPL_WIDTH - 1),
		4933 => to_unsigned(14926, LUT_AMPL_WIDTH - 1),
		4934 => to_unsigned(14929, LUT_AMPL_WIDTH - 1),
		4935 => to_unsigned(14931, LUT_AMPL_WIDTH - 1),
		4936 => to_unsigned(14934, LUT_AMPL_WIDTH - 1),
		4937 => to_unsigned(14937, LUT_AMPL_WIDTH - 1),
		4938 => to_unsigned(14940, LUT_AMPL_WIDTH - 1),
		4939 => to_unsigned(14942, LUT_AMPL_WIDTH - 1),
		4940 => to_unsigned(14945, LUT_AMPL_WIDTH - 1),
		4941 => to_unsigned(14948, LUT_AMPL_WIDTH - 1),
		4942 => to_unsigned(14951, LUT_AMPL_WIDTH - 1),
		4943 => to_unsigned(14954, LUT_AMPL_WIDTH - 1),
		4944 => to_unsigned(14956, LUT_AMPL_WIDTH - 1),
		4945 => to_unsigned(14959, LUT_AMPL_WIDTH - 1),
		4946 => to_unsigned(14962, LUT_AMPL_WIDTH - 1),
		4947 => to_unsigned(14965, LUT_AMPL_WIDTH - 1),
		4948 => to_unsigned(14968, LUT_AMPL_WIDTH - 1),
		4949 => to_unsigned(14970, LUT_AMPL_WIDTH - 1),
		4950 => to_unsigned(14973, LUT_AMPL_WIDTH - 1),
		4951 => to_unsigned(14976, LUT_AMPL_WIDTH - 1),
		4952 => to_unsigned(14979, LUT_AMPL_WIDTH - 1),
		4953 => to_unsigned(14982, LUT_AMPL_WIDTH - 1),
		4954 => to_unsigned(14984, LUT_AMPL_WIDTH - 1),
		4955 => to_unsigned(14987, LUT_AMPL_WIDTH - 1),
		4956 => to_unsigned(14990, LUT_AMPL_WIDTH - 1),
		4957 => to_unsigned(14993, LUT_AMPL_WIDTH - 1),
		4958 => to_unsigned(14996, LUT_AMPL_WIDTH - 1),
		4959 => to_unsigned(14998, LUT_AMPL_WIDTH - 1),
		4960 => to_unsigned(15001, LUT_AMPL_WIDTH - 1),
		4961 => to_unsigned(15004, LUT_AMPL_WIDTH - 1),
		4962 => to_unsigned(15007, LUT_AMPL_WIDTH - 1),
		4963 => to_unsigned(15010, LUT_AMPL_WIDTH - 1),
		4964 => to_unsigned(15012, LUT_AMPL_WIDTH - 1),
		4965 => to_unsigned(15015, LUT_AMPL_WIDTH - 1),
		4966 => to_unsigned(15018, LUT_AMPL_WIDTH - 1),
		4967 => to_unsigned(15021, LUT_AMPL_WIDTH - 1),
		4968 => to_unsigned(15024, LUT_AMPL_WIDTH - 1),
		4969 => to_unsigned(15026, LUT_AMPL_WIDTH - 1),
		4970 => to_unsigned(15029, LUT_AMPL_WIDTH - 1),
		4971 => to_unsigned(15032, LUT_AMPL_WIDTH - 1),
		4972 => to_unsigned(15035, LUT_AMPL_WIDTH - 1),
		4973 => to_unsigned(15037, LUT_AMPL_WIDTH - 1),
		4974 => to_unsigned(15040, LUT_AMPL_WIDTH - 1),
		4975 => to_unsigned(15043, LUT_AMPL_WIDTH - 1),
		4976 => to_unsigned(15046, LUT_AMPL_WIDTH - 1),
		4977 => to_unsigned(15049, LUT_AMPL_WIDTH - 1),
		4978 => to_unsigned(15051, LUT_AMPL_WIDTH - 1),
		4979 => to_unsigned(15054, LUT_AMPL_WIDTH - 1),
		4980 => to_unsigned(15057, LUT_AMPL_WIDTH - 1),
		4981 => to_unsigned(15060, LUT_AMPL_WIDTH - 1),
		4982 => to_unsigned(15063, LUT_AMPL_WIDTH - 1),
		4983 => to_unsigned(15065, LUT_AMPL_WIDTH - 1),
		4984 => to_unsigned(15068, LUT_AMPL_WIDTH - 1),
		4985 => to_unsigned(15071, LUT_AMPL_WIDTH - 1),
		4986 => to_unsigned(15074, LUT_AMPL_WIDTH - 1),
		4987 => to_unsigned(15077, LUT_AMPL_WIDTH - 1),
		4988 => to_unsigned(15079, LUT_AMPL_WIDTH - 1),
		4989 => to_unsigned(15082, LUT_AMPL_WIDTH - 1),
		4990 => to_unsigned(15085, LUT_AMPL_WIDTH - 1),
		4991 => to_unsigned(15088, LUT_AMPL_WIDTH - 1),
		4992 => to_unsigned(15090, LUT_AMPL_WIDTH - 1),
		4993 => to_unsigned(15093, LUT_AMPL_WIDTH - 1),
		4994 => to_unsigned(15096, LUT_AMPL_WIDTH - 1),
		4995 => to_unsigned(15099, LUT_AMPL_WIDTH - 1),
		4996 => to_unsigned(15102, LUT_AMPL_WIDTH - 1),
		4997 => to_unsigned(15104, LUT_AMPL_WIDTH - 1),
		4998 => to_unsigned(15107, LUT_AMPL_WIDTH - 1),
		4999 => to_unsigned(15110, LUT_AMPL_WIDTH - 1),
		5000 => to_unsigned(15113, LUT_AMPL_WIDTH - 1),
		5001 => to_unsigned(15116, LUT_AMPL_WIDTH - 1),
		5002 => to_unsigned(15118, LUT_AMPL_WIDTH - 1),
		5003 => to_unsigned(15121, LUT_AMPL_WIDTH - 1),
		5004 => to_unsigned(15124, LUT_AMPL_WIDTH - 1),
		5005 => to_unsigned(15127, LUT_AMPL_WIDTH - 1),
		5006 => to_unsigned(15129, LUT_AMPL_WIDTH - 1),
		5007 => to_unsigned(15132, LUT_AMPL_WIDTH - 1),
		5008 => to_unsigned(15135, LUT_AMPL_WIDTH - 1),
		5009 => to_unsigned(15138, LUT_AMPL_WIDTH - 1),
		5010 => to_unsigned(15141, LUT_AMPL_WIDTH - 1),
		5011 => to_unsigned(15143, LUT_AMPL_WIDTH - 1),
		5012 => to_unsigned(15146, LUT_AMPL_WIDTH - 1),
		5013 => to_unsigned(15149, LUT_AMPL_WIDTH - 1),
		5014 => to_unsigned(15152, LUT_AMPL_WIDTH - 1),
		5015 => to_unsigned(15155, LUT_AMPL_WIDTH - 1),
		5016 => to_unsigned(15157, LUT_AMPL_WIDTH - 1),
		5017 => to_unsigned(15160, LUT_AMPL_WIDTH - 1),
		5018 => to_unsigned(15163, LUT_AMPL_WIDTH - 1),
		5019 => to_unsigned(15166, LUT_AMPL_WIDTH - 1),
		5020 => to_unsigned(15168, LUT_AMPL_WIDTH - 1),
		5021 => to_unsigned(15171, LUT_AMPL_WIDTH - 1),
		5022 => to_unsigned(15174, LUT_AMPL_WIDTH - 1),
		5023 => to_unsigned(15177, LUT_AMPL_WIDTH - 1),
		5024 => to_unsigned(15180, LUT_AMPL_WIDTH - 1),
		5025 => to_unsigned(15182, LUT_AMPL_WIDTH - 1),
		5026 => to_unsigned(15185, LUT_AMPL_WIDTH - 1),
		5027 => to_unsigned(15188, LUT_AMPL_WIDTH - 1),
		5028 => to_unsigned(15191, LUT_AMPL_WIDTH - 1),
		5029 => to_unsigned(15194, LUT_AMPL_WIDTH - 1),
		5030 => to_unsigned(15196, LUT_AMPL_WIDTH - 1),
		5031 => to_unsigned(15199, LUT_AMPL_WIDTH - 1),
		5032 => to_unsigned(15202, LUT_AMPL_WIDTH - 1),
		5033 => to_unsigned(15205, LUT_AMPL_WIDTH - 1),
		5034 => to_unsigned(15207, LUT_AMPL_WIDTH - 1),
		5035 => to_unsigned(15210, LUT_AMPL_WIDTH - 1),
		5036 => to_unsigned(15213, LUT_AMPL_WIDTH - 1),
		5037 => to_unsigned(15216, LUT_AMPL_WIDTH - 1),
		5038 => to_unsigned(15219, LUT_AMPL_WIDTH - 1),
		5039 => to_unsigned(15221, LUT_AMPL_WIDTH - 1),
		5040 => to_unsigned(15224, LUT_AMPL_WIDTH - 1),
		5041 => to_unsigned(15227, LUT_AMPL_WIDTH - 1),
		5042 => to_unsigned(15230, LUT_AMPL_WIDTH - 1),
		5043 => to_unsigned(15233, LUT_AMPL_WIDTH - 1),
		5044 => to_unsigned(15235, LUT_AMPL_WIDTH - 1),
		5045 => to_unsigned(15238, LUT_AMPL_WIDTH - 1),
		5046 => to_unsigned(15241, LUT_AMPL_WIDTH - 1),
		5047 => to_unsigned(15244, LUT_AMPL_WIDTH - 1),
		5048 => to_unsigned(15246, LUT_AMPL_WIDTH - 1),
		5049 => to_unsigned(15249, LUT_AMPL_WIDTH - 1),
		5050 => to_unsigned(15252, LUT_AMPL_WIDTH - 1),
		5051 => to_unsigned(15255, LUT_AMPL_WIDTH - 1),
		5052 => to_unsigned(15258, LUT_AMPL_WIDTH - 1),
		5053 => to_unsigned(15260, LUT_AMPL_WIDTH - 1),
		5054 => to_unsigned(15263, LUT_AMPL_WIDTH - 1),
		5055 => to_unsigned(15266, LUT_AMPL_WIDTH - 1),
		5056 => to_unsigned(15269, LUT_AMPL_WIDTH - 1),
		5057 => to_unsigned(15271, LUT_AMPL_WIDTH - 1),
		5058 => to_unsigned(15274, LUT_AMPL_WIDTH - 1),
		5059 => to_unsigned(15277, LUT_AMPL_WIDTH - 1),
		5060 => to_unsigned(15280, LUT_AMPL_WIDTH - 1),
		5061 => to_unsigned(15283, LUT_AMPL_WIDTH - 1),
		5062 => to_unsigned(15285, LUT_AMPL_WIDTH - 1),
		5063 => to_unsigned(15288, LUT_AMPL_WIDTH - 1),
		5064 => to_unsigned(15291, LUT_AMPL_WIDTH - 1),
		5065 => to_unsigned(15294, LUT_AMPL_WIDTH - 1),
		5066 => to_unsigned(15296, LUT_AMPL_WIDTH - 1),
		5067 => to_unsigned(15299, LUT_AMPL_WIDTH - 1),
		5068 => to_unsigned(15302, LUT_AMPL_WIDTH - 1),
		5069 => to_unsigned(15305, LUT_AMPL_WIDTH - 1),
		5070 => to_unsigned(15308, LUT_AMPL_WIDTH - 1),
		5071 => to_unsigned(15310, LUT_AMPL_WIDTH - 1),
		5072 => to_unsigned(15313, LUT_AMPL_WIDTH - 1),
		5073 => to_unsigned(15316, LUT_AMPL_WIDTH - 1),
		5074 => to_unsigned(15319, LUT_AMPL_WIDTH - 1),
		5075 => to_unsigned(15321, LUT_AMPL_WIDTH - 1),
		5076 => to_unsigned(15324, LUT_AMPL_WIDTH - 1),
		5077 => to_unsigned(15327, LUT_AMPL_WIDTH - 1),
		5078 => to_unsigned(15330, LUT_AMPL_WIDTH - 1),
		5079 => to_unsigned(15333, LUT_AMPL_WIDTH - 1),
		5080 => to_unsigned(15335, LUT_AMPL_WIDTH - 1),
		5081 => to_unsigned(15338, LUT_AMPL_WIDTH - 1),
		5082 => to_unsigned(15341, LUT_AMPL_WIDTH - 1),
		5083 => to_unsigned(15344, LUT_AMPL_WIDTH - 1),
		5084 => to_unsigned(15346, LUT_AMPL_WIDTH - 1),
		5085 => to_unsigned(15349, LUT_AMPL_WIDTH - 1),
		5086 => to_unsigned(15352, LUT_AMPL_WIDTH - 1),
		5087 => to_unsigned(15355, LUT_AMPL_WIDTH - 1),
		5088 => to_unsigned(15358, LUT_AMPL_WIDTH - 1),
		5089 => to_unsigned(15360, LUT_AMPL_WIDTH - 1),
		5090 => to_unsigned(15363, LUT_AMPL_WIDTH - 1),
		5091 => to_unsigned(15366, LUT_AMPL_WIDTH - 1),
		5092 => to_unsigned(15369, LUT_AMPL_WIDTH - 1),
		5093 => to_unsigned(15371, LUT_AMPL_WIDTH - 1),
		5094 => to_unsigned(15374, LUT_AMPL_WIDTH - 1),
		5095 => to_unsigned(15377, LUT_AMPL_WIDTH - 1),
		5096 => to_unsigned(15380, LUT_AMPL_WIDTH - 1),
		5097 => to_unsigned(15382, LUT_AMPL_WIDTH - 1),
		5098 => to_unsigned(15385, LUT_AMPL_WIDTH - 1),
		5099 => to_unsigned(15388, LUT_AMPL_WIDTH - 1),
		5100 => to_unsigned(15391, LUT_AMPL_WIDTH - 1),
		5101 => to_unsigned(15394, LUT_AMPL_WIDTH - 1),
		5102 => to_unsigned(15396, LUT_AMPL_WIDTH - 1),
		5103 => to_unsigned(15399, LUT_AMPL_WIDTH - 1),
		5104 => to_unsigned(15402, LUT_AMPL_WIDTH - 1),
		5105 => to_unsigned(15405, LUT_AMPL_WIDTH - 1),
		5106 => to_unsigned(15407, LUT_AMPL_WIDTH - 1),
		5107 => to_unsigned(15410, LUT_AMPL_WIDTH - 1),
		5108 => to_unsigned(15413, LUT_AMPL_WIDTH - 1),
		5109 => to_unsigned(15416, LUT_AMPL_WIDTH - 1),
		5110 => to_unsigned(15419, LUT_AMPL_WIDTH - 1),
		5111 => to_unsigned(15421, LUT_AMPL_WIDTH - 1),
		5112 => to_unsigned(15424, LUT_AMPL_WIDTH - 1),
		5113 => to_unsigned(15427, LUT_AMPL_WIDTH - 1),
		5114 => to_unsigned(15430, LUT_AMPL_WIDTH - 1),
		5115 => to_unsigned(15432, LUT_AMPL_WIDTH - 1),
		5116 => to_unsigned(15435, LUT_AMPL_WIDTH - 1),
		5117 => to_unsigned(15438, LUT_AMPL_WIDTH - 1),
		5118 => to_unsigned(15441, LUT_AMPL_WIDTH - 1),
		5119 => to_unsigned(15443, LUT_AMPL_WIDTH - 1),
		5120 => to_unsigned(15446, LUT_AMPL_WIDTH - 1),
		5121 => to_unsigned(15449, LUT_AMPL_WIDTH - 1),
		5122 => to_unsigned(15452, LUT_AMPL_WIDTH - 1),
		5123 => to_unsigned(15455, LUT_AMPL_WIDTH - 1),
		5124 => to_unsigned(15457, LUT_AMPL_WIDTH - 1),
		5125 => to_unsigned(15460, LUT_AMPL_WIDTH - 1),
		5126 => to_unsigned(15463, LUT_AMPL_WIDTH - 1),
		5127 => to_unsigned(15466, LUT_AMPL_WIDTH - 1),
		5128 => to_unsigned(15468, LUT_AMPL_WIDTH - 1),
		5129 => to_unsigned(15471, LUT_AMPL_WIDTH - 1),
		5130 => to_unsigned(15474, LUT_AMPL_WIDTH - 1),
		5131 => to_unsigned(15477, LUT_AMPL_WIDTH - 1),
		5132 => to_unsigned(15479, LUT_AMPL_WIDTH - 1),
		5133 => to_unsigned(15482, LUT_AMPL_WIDTH - 1),
		5134 => to_unsigned(15485, LUT_AMPL_WIDTH - 1),
		5135 => to_unsigned(15488, LUT_AMPL_WIDTH - 1),
		5136 => to_unsigned(15491, LUT_AMPL_WIDTH - 1),
		5137 => to_unsigned(15493, LUT_AMPL_WIDTH - 1),
		5138 => to_unsigned(15496, LUT_AMPL_WIDTH - 1),
		5139 => to_unsigned(15499, LUT_AMPL_WIDTH - 1),
		5140 => to_unsigned(15502, LUT_AMPL_WIDTH - 1),
		5141 => to_unsigned(15504, LUT_AMPL_WIDTH - 1),
		5142 => to_unsigned(15507, LUT_AMPL_WIDTH - 1),
		5143 => to_unsigned(15510, LUT_AMPL_WIDTH - 1),
		5144 => to_unsigned(15513, LUT_AMPL_WIDTH - 1),
		5145 => to_unsigned(15515, LUT_AMPL_WIDTH - 1),
		5146 => to_unsigned(15518, LUT_AMPL_WIDTH - 1),
		5147 => to_unsigned(15521, LUT_AMPL_WIDTH - 1),
		5148 => to_unsigned(15524, LUT_AMPL_WIDTH - 1),
		5149 => to_unsigned(15527, LUT_AMPL_WIDTH - 1),
		5150 => to_unsigned(15529, LUT_AMPL_WIDTH - 1),
		5151 => to_unsigned(15532, LUT_AMPL_WIDTH - 1),
		5152 => to_unsigned(15535, LUT_AMPL_WIDTH - 1),
		5153 => to_unsigned(15538, LUT_AMPL_WIDTH - 1),
		5154 => to_unsigned(15540, LUT_AMPL_WIDTH - 1),
		5155 => to_unsigned(15543, LUT_AMPL_WIDTH - 1),
		5156 => to_unsigned(15546, LUT_AMPL_WIDTH - 1),
		5157 => to_unsigned(15549, LUT_AMPL_WIDTH - 1),
		5158 => to_unsigned(15551, LUT_AMPL_WIDTH - 1),
		5159 => to_unsigned(15554, LUT_AMPL_WIDTH - 1),
		5160 => to_unsigned(15557, LUT_AMPL_WIDTH - 1),
		5161 => to_unsigned(15560, LUT_AMPL_WIDTH - 1),
		5162 => to_unsigned(15562, LUT_AMPL_WIDTH - 1),
		5163 => to_unsigned(15565, LUT_AMPL_WIDTH - 1),
		5164 => to_unsigned(15568, LUT_AMPL_WIDTH - 1),
		5165 => to_unsigned(15571, LUT_AMPL_WIDTH - 1),
		5166 => to_unsigned(15574, LUT_AMPL_WIDTH - 1),
		5167 => to_unsigned(15576, LUT_AMPL_WIDTH - 1),
		5168 => to_unsigned(15579, LUT_AMPL_WIDTH - 1),
		5169 => to_unsigned(15582, LUT_AMPL_WIDTH - 1),
		5170 => to_unsigned(15585, LUT_AMPL_WIDTH - 1),
		5171 => to_unsigned(15587, LUT_AMPL_WIDTH - 1),
		5172 => to_unsigned(15590, LUT_AMPL_WIDTH - 1),
		5173 => to_unsigned(15593, LUT_AMPL_WIDTH - 1),
		5174 => to_unsigned(15596, LUT_AMPL_WIDTH - 1),
		5175 => to_unsigned(15598, LUT_AMPL_WIDTH - 1),
		5176 => to_unsigned(15601, LUT_AMPL_WIDTH - 1),
		5177 => to_unsigned(15604, LUT_AMPL_WIDTH - 1),
		5178 => to_unsigned(15607, LUT_AMPL_WIDTH - 1),
		5179 => to_unsigned(15609, LUT_AMPL_WIDTH - 1),
		5180 => to_unsigned(15612, LUT_AMPL_WIDTH - 1),
		5181 => to_unsigned(15615, LUT_AMPL_WIDTH - 1),
		5182 => to_unsigned(15618, LUT_AMPL_WIDTH - 1),
		5183 => to_unsigned(15621, LUT_AMPL_WIDTH - 1),
		5184 => to_unsigned(15623, LUT_AMPL_WIDTH - 1),
		5185 => to_unsigned(15626, LUT_AMPL_WIDTH - 1),
		5186 => to_unsigned(15629, LUT_AMPL_WIDTH - 1),
		5187 => to_unsigned(15632, LUT_AMPL_WIDTH - 1),
		5188 => to_unsigned(15634, LUT_AMPL_WIDTH - 1),
		5189 => to_unsigned(15637, LUT_AMPL_WIDTH - 1),
		5190 => to_unsigned(15640, LUT_AMPL_WIDTH - 1),
		5191 => to_unsigned(15643, LUT_AMPL_WIDTH - 1),
		5192 => to_unsigned(15645, LUT_AMPL_WIDTH - 1),
		5193 => to_unsigned(15648, LUT_AMPL_WIDTH - 1),
		5194 => to_unsigned(15651, LUT_AMPL_WIDTH - 1),
		5195 => to_unsigned(15654, LUT_AMPL_WIDTH - 1),
		5196 => to_unsigned(15656, LUT_AMPL_WIDTH - 1),
		5197 => to_unsigned(15659, LUT_AMPL_WIDTH - 1),
		5198 => to_unsigned(15662, LUT_AMPL_WIDTH - 1),
		5199 => to_unsigned(15665, LUT_AMPL_WIDTH - 1),
		5200 => to_unsigned(15667, LUT_AMPL_WIDTH - 1),
		5201 => to_unsigned(15670, LUT_AMPL_WIDTH - 1),
		5202 => to_unsigned(15673, LUT_AMPL_WIDTH - 1),
		5203 => to_unsigned(15676, LUT_AMPL_WIDTH - 1),
		5204 => to_unsigned(15678, LUT_AMPL_WIDTH - 1),
		5205 => to_unsigned(15681, LUT_AMPL_WIDTH - 1),
		5206 => to_unsigned(15684, LUT_AMPL_WIDTH - 1),
		5207 => to_unsigned(15687, LUT_AMPL_WIDTH - 1),
		5208 => to_unsigned(15690, LUT_AMPL_WIDTH - 1),
		5209 => to_unsigned(15692, LUT_AMPL_WIDTH - 1),
		5210 => to_unsigned(15695, LUT_AMPL_WIDTH - 1),
		5211 => to_unsigned(15698, LUT_AMPL_WIDTH - 1),
		5212 => to_unsigned(15701, LUT_AMPL_WIDTH - 1),
		5213 => to_unsigned(15703, LUT_AMPL_WIDTH - 1),
		5214 => to_unsigned(15706, LUT_AMPL_WIDTH - 1),
		5215 => to_unsigned(15709, LUT_AMPL_WIDTH - 1),
		5216 => to_unsigned(15712, LUT_AMPL_WIDTH - 1),
		5217 => to_unsigned(15714, LUT_AMPL_WIDTH - 1),
		5218 => to_unsigned(15717, LUT_AMPL_WIDTH - 1),
		5219 => to_unsigned(15720, LUT_AMPL_WIDTH - 1),
		5220 => to_unsigned(15723, LUT_AMPL_WIDTH - 1),
		5221 => to_unsigned(15725, LUT_AMPL_WIDTH - 1),
		5222 => to_unsigned(15728, LUT_AMPL_WIDTH - 1),
		5223 => to_unsigned(15731, LUT_AMPL_WIDTH - 1),
		5224 => to_unsigned(15734, LUT_AMPL_WIDTH - 1),
		5225 => to_unsigned(15736, LUT_AMPL_WIDTH - 1),
		5226 => to_unsigned(15739, LUT_AMPL_WIDTH - 1),
		5227 => to_unsigned(15742, LUT_AMPL_WIDTH - 1),
		5228 => to_unsigned(15745, LUT_AMPL_WIDTH - 1),
		5229 => to_unsigned(15747, LUT_AMPL_WIDTH - 1),
		5230 => to_unsigned(15750, LUT_AMPL_WIDTH - 1),
		5231 => to_unsigned(15753, LUT_AMPL_WIDTH - 1),
		5232 => to_unsigned(15756, LUT_AMPL_WIDTH - 1),
		5233 => to_unsigned(15758, LUT_AMPL_WIDTH - 1),
		5234 => to_unsigned(15761, LUT_AMPL_WIDTH - 1),
		5235 => to_unsigned(15764, LUT_AMPL_WIDTH - 1),
		5236 => to_unsigned(15767, LUT_AMPL_WIDTH - 1),
		5237 => to_unsigned(15769, LUT_AMPL_WIDTH - 1),
		5238 => to_unsigned(15772, LUT_AMPL_WIDTH - 1),
		5239 => to_unsigned(15775, LUT_AMPL_WIDTH - 1),
		5240 => to_unsigned(15778, LUT_AMPL_WIDTH - 1),
		5241 => to_unsigned(15780, LUT_AMPL_WIDTH - 1),
		5242 => to_unsigned(15783, LUT_AMPL_WIDTH - 1),
		5243 => to_unsigned(15786, LUT_AMPL_WIDTH - 1),
		5244 => to_unsigned(15789, LUT_AMPL_WIDTH - 1),
		5245 => to_unsigned(15791, LUT_AMPL_WIDTH - 1),
		5246 => to_unsigned(15794, LUT_AMPL_WIDTH - 1),
		5247 => to_unsigned(15797, LUT_AMPL_WIDTH - 1),
		5248 => to_unsigned(15800, LUT_AMPL_WIDTH - 1),
		5249 => to_unsigned(15802, LUT_AMPL_WIDTH - 1),
		5250 => to_unsigned(15805, LUT_AMPL_WIDTH - 1),
		5251 => to_unsigned(15808, LUT_AMPL_WIDTH - 1),
		5252 => to_unsigned(15811, LUT_AMPL_WIDTH - 1),
		5253 => to_unsigned(15813, LUT_AMPL_WIDTH - 1),
		5254 => to_unsigned(15816, LUT_AMPL_WIDTH - 1),
		5255 => to_unsigned(15819, LUT_AMPL_WIDTH - 1),
		5256 => to_unsigned(15822, LUT_AMPL_WIDTH - 1),
		5257 => to_unsigned(15824, LUT_AMPL_WIDTH - 1),
		5258 => to_unsigned(15827, LUT_AMPL_WIDTH - 1),
		5259 => to_unsigned(15830, LUT_AMPL_WIDTH - 1),
		5260 => to_unsigned(15833, LUT_AMPL_WIDTH - 1),
		5261 => to_unsigned(15835, LUT_AMPL_WIDTH - 1),
		5262 => to_unsigned(15838, LUT_AMPL_WIDTH - 1),
		5263 => to_unsigned(15841, LUT_AMPL_WIDTH - 1),
		5264 => to_unsigned(15844, LUT_AMPL_WIDTH - 1),
		5265 => to_unsigned(15846, LUT_AMPL_WIDTH - 1),
		5266 => to_unsigned(15849, LUT_AMPL_WIDTH - 1),
		5267 => to_unsigned(15852, LUT_AMPL_WIDTH - 1),
		5268 => to_unsigned(15855, LUT_AMPL_WIDTH - 1),
		5269 => to_unsigned(15857, LUT_AMPL_WIDTH - 1),
		5270 => to_unsigned(15860, LUT_AMPL_WIDTH - 1),
		5271 => to_unsigned(15863, LUT_AMPL_WIDTH - 1),
		5272 => to_unsigned(15866, LUT_AMPL_WIDTH - 1),
		5273 => to_unsigned(15868, LUT_AMPL_WIDTH - 1),
		5274 => to_unsigned(15871, LUT_AMPL_WIDTH - 1),
		5275 => to_unsigned(15874, LUT_AMPL_WIDTH - 1),
		5276 => to_unsigned(15877, LUT_AMPL_WIDTH - 1),
		5277 => to_unsigned(15879, LUT_AMPL_WIDTH - 1),
		5278 => to_unsigned(15882, LUT_AMPL_WIDTH - 1),
		5279 => to_unsigned(15885, LUT_AMPL_WIDTH - 1),
		5280 => to_unsigned(15888, LUT_AMPL_WIDTH - 1),
		5281 => to_unsigned(15890, LUT_AMPL_WIDTH - 1),
		5282 => to_unsigned(15893, LUT_AMPL_WIDTH - 1),
		5283 => to_unsigned(15896, LUT_AMPL_WIDTH - 1),
		5284 => to_unsigned(15899, LUT_AMPL_WIDTH - 1),
		5285 => to_unsigned(15901, LUT_AMPL_WIDTH - 1),
		5286 => to_unsigned(15904, LUT_AMPL_WIDTH - 1),
		5287 => to_unsigned(15907, LUT_AMPL_WIDTH - 1),
		5288 => to_unsigned(15910, LUT_AMPL_WIDTH - 1),
		5289 => to_unsigned(15912, LUT_AMPL_WIDTH - 1),
		5290 => to_unsigned(15915, LUT_AMPL_WIDTH - 1),
		5291 => to_unsigned(15918, LUT_AMPL_WIDTH - 1),
		5292 => to_unsigned(15921, LUT_AMPL_WIDTH - 1),
		5293 => to_unsigned(15923, LUT_AMPL_WIDTH - 1),
		5294 => to_unsigned(15926, LUT_AMPL_WIDTH - 1),
		5295 => to_unsigned(15929, LUT_AMPL_WIDTH - 1),
		5296 => to_unsigned(15932, LUT_AMPL_WIDTH - 1),
		5297 => to_unsigned(15934, LUT_AMPL_WIDTH - 1),
		5298 => to_unsigned(15937, LUT_AMPL_WIDTH - 1),
		5299 => to_unsigned(15940, LUT_AMPL_WIDTH - 1),
		5300 => to_unsigned(15943, LUT_AMPL_WIDTH - 1),
		5301 => to_unsigned(15945, LUT_AMPL_WIDTH - 1),
		5302 => to_unsigned(15948, LUT_AMPL_WIDTH - 1),
		5303 => to_unsigned(15951, LUT_AMPL_WIDTH - 1),
		5304 => to_unsigned(15954, LUT_AMPL_WIDTH - 1),
		5305 => to_unsigned(15956, LUT_AMPL_WIDTH - 1),
		5306 => to_unsigned(15959, LUT_AMPL_WIDTH - 1),
		5307 => to_unsigned(15962, LUT_AMPL_WIDTH - 1),
		5308 => to_unsigned(15965, LUT_AMPL_WIDTH - 1),
		5309 => to_unsigned(15967, LUT_AMPL_WIDTH - 1),
		5310 => to_unsigned(15970, LUT_AMPL_WIDTH - 1),
		5311 => to_unsigned(15973, LUT_AMPL_WIDTH - 1),
		5312 => to_unsigned(15976, LUT_AMPL_WIDTH - 1),
		5313 => to_unsigned(15978, LUT_AMPL_WIDTH - 1),
		5314 => to_unsigned(15981, LUT_AMPL_WIDTH - 1),
		5315 => to_unsigned(15984, LUT_AMPL_WIDTH - 1),
		5316 => to_unsigned(15987, LUT_AMPL_WIDTH - 1),
		5317 => to_unsigned(15989, LUT_AMPL_WIDTH - 1),
		5318 => to_unsigned(15992, LUT_AMPL_WIDTH - 1),
		5319 => to_unsigned(15995, LUT_AMPL_WIDTH - 1),
		5320 => to_unsigned(15997, LUT_AMPL_WIDTH - 1),
		5321 => to_unsigned(16000, LUT_AMPL_WIDTH - 1),
		5322 => to_unsigned(16003, LUT_AMPL_WIDTH - 1),
		5323 => to_unsigned(16006, LUT_AMPL_WIDTH - 1),
		5324 => to_unsigned(16008, LUT_AMPL_WIDTH - 1),
		5325 => to_unsigned(16011, LUT_AMPL_WIDTH - 1),
		5326 => to_unsigned(16014, LUT_AMPL_WIDTH - 1),
		5327 => to_unsigned(16017, LUT_AMPL_WIDTH - 1),
		5328 => to_unsigned(16019, LUT_AMPL_WIDTH - 1),
		5329 => to_unsigned(16022, LUT_AMPL_WIDTH - 1),
		5330 => to_unsigned(16025, LUT_AMPL_WIDTH - 1),
		5331 => to_unsigned(16028, LUT_AMPL_WIDTH - 1),
		5332 => to_unsigned(16030, LUT_AMPL_WIDTH - 1),
		5333 => to_unsigned(16033, LUT_AMPL_WIDTH - 1),
		5334 => to_unsigned(16036, LUT_AMPL_WIDTH - 1),
		5335 => to_unsigned(16039, LUT_AMPL_WIDTH - 1),
		5336 => to_unsigned(16041, LUT_AMPL_WIDTH - 1),
		5337 => to_unsigned(16044, LUT_AMPL_WIDTH - 1),
		5338 => to_unsigned(16047, LUT_AMPL_WIDTH - 1),
		5339 => to_unsigned(16050, LUT_AMPL_WIDTH - 1),
		5340 => to_unsigned(16052, LUT_AMPL_WIDTH - 1),
		5341 => to_unsigned(16055, LUT_AMPL_WIDTH - 1),
		5342 => to_unsigned(16058, LUT_AMPL_WIDTH - 1),
		5343 => to_unsigned(16061, LUT_AMPL_WIDTH - 1),
		5344 => to_unsigned(16063, LUT_AMPL_WIDTH - 1),
		5345 => to_unsigned(16066, LUT_AMPL_WIDTH - 1),
		5346 => to_unsigned(16069, LUT_AMPL_WIDTH - 1),
		5347 => to_unsigned(16071, LUT_AMPL_WIDTH - 1),
		5348 => to_unsigned(16074, LUT_AMPL_WIDTH - 1),
		5349 => to_unsigned(16077, LUT_AMPL_WIDTH - 1),
		5350 => to_unsigned(16080, LUT_AMPL_WIDTH - 1),
		5351 => to_unsigned(16082, LUT_AMPL_WIDTH - 1),
		5352 => to_unsigned(16085, LUT_AMPL_WIDTH - 1),
		5353 => to_unsigned(16088, LUT_AMPL_WIDTH - 1),
		5354 => to_unsigned(16091, LUT_AMPL_WIDTH - 1),
		5355 => to_unsigned(16093, LUT_AMPL_WIDTH - 1),
		5356 => to_unsigned(16096, LUT_AMPL_WIDTH - 1),
		5357 => to_unsigned(16099, LUT_AMPL_WIDTH - 1),
		5358 => to_unsigned(16102, LUT_AMPL_WIDTH - 1),
		5359 => to_unsigned(16104, LUT_AMPL_WIDTH - 1),
		5360 => to_unsigned(16107, LUT_AMPL_WIDTH - 1),
		5361 => to_unsigned(16110, LUT_AMPL_WIDTH - 1),
		5362 => to_unsigned(16113, LUT_AMPL_WIDTH - 1),
		5363 => to_unsigned(16115, LUT_AMPL_WIDTH - 1),
		5364 => to_unsigned(16118, LUT_AMPL_WIDTH - 1),
		5365 => to_unsigned(16121, LUT_AMPL_WIDTH - 1),
		5366 => to_unsigned(16123, LUT_AMPL_WIDTH - 1),
		5367 => to_unsigned(16126, LUT_AMPL_WIDTH - 1),
		5368 => to_unsigned(16129, LUT_AMPL_WIDTH - 1),
		5369 => to_unsigned(16132, LUT_AMPL_WIDTH - 1),
		5370 => to_unsigned(16134, LUT_AMPL_WIDTH - 1),
		5371 => to_unsigned(16137, LUT_AMPL_WIDTH - 1),
		5372 => to_unsigned(16140, LUT_AMPL_WIDTH - 1),
		5373 => to_unsigned(16143, LUT_AMPL_WIDTH - 1),
		5374 => to_unsigned(16145, LUT_AMPL_WIDTH - 1),
		5375 => to_unsigned(16148, LUT_AMPL_WIDTH - 1),
		5376 => to_unsigned(16151, LUT_AMPL_WIDTH - 1),
		5377 => to_unsigned(16154, LUT_AMPL_WIDTH - 1),
		5378 => to_unsigned(16156, LUT_AMPL_WIDTH - 1),
		5379 => to_unsigned(16159, LUT_AMPL_WIDTH - 1),
		5380 => to_unsigned(16162, LUT_AMPL_WIDTH - 1),
		5381 => to_unsigned(16164, LUT_AMPL_WIDTH - 1),
		5382 => to_unsigned(16167, LUT_AMPL_WIDTH - 1),
		5383 => to_unsigned(16170, LUT_AMPL_WIDTH - 1),
		5384 => to_unsigned(16173, LUT_AMPL_WIDTH - 1),
		5385 => to_unsigned(16175, LUT_AMPL_WIDTH - 1),
		5386 => to_unsigned(16178, LUT_AMPL_WIDTH - 1),
		5387 => to_unsigned(16181, LUT_AMPL_WIDTH - 1),
		5388 => to_unsigned(16184, LUT_AMPL_WIDTH - 1),
		5389 => to_unsigned(16186, LUT_AMPL_WIDTH - 1),
		5390 => to_unsigned(16189, LUT_AMPL_WIDTH - 1),
		5391 => to_unsigned(16192, LUT_AMPL_WIDTH - 1),
		5392 => to_unsigned(16195, LUT_AMPL_WIDTH - 1),
		5393 => to_unsigned(16197, LUT_AMPL_WIDTH - 1),
		5394 => to_unsigned(16200, LUT_AMPL_WIDTH - 1),
		5395 => to_unsigned(16203, LUT_AMPL_WIDTH - 1),
		5396 => to_unsigned(16205, LUT_AMPL_WIDTH - 1),
		5397 => to_unsigned(16208, LUT_AMPL_WIDTH - 1),
		5398 => to_unsigned(16211, LUT_AMPL_WIDTH - 1),
		5399 => to_unsigned(16214, LUT_AMPL_WIDTH - 1),
		5400 => to_unsigned(16216, LUT_AMPL_WIDTH - 1),
		5401 => to_unsigned(16219, LUT_AMPL_WIDTH - 1),
		5402 => to_unsigned(16222, LUT_AMPL_WIDTH - 1),
		5403 => to_unsigned(16225, LUT_AMPL_WIDTH - 1),
		5404 => to_unsigned(16227, LUT_AMPL_WIDTH - 1),
		5405 => to_unsigned(16230, LUT_AMPL_WIDTH - 1),
		5406 => to_unsigned(16233, LUT_AMPL_WIDTH - 1),
		5407 => to_unsigned(16235, LUT_AMPL_WIDTH - 1),
		5408 => to_unsigned(16238, LUT_AMPL_WIDTH - 1),
		5409 => to_unsigned(16241, LUT_AMPL_WIDTH - 1),
		5410 => to_unsigned(16244, LUT_AMPL_WIDTH - 1),
		5411 => to_unsigned(16246, LUT_AMPL_WIDTH - 1),
		5412 => to_unsigned(16249, LUT_AMPL_WIDTH - 1),
		5413 => to_unsigned(16252, LUT_AMPL_WIDTH - 1),
		5414 => to_unsigned(16255, LUT_AMPL_WIDTH - 1),
		5415 => to_unsigned(16257, LUT_AMPL_WIDTH - 1),
		5416 => to_unsigned(16260, LUT_AMPL_WIDTH - 1),
		5417 => to_unsigned(16263, LUT_AMPL_WIDTH - 1),
		5418 => to_unsigned(16265, LUT_AMPL_WIDTH - 1),
		5419 => to_unsigned(16268, LUT_AMPL_WIDTH - 1),
		5420 => to_unsigned(16271, LUT_AMPL_WIDTH - 1),
		5421 => to_unsigned(16274, LUT_AMPL_WIDTH - 1),
		5422 => to_unsigned(16276, LUT_AMPL_WIDTH - 1),
		5423 => to_unsigned(16279, LUT_AMPL_WIDTH - 1),
		5424 => to_unsigned(16282, LUT_AMPL_WIDTH - 1),
		5425 => to_unsigned(16285, LUT_AMPL_WIDTH - 1),
		5426 => to_unsigned(16287, LUT_AMPL_WIDTH - 1),
		5427 => to_unsigned(16290, LUT_AMPL_WIDTH - 1),
		5428 => to_unsigned(16293, LUT_AMPL_WIDTH - 1),
		5429 => to_unsigned(16295, LUT_AMPL_WIDTH - 1),
		5430 => to_unsigned(16298, LUT_AMPL_WIDTH - 1),
		5431 => to_unsigned(16301, LUT_AMPL_WIDTH - 1),
		5432 => to_unsigned(16304, LUT_AMPL_WIDTH - 1),
		5433 => to_unsigned(16306, LUT_AMPL_WIDTH - 1),
		5434 => to_unsigned(16309, LUT_AMPL_WIDTH - 1),
		5435 => to_unsigned(16312, LUT_AMPL_WIDTH - 1),
		5436 => to_unsigned(16315, LUT_AMPL_WIDTH - 1),
		5437 => to_unsigned(16317, LUT_AMPL_WIDTH - 1),
		5438 => to_unsigned(16320, LUT_AMPL_WIDTH - 1),
		5439 => to_unsigned(16323, LUT_AMPL_WIDTH - 1),
		5440 => to_unsigned(16325, LUT_AMPL_WIDTH - 1),
		5441 => to_unsigned(16328, LUT_AMPL_WIDTH - 1),
		5442 => to_unsigned(16331, LUT_AMPL_WIDTH - 1),
		5443 => to_unsigned(16334, LUT_AMPL_WIDTH - 1),
		5444 => to_unsigned(16336, LUT_AMPL_WIDTH - 1),
		5445 => to_unsigned(16339, LUT_AMPL_WIDTH - 1),
		5446 => to_unsigned(16342, LUT_AMPL_WIDTH - 1),
		5447 => to_unsigned(16344, LUT_AMPL_WIDTH - 1),
		5448 => to_unsigned(16347, LUT_AMPL_WIDTH - 1),
		5449 => to_unsigned(16350, LUT_AMPL_WIDTH - 1),
		5450 => to_unsigned(16353, LUT_AMPL_WIDTH - 1),
		5451 => to_unsigned(16355, LUT_AMPL_WIDTH - 1),
		5452 => to_unsigned(16358, LUT_AMPL_WIDTH - 1),
		5453 => to_unsigned(16361, LUT_AMPL_WIDTH - 1),
		5454 => to_unsigned(16364, LUT_AMPL_WIDTH - 1),
		5455 => to_unsigned(16366, LUT_AMPL_WIDTH - 1),
		5456 => to_unsigned(16369, LUT_AMPL_WIDTH - 1),
		5457 => to_unsigned(16372, LUT_AMPL_WIDTH - 1),
		5458 => to_unsigned(16374, LUT_AMPL_WIDTH - 1),
		5459 => to_unsigned(16377, LUT_AMPL_WIDTH - 1),
		5460 => to_unsigned(16380, LUT_AMPL_WIDTH - 1),
		5461 => to_unsigned(16383, LUT_AMPL_WIDTH - 1),
		5462 => to_unsigned(16385, LUT_AMPL_WIDTH - 1),
		5463 => to_unsigned(16388, LUT_AMPL_WIDTH - 1),
		5464 => to_unsigned(16391, LUT_AMPL_WIDTH - 1),
		5465 => to_unsigned(16393, LUT_AMPL_WIDTH - 1),
		5466 => to_unsigned(16396, LUT_AMPL_WIDTH - 1),
		5467 => to_unsigned(16399, LUT_AMPL_WIDTH - 1),
		5468 => to_unsigned(16402, LUT_AMPL_WIDTH - 1),
		5469 => to_unsigned(16404, LUT_AMPL_WIDTH - 1),
		5470 => to_unsigned(16407, LUT_AMPL_WIDTH - 1),
		5471 => to_unsigned(16410, LUT_AMPL_WIDTH - 1),
		5472 => to_unsigned(16413, LUT_AMPL_WIDTH - 1),
		5473 => to_unsigned(16415, LUT_AMPL_WIDTH - 1),
		5474 => to_unsigned(16418, LUT_AMPL_WIDTH - 1),
		5475 => to_unsigned(16421, LUT_AMPL_WIDTH - 1),
		5476 => to_unsigned(16423, LUT_AMPL_WIDTH - 1),
		5477 => to_unsigned(16426, LUT_AMPL_WIDTH - 1),
		5478 => to_unsigned(16429, LUT_AMPL_WIDTH - 1),
		5479 => to_unsigned(16432, LUT_AMPL_WIDTH - 1),
		5480 => to_unsigned(16434, LUT_AMPL_WIDTH - 1),
		5481 => to_unsigned(16437, LUT_AMPL_WIDTH - 1),
		5482 => to_unsigned(16440, LUT_AMPL_WIDTH - 1),
		5483 => to_unsigned(16442, LUT_AMPL_WIDTH - 1),
		5484 => to_unsigned(16445, LUT_AMPL_WIDTH - 1),
		5485 => to_unsigned(16448, LUT_AMPL_WIDTH - 1),
		5486 => to_unsigned(16451, LUT_AMPL_WIDTH - 1),
		5487 => to_unsigned(16453, LUT_AMPL_WIDTH - 1),
		5488 => to_unsigned(16456, LUT_AMPL_WIDTH - 1),
		5489 => to_unsigned(16459, LUT_AMPL_WIDTH - 1),
		5490 => to_unsigned(16461, LUT_AMPL_WIDTH - 1),
		5491 => to_unsigned(16464, LUT_AMPL_WIDTH - 1),
		5492 => to_unsigned(16467, LUT_AMPL_WIDTH - 1),
		5493 => to_unsigned(16470, LUT_AMPL_WIDTH - 1),
		5494 => to_unsigned(16472, LUT_AMPL_WIDTH - 1),
		5495 => to_unsigned(16475, LUT_AMPL_WIDTH - 1),
		5496 => to_unsigned(16478, LUT_AMPL_WIDTH - 1),
		5497 => to_unsigned(16480, LUT_AMPL_WIDTH - 1),
		5498 => to_unsigned(16483, LUT_AMPL_WIDTH - 1),
		5499 => to_unsigned(16486, LUT_AMPL_WIDTH - 1),
		5500 => to_unsigned(16489, LUT_AMPL_WIDTH - 1),
		5501 => to_unsigned(16491, LUT_AMPL_WIDTH - 1),
		5502 => to_unsigned(16494, LUT_AMPL_WIDTH - 1),
		5503 => to_unsigned(16497, LUT_AMPL_WIDTH - 1),
		5504 => to_unsigned(16499, LUT_AMPL_WIDTH - 1),
		5505 => to_unsigned(16502, LUT_AMPL_WIDTH - 1),
		5506 => to_unsigned(16505, LUT_AMPL_WIDTH - 1),
		5507 => to_unsigned(16508, LUT_AMPL_WIDTH - 1),
		5508 => to_unsigned(16510, LUT_AMPL_WIDTH - 1),
		5509 => to_unsigned(16513, LUT_AMPL_WIDTH - 1),
		5510 => to_unsigned(16516, LUT_AMPL_WIDTH - 1),
		5511 => to_unsigned(16518, LUT_AMPL_WIDTH - 1),
		5512 => to_unsigned(16521, LUT_AMPL_WIDTH - 1),
		5513 => to_unsigned(16524, LUT_AMPL_WIDTH - 1),
		5514 => to_unsigned(16527, LUT_AMPL_WIDTH - 1),
		5515 => to_unsigned(16529, LUT_AMPL_WIDTH - 1),
		5516 => to_unsigned(16532, LUT_AMPL_WIDTH - 1),
		5517 => to_unsigned(16535, LUT_AMPL_WIDTH - 1),
		5518 => to_unsigned(16537, LUT_AMPL_WIDTH - 1),
		5519 => to_unsigned(16540, LUT_AMPL_WIDTH - 1),
		5520 => to_unsigned(16543, LUT_AMPL_WIDTH - 1),
		5521 => to_unsigned(16546, LUT_AMPL_WIDTH - 1),
		5522 => to_unsigned(16548, LUT_AMPL_WIDTH - 1),
		5523 => to_unsigned(16551, LUT_AMPL_WIDTH - 1),
		5524 => to_unsigned(16554, LUT_AMPL_WIDTH - 1),
		5525 => to_unsigned(16556, LUT_AMPL_WIDTH - 1),
		5526 => to_unsigned(16559, LUT_AMPL_WIDTH - 1),
		5527 => to_unsigned(16562, LUT_AMPL_WIDTH - 1),
		5528 => to_unsigned(16565, LUT_AMPL_WIDTH - 1),
		5529 => to_unsigned(16567, LUT_AMPL_WIDTH - 1),
		5530 => to_unsigned(16570, LUT_AMPL_WIDTH - 1),
		5531 => to_unsigned(16573, LUT_AMPL_WIDTH - 1),
		5532 => to_unsigned(16575, LUT_AMPL_WIDTH - 1),
		5533 => to_unsigned(16578, LUT_AMPL_WIDTH - 1),
		5534 => to_unsigned(16581, LUT_AMPL_WIDTH - 1),
		5535 => to_unsigned(16584, LUT_AMPL_WIDTH - 1),
		5536 => to_unsigned(16586, LUT_AMPL_WIDTH - 1),
		5537 => to_unsigned(16589, LUT_AMPL_WIDTH - 1),
		5538 => to_unsigned(16592, LUT_AMPL_WIDTH - 1),
		5539 => to_unsigned(16594, LUT_AMPL_WIDTH - 1),
		5540 => to_unsigned(16597, LUT_AMPL_WIDTH - 1),
		5541 => to_unsigned(16600, LUT_AMPL_WIDTH - 1),
		5542 => to_unsigned(16602, LUT_AMPL_WIDTH - 1),
		5543 => to_unsigned(16605, LUT_AMPL_WIDTH - 1),
		5544 => to_unsigned(16608, LUT_AMPL_WIDTH - 1),
		5545 => to_unsigned(16611, LUT_AMPL_WIDTH - 1),
		5546 => to_unsigned(16613, LUT_AMPL_WIDTH - 1),
		5547 => to_unsigned(16616, LUT_AMPL_WIDTH - 1),
		5548 => to_unsigned(16619, LUT_AMPL_WIDTH - 1),
		5549 => to_unsigned(16621, LUT_AMPL_WIDTH - 1),
		5550 => to_unsigned(16624, LUT_AMPL_WIDTH - 1),
		5551 => to_unsigned(16627, LUT_AMPL_WIDTH - 1),
		5552 => to_unsigned(16630, LUT_AMPL_WIDTH - 1),
		5553 => to_unsigned(16632, LUT_AMPL_WIDTH - 1),
		5554 => to_unsigned(16635, LUT_AMPL_WIDTH - 1),
		5555 => to_unsigned(16638, LUT_AMPL_WIDTH - 1),
		5556 => to_unsigned(16640, LUT_AMPL_WIDTH - 1),
		5557 => to_unsigned(16643, LUT_AMPL_WIDTH - 1),
		5558 => to_unsigned(16646, LUT_AMPL_WIDTH - 1),
		5559 => to_unsigned(16648, LUT_AMPL_WIDTH - 1),
		5560 => to_unsigned(16651, LUT_AMPL_WIDTH - 1),
		5561 => to_unsigned(16654, LUT_AMPL_WIDTH - 1),
		5562 => to_unsigned(16657, LUT_AMPL_WIDTH - 1),
		5563 => to_unsigned(16659, LUT_AMPL_WIDTH - 1),
		5564 => to_unsigned(16662, LUT_AMPL_WIDTH - 1),
		5565 => to_unsigned(16665, LUT_AMPL_WIDTH - 1),
		5566 => to_unsigned(16667, LUT_AMPL_WIDTH - 1),
		5567 => to_unsigned(16670, LUT_AMPL_WIDTH - 1),
		5568 => to_unsigned(16673, LUT_AMPL_WIDTH - 1),
		5569 => to_unsigned(16676, LUT_AMPL_WIDTH - 1),
		5570 => to_unsigned(16678, LUT_AMPL_WIDTH - 1),
		5571 => to_unsigned(16681, LUT_AMPL_WIDTH - 1),
		5572 => to_unsigned(16684, LUT_AMPL_WIDTH - 1),
		5573 => to_unsigned(16686, LUT_AMPL_WIDTH - 1),
		5574 => to_unsigned(16689, LUT_AMPL_WIDTH - 1),
		5575 => to_unsigned(16692, LUT_AMPL_WIDTH - 1),
		5576 => to_unsigned(16694, LUT_AMPL_WIDTH - 1),
		5577 => to_unsigned(16697, LUT_AMPL_WIDTH - 1),
		5578 => to_unsigned(16700, LUT_AMPL_WIDTH - 1),
		5579 => to_unsigned(16703, LUT_AMPL_WIDTH - 1),
		5580 => to_unsigned(16705, LUT_AMPL_WIDTH - 1),
		5581 => to_unsigned(16708, LUT_AMPL_WIDTH - 1),
		5582 => to_unsigned(16711, LUT_AMPL_WIDTH - 1),
		5583 => to_unsigned(16713, LUT_AMPL_WIDTH - 1),
		5584 => to_unsigned(16716, LUT_AMPL_WIDTH - 1),
		5585 => to_unsigned(16719, LUT_AMPL_WIDTH - 1),
		5586 => to_unsigned(16721, LUT_AMPL_WIDTH - 1),
		5587 => to_unsigned(16724, LUT_AMPL_WIDTH - 1),
		5588 => to_unsigned(16727, LUT_AMPL_WIDTH - 1),
		5589 => to_unsigned(16730, LUT_AMPL_WIDTH - 1),
		5590 => to_unsigned(16732, LUT_AMPL_WIDTH - 1),
		5591 => to_unsigned(16735, LUT_AMPL_WIDTH - 1),
		5592 => to_unsigned(16738, LUT_AMPL_WIDTH - 1),
		5593 => to_unsigned(16740, LUT_AMPL_WIDTH - 1),
		5594 => to_unsigned(16743, LUT_AMPL_WIDTH - 1),
		5595 => to_unsigned(16746, LUT_AMPL_WIDTH - 1),
		5596 => to_unsigned(16749, LUT_AMPL_WIDTH - 1),
		5597 => to_unsigned(16751, LUT_AMPL_WIDTH - 1),
		5598 => to_unsigned(16754, LUT_AMPL_WIDTH - 1),
		5599 => to_unsigned(16757, LUT_AMPL_WIDTH - 1),
		5600 => to_unsigned(16759, LUT_AMPL_WIDTH - 1),
		5601 => to_unsigned(16762, LUT_AMPL_WIDTH - 1),
		5602 => to_unsigned(16765, LUT_AMPL_WIDTH - 1),
		5603 => to_unsigned(16767, LUT_AMPL_WIDTH - 1),
		5604 => to_unsigned(16770, LUT_AMPL_WIDTH - 1),
		5605 => to_unsigned(16773, LUT_AMPL_WIDTH - 1),
		5606 => to_unsigned(16775, LUT_AMPL_WIDTH - 1),
		5607 => to_unsigned(16778, LUT_AMPL_WIDTH - 1),
		5608 => to_unsigned(16781, LUT_AMPL_WIDTH - 1),
		5609 => to_unsigned(16784, LUT_AMPL_WIDTH - 1),
		5610 => to_unsigned(16786, LUT_AMPL_WIDTH - 1),
		5611 => to_unsigned(16789, LUT_AMPL_WIDTH - 1),
		5612 => to_unsigned(16792, LUT_AMPL_WIDTH - 1),
		5613 => to_unsigned(16794, LUT_AMPL_WIDTH - 1),
		5614 => to_unsigned(16797, LUT_AMPL_WIDTH - 1),
		5615 => to_unsigned(16800, LUT_AMPL_WIDTH - 1),
		5616 => to_unsigned(16802, LUT_AMPL_WIDTH - 1),
		5617 => to_unsigned(16805, LUT_AMPL_WIDTH - 1),
		5618 => to_unsigned(16808, LUT_AMPL_WIDTH - 1),
		5619 => to_unsigned(16811, LUT_AMPL_WIDTH - 1),
		5620 => to_unsigned(16813, LUT_AMPL_WIDTH - 1),
		5621 => to_unsigned(16816, LUT_AMPL_WIDTH - 1),
		5622 => to_unsigned(16819, LUT_AMPL_WIDTH - 1),
		5623 => to_unsigned(16821, LUT_AMPL_WIDTH - 1),
		5624 => to_unsigned(16824, LUT_AMPL_WIDTH - 1),
		5625 => to_unsigned(16827, LUT_AMPL_WIDTH - 1),
		5626 => to_unsigned(16829, LUT_AMPL_WIDTH - 1),
		5627 => to_unsigned(16832, LUT_AMPL_WIDTH - 1),
		5628 => to_unsigned(16835, LUT_AMPL_WIDTH - 1),
		5629 => to_unsigned(16838, LUT_AMPL_WIDTH - 1),
		5630 => to_unsigned(16840, LUT_AMPL_WIDTH - 1),
		5631 => to_unsigned(16843, LUT_AMPL_WIDTH - 1),
		5632 => to_unsigned(16846, LUT_AMPL_WIDTH - 1),
		5633 => to_unsigned(16848, LUT_AMPL_WIDTH - 1),
		5634 => to_unsigned(16851, LUT_AMPL_WIDTH - 1),
		5635 => to_unsigned(16854, LUT_AMPL_WIDTH - 1),
		5636 => to_unsigned(16856, LUT_AMPL_WIDTH - 1),
		5637 => to_unsigned(16859, LUT_AMPL_WIDTH - 1),
		5638 => to_unsigned(16862, LUT_AMPL_WIDTH - 1),
		5639 => to_unsigned(16864, LUT_AMPL_WIDTH - 1),
		5640 => to_unsigned(16867, LUT_AMPL_WIDTH - 1),
		5641 => to_unsigned(16870, LUT_AMPL_WIDTH - 1),
		5642 => to_unsigned(16873, LUT_AMPL_WIDTH - 1),
		5643 => to_unsigned(16875, LUT_AMPL_WIDTH - 1),
		5644 => to_unsigned(16878, LUT_AMPL_WIDTH - 1),
		5645 => to_unsigned(16881, LUT_AMPL_WIDTH - 1),
		5646 => to_unsigned(16883, LUT_AMPL_WIDTH - 1),
		5647 => to_unsigned(16886, LUT_AMPL_WIDTH - 1),
		5648 => to_unsigned(16889, LUT_AMPL_WIDTH - 1),
		5649 => to_unsigned(16891, LUT_AMPL_WIDTH - 1),
		5650 => to_unsigned(16894, LUT_AMPL_WIDTH - 1),
		5651 => to_unsigned(16897, LUT_AMPL_WIDTH - 1),
		5652 => to_unsigned(16899, LUT_AMPL_WIDTH - 1),
		5653 => to_unsigned(16902, LUT_AMPL_WIDTH - 1),
		5654 => to_unsigned(16905, LUT_AMPL_WIDTH - 1),
		5655 => to_unsigned(16908, LUT_AMPL_WIDTH - 1),
		5656 => to_unsigned(16910, LUT_AMPL_WIDTH - 1),
		5657 => to_unsigned(16913, LUT_AMPL_WIDTH - 1),
		5658 => to_unsigned(16916, LUT_AMPL_WIDTH - 1),
		5659 => to_unsigned(16918, LUT_AMPL_WIDTH - 1),
		5660 => to_unsigned(16921, LUT_AMPL_WIDTH - 1),
		5661 => to_unsigned(16924, LUT_AMPL_WIDTH - 1),
		5662 => to_unsigned(16926, LUT_AMPL_WIDTH - 1),
		5663 => to_unsigned(16929, LUT_AMPL_WIDTH - 1),
		5664 => to_unsigned(16932, LUT_AMPL_WIDTH - 1),
		5665 => to_unsigned(16934, LUT_AMPL_WIDTH - 1),
		5666 => to_unsigned(16937, LUT_AMPL_WIDTH - 1),
		5667 => to_unsigned(16940, LUT_AMPL_WIDTH - 1),
		5668 => to_unsigned(16943, LUT_AMPL_WIDTH - 1),
		5669 => to_unsigned(16945, LUT_AMPL_WIDTH - 1),
		5670 => to_unsigned(16948, LUT_AMPL_WIDTH - 1),
		5671 => to_unsigned(16951, LUT_AMPL_WIDTH - 1),
		5672 => to_unsigned(16953, LUT_AMPL_WIDTH - 1),
		5673 => to_unsigned(16956, LUT_AMPL_WIDTH - 1),
		5674 => to_unsigned(16959, LUT_AMPL_WIDTH - 1),
		5675 => to_unsigned(16961, LUT_AMPL_WIDTH - 1),
		5676 => to_unsigned(16964, LUT_AMPL_WIDTH - 1),
		5677 => to_unsigned(16967, LUT_AMPL_WIDTH - 1),
		5678 => to_unsigned(16969, LUT_AMPL_WIDTH - 1),
		5679 => to_unsigned(16972, LUT_AMPL_WIDTH - 1),
		5680 => to_unsigned(16975, LUT_AMPL_WIDTH - 1),
		5681 => to_unsigned(16977, LUT_AMPL_WIDTH - 1),
		5682 => to_unsigned(16980, LUT_AMPL_WIDTH - 1),
		5683 => to_unsigned(16983, LUT_AMPL_WIDTH - 1),
		5684 => to_unsigned(16986, LUT_AMPL_WIDTH - 1),
		5685 => to_unsigned(16988, LUT_AMPL_WIDTH - 1),
		5686 => to_unsigned(16991, LUT_AMPL_WIDTH - 1),
		5687 => to_unsigned(16994, LUT_AMPL_WIDTH - 1),
		5688 => to_unsigned(16996, LUT_AMPL_WIDTH - 1),
		5689 => to_unsigned(16999, LUT_AMPL_WIDTH - 1),
		5690 => to_unsigned(17002, LUT_AMPL_WIDTH - 1),
		5691 => to_unsigned(17004, LUT_AMPL_WIDTH - 1),
		5692 => to_unsigned(17007, LUT_AMPL_WIDTH - 1),
		5693 => to_unsigned(17010, LUT_AMPL_WIDTH - 1),
		5694 => to_unsigned(17012, LUT_AMPL_WIDTH - 1),
		5695 => to_unsigned(17015, LUT_AMPL_WIDTH - 1),
		5696 => to_unsigned(17018, LUT_AMPL_WIDTH - 1),
		5697 => to_unsigned(17020, LUT_AMPL_WIDTH - 1),
		5698 => to_unsigned(17023, LUT_AMPL_WIDTH - 1),
		5699 => to_unsigned(17026, LUT_AMPL_WIDTH - 1),
		5700 => to_unsigned(17028, LUT_AMPL_WIDTH - 1),
		5701 => to_unsigned(17031, LUT_AMPL_WIDTH - 1),
		5702 => to_unsigned(17034, LUT_AMPL_WIDTH - 1),
		5703 => to_unsigned(17037, LUT_AMPL_WIDTH - 1),
		5704 => to_unsigned(17039, LUT_AMPL_WIDTH - 1),
		5705 => to_unsigned(17042, LUT_AMPL_WIDTH - 1),
		5706 => to_unsigned(17045, LUT_AMPL_WIDTH - 1),
		5707 => to_unsigned(17047, LUT_AMPL_WIDTH - 1),
		5708 => to_unsigned(17050, LUT_AMPL_WIDTH - 1),
		5709 => to_unsigned(17053, LUT_AMPL_WIDTH - 1),
		5710 => to_unsigned(17055, LUT_AMPL_WIDTH - 1),
		5711 => to_unsigned(17058, LUT_AMPL_WIDTH - 1),
		5712 => to_unsigned(17061, LUT_AMPL_WIDTH - 1),
		5713 => to_unsigned(17063, LUT_AMPL_WIDTH - 1),
		5714 => to_unsigned(17066, LUT_AMPL_WIDTH - 1),
		5715 => to_unsigned(17069, LUT_AMPL_WIDTH - 1),
		5716 => to_unsigned(17071, LUT_AMPL_WIDTH - 1),
		5717 => to_unsigned(17074, LUT_AMPL_WIDTH - 1),
		5718 => to_unsigned(17077, LUT_AMPL_WIDTH - 1),
		5719 => to_unsigned(17079, LUT_AMPL_WIDTH - 1),
		5720 => to_unsigned(17082, LUT_AMPL_WIDTH - 1),
		5721 => to_unsigned(17085, LUT_AMPL_WIDTH - 1),
		5722 => to_unsigned(17087, LUT_AMPL_WIDTH - 1),
		5723 => to_unsigned(17090, LUT_AMPL_WIDTH - 1),
		5724 => to_unsigned(17093, LUT_AMPL_WIDTH - 1),
		5725 => to_unsigned(17096, LUT_AMPL_WIDTH - 1),
		5726 => to_unsigned(17098, LUT_AMPL_WIDTH - 1),
		5727 => to_unsigned(17101, LUT_AMPL_WIDTH - 1),
		5728 => to_unsigned(17104, LUT_AMPL_WIDTH - 1),
		5729 => to_unsigned(17106, LUT_AMPL_WIDTH - 1),
		5730 => to_unsigned(17109, LUT_AMPL_WIDTH - 1),
		5731 => to_unsigned(17112, LUT_AMPL_WIDTH - 1),
		5732 => to_unsigned(17114, LUT_AMPL_WIDTH - 1),
		5733 => to_unsigned(17117, LUT_AMPL_WIDTH - 1),
		5734 => to_unsigned(17120, LUT_AMPL_WIDTH - 1),
		5735 => to_unsigned(17122, LUT_AMPL_WIDTH - 1),
		5736 => to_unsigned(17125, LUT_AMPL_WIDTH - 1),
		5737 => to_unsigned(17128, LUT_AMPL_WIDTH - 1),
		5738 => to_unsigned(17130, LUT_AMPL_WIDTH - 1),
		5739 => to_unsigned(17133, LUT_AMPL_WIDTH - 1),
		5740 => to_unsigned(17136, LUT_AMPL_WIDTH - 1),
		5741 => to_unsigned(17138, LUT_AMPL_WIDTH - 1),
		5742 => to_unsigned(17141, LUT_AMPL_WIDTH - 1),
		5743 => to_unsigned(17144, LUT_AMPL_WIDTH - 1),
		5744 => to_unsigned(17146, LUT_AMPL_WIDTH - 1),
		5745 => to_unsigned(17149, LUT_AMPL_WIDTH - 1),
		5746 => to_unsigned(17152, LUT_AMPL_WIDTH - 1),
		5747 => to_unsigned(17154, LUT_AMPL_WIDTH - 1),
		5748 => to_unsigned(17157, LUT_AMPL_WIDTH - 1),
		5749 => to_unsigned(17160, LUT_AMPL_WIDTH - 1),
		5750 => to_unsigned(17162, LUT_AMPL_WIDTH - 1),
		5751 => to_unsigned(17165, LUT_AMPL_WIDTH - 1),
		5752 => to_unsigned(17168, LUT_AMPL_WIDTH - 1),
		5753 => to_unsigned(17171, LUT_AMPL_WIDTH - 1),
		5754 => to_unsigned(17173, LUT_AMPL_WIDTH - 1),
		5755 => to_unsigned(17176, LUT_AMPL_WIDTH - 1),
		5756 => to_unsigned(17179, LUT_AMPL_WIDTH - 1),
		5757 => to_unsigned(17181, LUT_AMPL_WIDTH - 1),
		5758 => to_unsigned(17184, LUT_AMPL_WIDTH - 1),
		5759 => to_unsigned(17187, LUT_AMPL_WIDTH - 1),
		5760 => to_unsigned(17189, LUT_AMPL_WIDTH - 1),
		5761 => to_unsigned(17192, LUT_AMPL_WIDTH - 1),
		5762 => to_unsigned(17195, LUT_AMPL_WIDTH - 1),
		5763 => to_unsigned(17197, LUT_AMPL_WIDTH - 1),
		5764 => to_unsigned(17200, LUT_AMPL_WIDTH - 1),
		5765 => to_unsigned(17203, LUT_AMPL_WIDTH - 1),
		5766 => to_unsigned(17205, LUT_AMPL_WIDTH - 1),
		5767 => to_unsigned(17208, LUT_AMPL_WIDTH - 1),
		5768 => to_unsigned(17211, LUT_AMPL_WIDTH - 1),
		5769 => to_unsigned(17213, LUT_AMPL_WIDTH - 1),
		5770 => to_unsigned(17216, LUT_AMPL_WIDTH - 1),
		5771 => to_unsigned(17219, LUT_AMPL_WIDTH - 1),
		5772 => to_unsigned(17221, LUT_AMPL_WIDTH - 1),
		5773 => to_unsigned(17224, LUT_AMPL_WIDTH - 1),
		5774 => to_unsigned(17227, LUT_AMPL_WIDTH - 1),
		5775 => to_unsigned(17229, LUT_AMPL_WIDTH - 1),
		5776 => to_unsigned(17232, LUT_AMPL_WIDTH - 1),
		5777 => to_unsigned(17235, LUT_AMPL_WIDTH - 1),
		5778 => to_unsigned(17237, LUT_AMPL_WIDTH - 1),
		5779 => to_unsigned(17240, LUT_AMPL_WIDTH - 1),
		5780 => to_unsigned(17243, LUT_AMPL_WIDTH - 1),
		5781 => to_unsigned(17245, LUT_AMPL_WIDTH - 1),
		5782 => to_unsigned(17248, LUT_AMPL_WIDTH - 1),
		5783 => to_unsigned(17251, LUT_AMPL_WIDTH - 1),
		5784 => to_unsigned(17253, LUT_AMPL_WIDTH - 1),
		5785 => to_unsigned(17256, LUT_AMPL_WIDTH - 1),
		5786 => to_unsigned(17259, LUT_AMPL_WIDTH - 1),
		5787 => to_unsigned(17261, LUT_AMPL_WIDTH - 1),
		5788 => to_unsigned(17264, LUT_AMPL_WIDTH - 1),
		5789 => to_unsigned(17267, LUT_AMPL_WIDTH - 1),
		5790 => to_unsigned(17269, LUT_AMPL_WIDTH - 1),
		5791 => to_unsigned(17272, LUT_AMPL_WIDTH - 1),
		5792 => to_unsigned(17275, LUT_AMPL_WIDTH - 1),
		5793 => to_unsigned(17277, LUT_AMPL_WIDTH - 1),
		5794 => to_unsigned(17280, LUT_AMPL_WIDTH - 1),
		5795 => to_unsigned(17283, LUT_AMPL_WIDTH - 1),
		5796 => to_unsigned(17285, LUT_AMPL_WIDTH - 1),
		5797 => to_unsigned(17288, LUT_AMPL_WIDTH - 1),
		5798 => to_unsigned(17291, LUT_AMPL_WIDTH - 1),
		5799 => to_unsigned(17293, LUT_AMPL_WIDTH - 1),
		5800 => to_unsigned(17296, LUT_AMPL_WIDTH - 1),
		5801 => to_unsigned(17299, LUT_AMPL_WIDTH - 1),
		5802 => to_unsigned(17301, LUT_AMPL_WIDTH - 1),
		5803 => to_unsigned(17304, LUT_AMPL_WIDTH - 1),
		5804 => to_unsigned(17307, LUT_AMPL_WIDTH - 1),
		5805 => to_unsigned(17309, LUT_AMPL_WIDTH - 1),
		5806 => to_unsigned(17312, LUT_AMPL_WIDTH - 1),
		5807 => to_unsigned(17315, LUT_AMPL_WIDTH - 1),
		5808 => to_unsigned(17317, LUT_AMPL_WIDTH - 1),
		5809 => to_unsigned(17320, LUT_AMPL_WIDTH - 1),
		5810 => to_unsigned(17323, LUT_AMPL_WIDTH - 1),
		5811 => to_unsigned(17325, LUT_AMPL_WIDTH - 1),
		5812 => to_unsigned(17328, LUT_AMPL_WIDTH - 1),
		5813 => to_unsigned(17331, LUT_AMPL_WIDTH - 1),
		5814 => to_unsigned(17333, LUT_AMPL_WIDTH - 1),
		5815 => to_unsigned(17336, LUT_AMPL_WIDTH - 1),
		5816 => to_unsigned(17339, LUT_AMPL_WIDTH - 1),
		5817 => to_unsigned(17341, LUT_AMPL_WIDTH - 1),
		5818 => to_unsigned(17344, LUT_AMPL_WIDTH - 1),
		5819 => to_unsigned(17347, LUT_AMPL_WIDTH - 1),
		5820 => to_unsigned(17349, LUT_AMPL_WIDTH - 1),
		5821 => to_unsigned(17352, LUT_AMPL_WIDTH - 1),
		5822 => to_unsigned(17355, LUT_AMPL_WIDTH - 1),
		5823 => to_unsigned(17357, LUT_AMPL_WIDTH - 1),
		5824 => to_unsigned(17360, LUT_AMPL_WIDTH - 1),
		5825 => to_unsigned(17363, LUT_AMPL_WIDTH - 1),
		5826 => to_unsigned(17365, LUT_AMPL_WIDTH - 1),
		5827 => to_unsigned(17368, LUT_AMPL_WIDTH - 1),
		5828 => to_unsigned(17371, LUT_AMPL_WIDTH - 1),
		5829 => to_unsigned(17373, LUT_AMPL_WIDTH - 1),
		5830 => to_unsigned(17376, LUT_AMPL_WIDTH - 1),
		5831 => to_unsigned(17379, LUT_AMPL_WIDTH - 1),
		5832 => to_unsigned(17381, LUT_AMPL_WIDTH - 1),
		5833 => to_unsigned(17384, LUT_AMPL_WIDTH - 1),
		5834 => to_unsigned(17387, LUT_AMPL_WIDTH - 1),
		5835 => to_unsigned(17389, LUT_AMPL_WIDTH - 1),
		5836 => to_unsigned(17392, LUT_AMPL_WIDTH - 1),
		5837 => to_unsigned(17395, LUT_AMPL_WIDTH - 1),
		5838 => to_unsigned(17397, LUT_AMPL_WIDTH - 1),
		5839 => to_unsigned(17400, LUT_AMPL_WIDTH - 1),
		5840 => to_unsigned(17403, LUT_AMPL_WIDTH - 1),
		5841 => to_unsigned(17405, LUT_AMPL_WIDTH - 1),
		5842 => to_unsigned(17408, LUT_AMPL_WIDTH - 1),
		5843 => to_unsigned(17411, LUT_AMPL_WIDTH - 1),
		5844 => to_unsigned(17413, LUT_AMPL_WIDTH - 1),
		5845 => to_unsigned(17416, LUT_AMPL_WIDTH - 1),
		5846 => to_unsigned(17419, LUT_AMPL_WIDTH - 1),
		5847 => to_unsigned(17421, LUT_AMPL_WIDTH - 1),
		5848 => to_unsigned(17424, LUT_AMPL_WIDTH - 1),
		5849 => to_unsigned(17427, LUT_AMPL_WIDTH - 1),
		5850 => to_unsigned(17429, LUT_AMPL_WIDTH - 1),
		5851 => to_unsigned(17432, LUT_AMPL_WIDTH - 1),
		5852 => to_unsigned(17435, LUT_AMPL_WIDTH - 1),
		5853 => to_unsigned(17437, LUT_AMPL_WIDTH - 1),
		5854 => to_unsigned(17440, LUT_AMPL_WIDTH - 1),
		5855 => to_unsigned(17443, LUT_AMPL_WIDTH - 1),
		5856 => to_unsigned(17445, LUT_AMPL_WIDTH - 1),
		5857 => to_unsigned(17448, LUT_AMPL_WIDTH - 1),
		5858 => to_unsigned(17451, LUT_AMPL_WIDTH - 1),
		5859 => to_unsigned(17453, LUT_AMPL_WIDTH - 1),
		5860 => to_unsigned(17456, LUT_AMPL_WIDTH - 1),
		5861 => to_unsigned(17459, LUT_AMPL_WIDTH - 1),
		5862 => to_unsigned(17461, LUT_AMPL_WIDTH - 1),
		5863 => to_unsigned(17464, LUT_AMPL_WIDTH - 1),
		5864 => to_unsigned(17467, LUT_AMPL_WIDTH - 1),
		5865 => to_unsigned(17469, LUT_AMPL_WIDTH - 1),
		5866 => to_unsigned(17472, LUT_AMPL_WIDTH - 1),
		5867 => to_unsigned(17474, LUT_AMPL_WIDTH - 1),
		5868 => to_unsigned(17477, LUT_AMPL_WIDTH - 1),
		5869 => to_unsigned(17480, LUT_AMPL_WIDTH - 1),
		5870 => to_unsigned(17482, LUT_AMPL_WIDTH - 1),
		5871 => to_unsigned(17485, LUT_AMPL_WIDTH - 1),
		5872 => to_unsigned(17488, LUT_AMPL_WIDTH - 1),
		5873 => to_unsigned(17490, LUT_AMPL_WIDTH - 1),
		5874 => to_unsigned(17493, LUT_AMPL_WIDTH - 1),
		5875 => to_unsigned(17496, LUT_AMPL_WIDTH - 1),
		5876 => to_unsigned(17498, LUT_AMPL_WIDTH - 1),
		5877 => to_unsigned(17501, LUT_AMPL_WIDTH - 1),
		5878 => to_unsigned(17504, LUT_AMPL_WIDTH - 1),
		5879 => to_unsigned(17506, LUT_AMPL_WIDTH - 1),
		5880 => to_unsigned(17509, LUT_AMPL_WIDTH - 1),
		5881 => to_unsigned(17512, LUT_AMPL_WIDTH - 1),
		5882 => to_unsigned(17514, LUT_AMPL_WIDTH - 1),
		5883 => to_unsigned(17517, LUT_AMPL_WIDTH - 1),
		5884 => to_unsigned(17520, LUT_AMPL_WIDTH - 1),
		5885 => to_unsigned(17522, LUT_AMPL_WIDTH - 1),
		5886 => to_unsigned(17525, LUT_AMPL_WIDTH - 1),
		5887 => to_unsigned(17528, LUT_AMPL_WIDTH - 1),
		5888 => to_unsigned(17530, LUT_AMPL_WIDTH - 1),
		5889 => to_unsigned(17533, LUT_AMPL_WIDTH - 1),
		5890 => to_unsigned(17536, LUT_AMPL_WIDTH - 1),
		5891 => to_unsigned(17538, LUT_AMPL_WIDTH - 1),
		5892 => to_unsigned(17541, LUT_AMPL_WIDTH - 1),
		5893 => to_unsigned(17544, LUT_AMPL_WIDTH - 1),
		5894 => to_unsigned(17546, LUT_AMPL_WIDTH - 1),
		5895 => to_unsigned(17549, LUT_AMPL_WIDTH - 1),
		5896 => to_unsigned(17551, LUT_AMPL_WIDTH - 1),
		5897 => to_unsigned(17554, LUT_AMPL_WIDTH - 1),
		5898 => to_unsigned(17557, LUT_AMPL_WIDTH - 1),
		5899 => to_unsigned(17559, LUT_AMPL_WIDTH - 1),
		5900 => to_unsigned(17562, LUT_AMPL_WIDTH - 1),
		5901 => to_unsigned(17565, LUT_AMPL_WIDTH - 1),
		5902 => to_unsigned(17567, LUT_AMPL_WIDTH - 1),
		5903 => to_unsigned(17570, LUT_AMPL_WIDTH - 1),
		5904 => to_unsigned(17573, LUT_AMPL_WIDTH - 1),
		5905 => to_unsigned(17575, LUT_AMPL_WIDTH - 1),
		5906 => to_unsigned(17578, LUT_AMPL_WIDTH - 1),
		5907 => to_unsigned(17581, LUT_AMPL_WIDTH - 1),
		5908 => to_unsigned(17583, LUT_AMPL_WIDTH - 1),
		5909 => to_unsigned(17586, LUT_AMPL_WIDTH - 1),
		5910 => to_unsigned(17589, LUT_AMPL_WIDTH - 1),
		5911 => to_unsigned(17591, LUT_AMPL_WIDTH - 1),
		5912 => to_unsigned(17594, LUT_AMPL_WIDTH - 1),
		5913 => to_unsigned(17597, LUT_AMPL_WIDTH - 1),
		5914 => to_unsigned(17599, LUT_AMPL_WIDTH - 1),
		5915 => to_unsigned(17602, LUT_AMPL_WIDTH - 1),
		5916 => to_unsigned(17605, LUT_AMPL_WIDTH - 1),
		5917 => to_unsigned(17607, LUT_AMPL_WIDTH - 1),
		5918 => to_unsigned(17610, LUT_AMPL_WIDTH - 1),
		5919 => to_unsigned(17612, LUT_AMPL_WIDTH - 1),
		5920 => to_unsigned(17615, LUT_AMPL_WIDTH - 1),
		5921 => to_unsigned(17618, LUT_AMPL_WIDTH - 1),
		5922 => to_unsigned(17620, LUT_AMPL_WIDTH - 1),
		5923 => to_unsigned(17623, LUT_AMPL_WIDTH - 1),
		5924 => to_unsigned(17626, LUT_AMPL_WIDTH - 1),
		5925 => to_unsigned(17628, LUT_AMPL_WIDTH - 1),
		5926 => to_unsigned(17631, LUT_AMPL_WIDTH - 1),
		5927 => to_unsigned(17634, LUT_AMPL_WIDTH - 1),
		5928 => to_unsigned(17636, LUT_AMPL_WIDTH - 1),
		5929 => to_unsigned(17639, LUT_AMPL_WIDTH - 1),
		5930 => to_unsigned(17642, LUT_AMPL_WIDTH - 1),
		5931 => to_unsigned(17644, LUT_AMPL_WIDTH - 1),
		5932 => to_unsigned(17647, LUT_AMPL_WIDTH - 1),
		5933 => to_unsigned(17650, LUT_AMPL_WIDTH - 1),
		5934 => to_unsigned(17652, LUT_AMPL_WIDTH - 1),
		5935 => to_unsigned(17655, LUT_AMPL_WIDTH - 1),
		5936 => to_unsigned(17657, LUT_AMPL_WIDTH - 1),
		5937 => to_unsigned(17660, LUT_AMPL_WIDTH - 1),
		5938 => to_unsigned(17663, LUT_AMPL_WIDTH - 1),
		5939 => to_unsigned(17665, LUT_AMPL_WIDTH - 1),
		5940 => to_unsigned(17668, LUT_AMPL_WIDTH - 1),
		5941 => to_unsigned(17671, LUT_AMPL_WIDTH - 1),
		5942 => to_unsigned(17673, LUT_AMPL_WIDTH - 1),
		5943 => to_unsigned(17676, LUT_AMPL_WIDTH - 1),
		5944 => to_unsigned(17679, LUT_AMPL_WIDTH - 1),
		5945 => to_unsigned(17681, LUT_AMPL_WIDTH - 1),
		5946 => to_unsigned(17684, LUT_AMPL_WIDTH - 1),
		5947 => to_unsigned(17687, LUT_AMPL_WIDTH - 1),
		5948 => to_unsigned(17689, LUT_AMPL_WIDTH - 1),
		5949 => to_unsigned(17692, LUT_AMPL_WIDTH - 1),
		5950 => to_unsigned(17695, LUT_AMPL_WIDTH - 1),
		5951 => to_unsigned(17697, LUT_AMPL_WIDTH - 1),
		5952 => to_unsigned(17700, LUT_AMPL_WIDTH - 1),
		5953 => to_unsigned(17702, LUT_AMPL_WIDTH - 1),
		5954 => to_unsigned(17705, LUT_AMPL_WIDTH - 1),
		5955 => to_unsigned(17708, LUT_AMPL_WIDTH - 1),
		5956 => to_unsigned(17710, LUT_AMPL_WIDTH - 1),
		5957 => to_unsigned(17713, LUT_AMPL_WIDTH - 1),
		5958 => to_unsigned(17716, LUT_AMPL_WIDTH - 1),
		5959 => to_unsigned(17718, LUT_AMPL_WIDTH - 1),
		5960 => to_unsigned(17721, LUT_AMPL_WIDTH - 1),
		5961 => to_unsigned(17724, LUT_AMPL_WIDTH - 1),
		5962 => to_unsigned(17726, LUT_AMPL_WIDTH - 1),
		5963 => to_unsigned(17729, LUT_AMPL_WIDTH - 1),
		5964 => to_unsigned(17732, LUT_AMPL_WIDTH - 1),
		5965 => to_unsigned(17734, LUT_AMPL_WIDTH - 1),
		5966 => to_unsigned(17737, LUT_AMPL_WIDTH - 1),
		5967 => to_unsigned(17739, LUT_AMPL_WIDTH - 1),
		5968 => to_unsigned(17742, LUT_AMPL_WIDTH - 1),
		5969 => to_unsigned(17745, LUT_AMPL_WIDTH - 1),
		5970 => to_unsigned(17747, LUT_AMPL_WIDTH - 1),
		5971 => to_unsigned(17750, LUT_AMPL_WIDTH - 1),
		5972 => to_unsigned(17753, LUT_AMPL_WIDTH - 1),
		5973 => to_unsigned(17755, LUT_AMPL_WIDTH - 1),
		5974 => to_unsigned(17758, LUT_AMPL_WIDTH - 1),
		5975 => to_unsigned(17761, LUT_AMPL_WIDTH - 1),
		5976 => to_unsigned(17763, LUT_AMPL_WIDTH - 1),
		5977 => to_unsigned(17766, LUT_AMPL_WIDTH - 1),
		5978 => to_unsigned(17768, LUT_AMPL_WIDTH - 1),
		5979 => to_unsigned(17771, LUT_AMPL_WIDTH - 1),
		5980 => to_unsigned(17774, LUT_AMPL_WIDTH - 1),
		5981 => to_unsigned(17776, LUT_AMPL_WIDTH - 1),
		5982 => to_unsigned(17779, LUT_AMPL_WIDTH - 1),
		5983 => to_unsigned(17782, LUT_AMPL_WIDTH - 1),
		5984 => to_unsigned(17784, LUT_AMPL_WIDTH - 1),
		5985 => to_unsigned(17787, LUT_AMPL_WIDTH - 1),
		5986 => to_unsigned(17790, LUT_AMPL_WIDTH - 1),
		5987 => to_unsigned(17792, LUT_AMPL_WIDTH - 1),
		5988 => to_unsigned(17795, LUT_AMPL_WIDTH - 1),
		5989 => to_unsigned(17798, LUT_AMPL_WIDTH - 1),
		5990 => to_unsigned(17800, LUT_AMPL_WIDTH - 1),
		5991 => to_unsigned(17803, LUT_AMPL_WIDTH - 1),
		5992 => to_unsigned(17805, LUT_AMPL_WIDTH - 1),
		5993 => to_unsigned(17808, LUT_AMPL_WIDTH - 1),
		5994 => to_unsigned(17811, LUT_AMPL_WIDTH - 1),
		5995 => to_unsigned(17813, LUT_AMPL_WIDTH - 1),
		5996 => to_unsigned(17816, LUT_AMPL_WIDTH - 1),
		5997 => to_unsigned(17819, LUT_AMPL_WIDTH - 1),
		5998 => to_unsigned(17821, LUT_AMPL_WIDTH - 1),
		5999 => to_unsigned(17824, LUT_AMPL_WIDTH - 1),
		6000 => to_unsigned(17827, LUT_AMPL_WIDTH - 1),
		6001 => to_unsigned(17829, LUT_AMPL_WIDTH - 1),
		6002 => to_unsigned(17832, LUT_AMPL_WIDTH - 1),
		6003 => to_unsigned(17834, LUT_AMPL_WIDTH - 1),
		6004 => to_unsigned(17837, LUT_AMPL_WIDTH - 1),
		6005 => to_unsigned(17840, LUT_AMPL_WIDTH - 1),
		6006 => to_unsigned(17842, LUT_AMPL_WIDTH - 1),
		6007 => to_unsigned(17845, LUT_AMPL_WIDTH - 1),
		6008 => to_unsigned(17848, LUT_AMPL_WIDTH - 1),
		6009 => to_unsigned(17850, LUT_AMPL_WIDTH - 1),
		6010 => to_unsigned(17853, LUT_AMPL_WIDTH - 1),
		6011 => to_unsigned(17855, LUT_AMPL_WIDTH - 1),
		6012 => to_unsigned(17858, LUT_AMPL_WIDTH - 1),
		6013 => to_unsigned(17861, LUT_AMPL_WIDTH - 1),
		6014 => to_unsigned(17863, LUT_AMPL_WIDTH - 1),
		6015 => to_unsigned(17866, LUT_AMPL_WIDTH - 1),
		6016 => to_unsigned(17869, LUT_AMPL_WIDTH - 1),
		6017 => to_unsigned(17871, LUT_AMPL_WIDTH - 1),
		6018 => to_unsigned(17874, LUT_AMPL_WIDTH - 1),
		6019 => to_unsigned(17877, LUT_AMPL_WIDTH - 1),
		6020 => to_unsigned(17879, LUT_AMPL_WIDTH - 1),
		6021 => to_unsigned(17882, LUT_AMPL_WIDTH - 1),
		6022 => to_unsigned(17884, LUT_AMPL_WIDTH - 1),
		6023 => to_unsigned(17887, LUT_AMPL_WIDTH - 1),
		6024 => to_unsigned(17890, LUT_AMPL_WIDTH - 1),
		6025 => to_unsigned(17892, LUT_AMPL_WIDTH - 1),
		6026 => to_unsigned(17895, LUT_AMPL_WIDTH - 1),
		6027 => to_unsigned(17898, LUT_AMPL_WIDTH - 1),
		6028 => to_unsigned(17900, LUT_AMPL_WIDTH - 1),
		6029 => to_unsigned(17903, LUT_AMPL_WIDTH - 1),
		6030 => to_unsigned(17906, LUT_AMPL_WIDTH - 1),
		6031 => to_unsigned(17908, LUT_AMPL_WIDTH - 1),
		6032 => to_unsigned(17911, LUT_AMPL_WIDTH - 1),
		6033 => to_unsigned(17913, LUT_AMPL_WIDTH - 1),
		6034 => to_unsigned(17916, LUT_AMPL_WIDTH - 1),
		6035 => to_unsigned(17919, LUT_AMPL_WIDTH - 1),
		6036 => to_unsigned(17921, LUT_AMPL_WIDTH - 1),
		6037 => to_unsigned(17924, LUT_AMPL_WIDTH - 1),
		6038 => to_unsigned(17927, LUT_AMPL_WIDTH - 1),
		6039 => to_unsigned(17929, LUT_AMPL_WIDTH - 1),
		6040 => to_unsigned(17932, LUT_AMPL_WIDTH - 1),
		6041 => to_unsigned(17934, LUT_AMPL_WIDTH - 1),
		6042 => to_unsigned(17937, LUT_AMPL_WIDTH - 1),
		6043 => to_unsigned(17940, LUT_AMPL_WIDTH - 1),
		6044 => to_unsigned(17942, LUT_AMPL_WIDTH - 1),
		6045 => to_unsigned(17945, LUT_AMPL_WIDTH - 1),
		6046 => to_unsigned(17948, LUT_AMPL_WIDTH - 1),
		6047 => to_unsigned(17950, LUT_AMPL_WIDTH - 1),
		6048 => to_unsigned(17953, LUT_AMPL_WIDTH - 1),
		6049 => to_unsigned(17955, LUT_AMPL_WIDTH - 1),
		6050 => to_unsigned(17958, LUT_AMPL_WIDTH - 1),
		6051 => to_unsigned(17961, LUT_AMPL_WIDTH - 1),
		6052 => to_unsigned(17963, LUT_AMPL_WIDTH - 1),
		6053 => to_unsigned(17966, LUT_AMPL_WIDTH - 1),
		6054 => to_unsigned(17969, LUT_AMPL_WIDTH - 1),
		6055 => to_unsigned(17971, LUT_AMPL_WIDTH - 1),
		6056 => to_unsigned(17974, LUT_AMPL_WIDTH - 1),
		6057 => to_unsigned(17976, LUT_AMPL_WIDTH - 1),
		6058 => to_unsigned(17979, LUT_AMPL_WIDTH - 1),
		6059 => to_unsigned(17982, LUT_AMPL_WIDTH - 1),
		6060 => to_unsigned(17984, LUT_AMPL_WIDTH - 1),
		6061 => to_unsigned(17987, LUT_AMPL_WIDTH - 1),
		6062 => to_unsigned(17990, LUT_AMPL_WIDTH - 1),
		6063 => to_unsigned(17992, LUT_AMPL_WIDTH - 1),
		6064 => to_unsigned(17995, LUT_AMPL_WIDTH - 1),
		6065 => to_unsigned(17997, LUT_AMPL_WIDTH - 1),
		6066 => to_unsigned(18000, LUT_AMPL_WIDTH - 1),
		6067 => to_unsigned(18003, LUT_AMPL_WIDTH - 1),
		6068 => to_unsigned(18005, LUT_AMPL_WIDTH - 1),
		6069 => to_unsigned(18008, LUT_AMPL_WIDTH - 1),
		6070 => to_unsigned(18011, LUT_AMPL_WIDTH - 1),
		6071 => to_unsigned(18013, LUT_AMPL_WIDTH - 1),
		6072 => to_unsigned(18016, LUT_AMPL_WIDTH - 1),
		6073 => to_unsigned(18018, LUT_AMPL_WIDTH - 1),
		6074 => to_unsigned(18021, LUT_AMPL_WIDTH - 1),
		6075 => to_unsigned(18024, LUT_AMPL_WIDTH - 1),
		6076 => to_unsigned(18026, LUT_AMPL_WIDTH - 1),
		6077 => to_unsigned(18029, LUT_AMPL_WIDTH - 1),
		6078 => to_unsigned(18032, LUT_AMPL_WIDTH - 1),
		6079 => to_unsigned(18034, LUT_AMPL_WIDTH - 1),
		6080 => to_unsigned(18037, LUT_AMPL_WIDTH - 1),
		6081 => to_unsigned(18039, LUT_AMPL_WIDTH - 1),
		6082 => to_unsigned(18042, LUT_AMPL_WIDTH - 1),
		6083 => to_unsigned(18045, LUT_AMPL_WIDTH - 1),
		6084 => to_unsigned(18047, LUT_AMPL_WIDTH - 1),
		6085 => to_unsigned(18050, LUT_AMPL_WIDTH - 1),
		6086 => to_unsigned(18053, LUT_AMPL_WIDTH - 1),
		6087 => to_unsigned(18055, LUT_AMPL_WIDTH - 1),
		6088 => to_unsigned(18058, LUT_AMPL_WIDTH - 1),
		6089 => to_unsigned(18060, LUT_AMPL_WIDTH - 1),
		6090 => to_unsigned(18063, LUT_AMPL_WIDTH - 1),
		6091 => to_unsigned(18066, LUT_AMPL_WIDTH - 1),
		6092 => to_unsigned(18068, LUT_AMPL_WIDTH - 1),
		6093 => to_unsigned(18071, LUT_AMPL_WIDTH - 1),
		6094 => to_unsigned(18074, LUT_AMPL_WIDTH - 1),
		6095 => to_unsigned(18076, LUT_AMPL_WIDTH - 1),
		6096 => to_unsigned(18079, LUT_AMPL_WIDTH - 1),
		6097 => to_unsigned(18081, LUT_AMPL_WIDTH - 1),
		6098 => to_unsigned(18084, LUT_AMPL_WIDTH - 1),
		6099 => to_unsigned(18087, LUT_AMPL_WIDTH - 1),
		6100 => to_unsigned(18089, LUT_AMPL_WIDTH - 1),
		6101 => to_unsigned(18092, LUT_AMPL_WIDTH - 1),
		6102 => to_unsigned(18095, LUT_AMPL_WIDTH - 1),
		6103 => to_unsigned(18097, LUT_AMPL_WIDTH - 1),
		6104 => to_unsigned(18100, LUT_AMPL_WIDTH - 1),
		6105 => to_unsigned(18102, LUT_AMPL_WIDTH - 1),
		6106 => to_unsigned(18105, LUT_AMPL_WIDTH - 1),
		6107 => to_unsigned(18108, LUT_AMPL_WIDTH - 1),
		6108 => to_unsigned(18110, LUT_AMPL_WIDTH - 1),
		6109 => to_unsigned(18113, LUT_AMPL_WIDTH - 1),
		6110 => to_unsigned(18115, LUT_AMPL_WIDTH - 1),
		6111 => to_unsigned(18118, LUT_AMPL_WIDTH - 1),
		6112 => to_unsigned(18121, LUT_AMPL_WIDTH - 1),
		6113 => to_unsigned(18123, LUT_AMPL_WIDTH - 1),
		6114 => to_unsigned(18126, LUT_AMPL_WIDTH - 1),
		6115 => to_unsigned(18129, LUT_AMPL_WIDTH - 1),
		6116 => to_unsigned(18131, LUT_AMPL_WIDTH - 1),
		6117 => to_unsigned(18134, LUT_AMPL_WIDTH - 1),
		6118 => to_unsigned(18136, LUT_AMPL_WIDTH - 1),
		6119 => to_unsigned(18139, LUT_AMPL_WIDTH - 1),
		6120 => to_unsigned(18142, LUT_AMPL_WIDTH - 1),
		6121 => to_unsigned(18144, LUT_AMPL_WIDTH - 1),
		6122 => to_unsigned(18147, LUT_AMPL_WIDTH - 1),
		6123 => to_unsigned(18149, LUT_AMPL_WIDTH - 1),
		6124 => to_unsigned(18152, LUT_AMPL_WIDTH - 1),
		6125 => to_unsigned(18155, LUT_AMPL_WIDTH - 1),
		6126 => to_unsigned(18157, LUT_AMPL_WIDTH - 1),
		6127 => to_unsigned(18160, LUT_AMPL_WIDTH - 1),
		6128 => to_unsigned(18163, LUT_AMPL_WIDTH - 1),
		6129 => to_unsigned(18165, LUT_AMPL_WIDTH - 1),
		6130 => to_unsigned(18168, LUT_AMPL_WIDTH - 1),
		6131 => to_unsigned(18170, LUT_AMPL_WIDTH - 1),
		6132 => to_unsigned(18173, LUT_AMPL_WIDTH - 1),
		6133 => to_unsigned(18176, LUT_AMPL_WIDTH - 1),
		6134 => to_unsigned(18178, LUT_AMPL_WIDTH - 1),
		6135 => to_unsigned(18181, LUT_AMPL_WIDTH - 1),
		6136 => to_unsigned(18183, LUT_AMPL_WIDTH - 1),
		6137 => to_unsigned(18186, LUT_AMPL_WIDTH - 1),
		6138 => to_unsigned(18189, LUT_AMPL_WIDTH - 1),
		6139 => to_unsigned(18191, LUT_AMPL_WIDTH - 1),
		6140 => to_unsigned(18194, LUT_AMPL_WIDTH - 1),
		6141 => to_unsigned(18197, LUT_AMPL_WIDTH - 1),
		6142 => to_unsigned(18199, LUT_AMPL_WIDTH - 1),
		6143 => to_unsigned(18202, LUT_AMPL_WIDTH - 1),
		6144 => to_unsigned(18204, LUT_AMPL_WIDTH - 1),
		6145 => to_unsigned(18207, LUT_AMPL_WIDTH - 1),
		6146 => to_unsigned(18210, LUT_AMPL_WIDTH - 1),
		6147 => to_unsigned(18212, LUT_AMPL_WIDTH - 1),
		6148 => to_unsigned(18215, LUT_AMPL_WIDTH - 1),
		6149 => to_unsigned(18217, LUT_AMPL_WIDTH - 1),
		6150 => to_unsigned(18220, LUT_AMPL_WIDTH - 1),
		6151 => to_unsigned(18223, LUT_AMPL_WIDTH - 1),
		6152 => to_unsigned(18225, LUT_AMPL_WIDTH - 1),
		6153 => to_unsigned(18228, LUT_AMPL_WIDTH - 1),
		6154 => to_unsigned(18230, LUT_AMPL_WIDTH - 1),
		6155 => to_unsigned(18233, LUT_AMPL_WIDTH - 1),
		6156 => to_unsigned(18236, LUT_AMPL_WIDTH - 1),
		6157 => to_unsigned(18238, LUT_AMPL_WIDTH - 1),
		6158 => to_unsigned(18241, LUT_AMPL_WIDTH - 1),
		6159 => to_unsigned(18244, LUT_AMPL_WIDTH - 1),
		6160 => to_unsigned(18246, LUT_AMPL_WIDTH - 1),
		6161 => to_unsigned(18249, LUT_AMPL_WIDTH - 1),
		6162 => to_unsigned(18251, LUT_AMPL_WIDTH - 1),
		6163 => to_unsigned(18254, LUT_AMPL_WIDTH - 1),
		6164 => to_unsigned(18257, LUT_AMPL_WIDTH - 1),
		6165 => to_unsigned(18259, LUT_AMPL_WIDTH - 1),
		6166 => to_unsigned(18262, LUT_AMPL_WIDTH - 1),
		6167 => to_unsigned(18264, LUT_AMPL_WIDTH - 1),
		6168 => to_unsigned(18267, LUT_AMPL_WIDTH - 1),
		6169 => to_unsigned(18270, LUT_AMPL_WIDTH - 1),
		6170 => to_unsigned(18272, LUT_AMPL_WIDTH - 1),
		6171 => to_unsigned(18275, LUT_AMPL_WIDTH - 1),
		6172 => to_unsigned(18277, LUT_AMPL_WIDTH - 1),
		6173 => to_unsigned(18280, LUT_AMPL_WIDTH - 1),
		6174 => to_unsigned(18283, LUT_AMPL_WIDTH - 1),
		6175 => to_unsigned(18285, LUT_AMPL_WIDTH - 1),
		6176 => to_unsigned(18288, LUT_AMPL_WIDTH - 1),
		6177 => to_unsigned(18290, LUT_AMPL_WIDTH - 1),
		6178 => to_unsigned(18293, LUT_AMPL_WIDTH - 1),
		6179 => to_unsigned(18296, LUT_AMPL_WIDTH - 1),
		6180 => to_unsigned(18298, LUT_AMPL_WIDTH - 1),
		6181 => to_unsigned(18301, LUT_AMPL_WIDTH - 1),
		6182 => to_unsigned(18304, LUT_AMPL_WIDTH - 1),
		6183 => to_unsigned(18306, LUT_AMPL_WIDTH - 1),
		6184 => to_unsigned(18309, LUT_AMPL_WIDTH - 1),
		6185 => to_unsigned(18311, LUT_AMPL_WIDTH - 1),
		6186 => to_unsigned(18314, LUT_AMPL_WIDTH - 1),
		6187 => to_unsigned(18317, LUT_AMPL_WIDTH - 1),
		6188 => to_unsigned(18319, LUT_AMPL_WIDTH - 1),
		6189 => to_unsigned(18322, LUT_AMPL_WIDTH - 1),
		6190 => to_unsigned(18324, LUT_AMPL_WIDTH - 1),
		6191 => to_unsigned(18327, LUT_AMPL_WIDTH - 1),
		6192 => to_unsigned(18330, LUT_AMPL_WIDTH - 1),
		6193 => to_unsigned(18332, LUT_AMPL_WIDTH - 1),
		6194 => to_unsigned(18335, LUT_AMPL_WIDTH - 1),
		6195 => to_unsigned(18337, LUT_AMPL_WIDTH - 1),
		6196 => to_unsigned(18340, LUT_AMPL_WIDTH - 1),
		6197 => to_unsigned(18343, LUT_AMPL_WIDTH - 1),
		6198 => to_unsigned(18345, LUT_AMPL_WIDTH - 1),
		6199 => to_unsigned(18348, LUT_AMPL_WIDTH - 1),
		6200 => to_unsigned(18350, LUT_AMPL_WIDTH - 1),
		6201 => to_unsigned(18353, LUT_AMPL_WIDTH - 1),
		6202 => to_unsigned(18356, LUT_AMPL_WIDTH - 1),
		6203 => to_unsigned(18358, LUT_AMPL_WIDTH - 1),
		6204 => to_unsigned(18361, LUT_AMPL_WIDTH - 1),
		6205 => to_unsigned(18363, LUT_AMPL_WIDTH - 1),
		6206 => to_unsigned(18366, LUT_AMPL_WIDTH - 1),
		6207 => to_unsigned(18369, LUT_AMPL_WIDTH - 1),
		6208 => to_unsigned(18371, LUT_AMPL_WIDTH - 1),
		6209 => to_unsigned(18374, LUT_AMPL_WIDTH - 1),
		6210 => to_unsigned(18376, LUT_AMPL_WIDTH - 1),
		6211 => to_unsigned(18379, LUT_AMPL_WIDTH - 1),
		6212 => to_unsigned(18382, LUT_AMPL_WIDTH - 1),
		6213 => to_unsigned(18384, LUT_AMPL_WIDTH - 1),
		6214 => to_unsigned(18387, LUT_AMPL_WIDTH - 1),
		6215 => to_unsigned(18389, LUT_AMPL_WIDTH - 1),
		6216 => to_unsigned(18392, LUT_AMPL_WIDTH - 1),
		6217 => to_unsigned(18395, LUT_AMPL_WIDTH - 1),
		6218 => to_unsigned(18397, LUT_AMPL_WIDTH - 1),
		6219 => to_unsigned(18400, LUT_AMPL_WIDTH - 1),
		6220 => to_unsigned(18402, LUT_AMPL_WIDTH - 1),
		6221 => to_unsigned(18405, LUT_AMPL_WIDTH - 1),
		6222 => to_unsigned(18408, LUT_AMPL_WIDTH - 1),
		6223 => to_unsigned(18410, LUT_AMPL_WIDTH - 1),
		6224 => to_unsigned(18413, LUT_AMPL_WIDTH - 1),
		6225 => to_unsigned(18415, LUT_AMPL_WIDTH - 1),
		6226 => to_unsigned(18418, LUT_AMPL_WIDTH - 1),
		6227 => to_unsigned(18421, LUT_AMPL_WIDTH - 1),
		6228 => to_unsigned(18423, LUT_AMPL_WIDTH - 1),
		6229 => to_unsigned(18426, LUT_AMPL_WIDTH - 1),
		6230 => to_unsigned(18428, LUT_AMPL_WIDTH - 1),
		6231 => to_unsigned(18431, LUT_AMPL_WIDTH - 1),
		6232 => to_unsigned(18434, LUT_AMPL_WIDTH - 1),
		6233 => to_unsigned(18436, LUT_AMPL_WIDTH - 1),
		6234 => to_unsigned(18439, LUT_AMPL_WIDTH - 1),
		6235 => to_unsigned(18441, LUT_AMPL_WIDTH - 1),
		6236 => to_unsigned(18444, LUT_AMPL_WIDTH - 1),
		6237 => to_unsigned(18447, LUT_AMPL_WIDTH - 1),
		6238 => to_unsigned(18449, LUT_AMPL_WIDTH - 1),
		6239 => to_unsigned(18452, LUT_AMPL_WIDTH - 1),
		6240 => to_unsigned(18454, LUT_AMPL_WIDTH - 1),
		6241 => to_unsigned(18457, LUT_AMPL_WIDTH - 1),
		6242 => to_unsigned(18460, LUT_AMPL_WIDTH - 1),
		6243 => to_unsigned(18462, LUT_AMPL_WIDTH - 1),
		6244 => to_unsigned(18465, LUT_AMPL_WIDTH - 1),
		6245 => to_unsigned(18467, LUT_AMPL_WIDTH - 1),
		6246 => to_unsigned(18470, LUT_AMPL_WIDTH - 1),
		6247 => to_unsigned(18473, LUT_AMPL_WIDTH - 1),
		6248 => to_unsigned(18475, LUT_AMPL_WIDTH - 1),
		6249 => to_unsigned(18478, LUT_AMPL_WIDTH - 1),
		6250 => to_unsigned(18480, LUT_AMPL_WIDTH - 1),
		6251 => to_unsigned(18483, LUT_AMPL_WIDTH - 1),
		6252 => to_unsigned(18485, LUT_AMPL_WIDTH - 1),
		6253 => to_unsigned(18488, LUT_AMPL_WIDTH - 1),
		6254 => to_unsigned(18491, LUT_AMPL_WIDTH - 1),
		6255 => to_unsigned(18493, LUT_AMPL_WIDTH - 1),
		6256 => to_unsigned(18496, LUT_AMPL_WIDTH - 1),
		6257 => to_unsigned(18498, LUT_AMPL_WIDTH - 1),
		6258 => to_unsigned(18501, LUT_AMPL_WIDTH - 1),
		6259 => to_unsigned(18504, LUT_AMPL_WIDTH - 1),
		6260 => to_unsigned(18506, LUT_AMPL_WIDTH - 1),
		6261 => to_unsigned(18509, LUT_AMPL_WIDTH - 1),
		6262 => to_unsigned(18511, LUT_AMPL_WIDTH - 1),
		6263 => to_unsigned(18514, LUT_AMPL_WIDTH - 1),
		6264 => to_unsigned(18517, LUT_AMPL_WIDTH - 1),
		6265 => to_unsigned(18519, LUT_AMPL_WIDTH - 1),
		6266 => to_unsigned(18522, LUT_AMPL_WIDTH - 1),
		6267 => to_unsigned(18524, LUT_AMPL_WIDTH - 1),
		6268 => to_unsigned(18527, LUT_AMPL_WIDTH - 1),
		6269 => to_unsigned(18530, LUT_AMPL_WIDTH - 1),
		6270 => to_unsigned(18532, LUT_AMPL_WIDTH - 1),
		6271 => to_unsigned(18535, LUT_AMPL_WIDTH - 1),
		6272 => to_unsigned(18537, LUT_AMPL_WIDTH - 1),
		6273 => to_unsigned(18540, LUT_AMPL_WIDTH - 1),
		6274 => to_unsigned(18543, LUT_AMPL_WIDTH - 1),
		6275 => to_unsigned(18545, LUT_AMPL_WIDTH - 1),
		6276 => to_unsigned(18548, LUT_AMPL_WIDTH - 1),
		6277 => to_unsigned(18550, LUT_AMPL_WIDTH - 1),
		6278 => to_unsigned(18553, LUT_AMPL_WIDTH - 1),
		6279 => to_unsigned(18555, LUT_AMPL_WIDTH - 1),
		6280 => to_unsigned(18558, LUT_AMPL_WIDTH - 1),
		6281 => to_unsigned(18561, LUT_AMPL_WIDTH - 1),
		6282 => to_unsigned(18563, LUT_AMPL_WIDTH - 1),
		6283 => to_unsigned(18566, LUT_AMPL_WIDTH - 1),
		6284 => to_unsigned(18568, LUT_AMPL_WIDTH - 1),
		6285 => to_unsigned(18571, LUT_AMPL_WIDTH - 1),
		6286 => to_unsigned(18574, LUT_AMPL_WIDTH - 1),
		6287 => to_unsigned(18576, LUT_AMPL_WIDTH - 1),
		6288 => to_unsigned(18579, LUT_AMPL_WIDTH - 1),
		6289 => to_unsigned(18581, LUT_AMPL_WIDTH - 1),
		6290 => to_unsigned(18584, LUT_AMPL_WIDTH - 1),
		6291 => to_unsigned(18587, LUT_AMPL_WIDTH - 1),
		6292 => to_unsigned(18589, LUT_AMPL_WIDTH - 1),
		6293 => to_unsigned(18592, LUT_AMPL_WIDTH - 1),
		6294 => to_unsigned(18594, LUT_AMPL_WIDTH - 1),
		6295 => to_unsigned(18597, LUT_AMPL_WIDTH - 1),
		6296 => to_unsigned(18599, LUT_AMPL_WIDTH - 1),
		6297 => to_unsigned(18602, LUT_AMPL_WIDTH - 1),
		6298 => to_unsigned(18605, LUT_AMPL_WIDTH - 1),
		6299 => to_unsigned(18607, LUT_AMPL_WIDTH - 1),
		6300 => to_unsigned(18610, LUT_AMPL_WIDTH - 1),
		6301 => to_unsigned(18612, LUT_AMPL_WIDTH - 1),
		6302 => to_unsigned(18615, LUT_AMPL_WIDTH - 1),
		6303 => to_unsigned(18618, LUT_AMPL_WIDTH - 1),
		6304 => to_unsigned(18620, LUT_AMPL_WIDTH - 1),
		6305 => to_unsigned(18623, LUT_AMPL_WIDTH - 1),
		6306 => to_unsigned(18625, LUT_AMPL_WIDTH - 1),
		6307 => to_unsigned(18628, LUT_AMPL_WIDTH - 1),
		6308 => to_unsigned(18630, LUT_AMPL_WIDTH - 1),
		6309 => to_unsigned(18633, LUT_AMPL_WIDTH - 1),
		6310 => to_unsigned(18636, LUT_AMPL_WIDTH - 1),
		6311 => to_unsigned(18638, LUT_AMPL_WIDTH - 1),
		6312 => to_unsigned(18641, LUT_AMPL_WIDTH - 1),
		6313 => to_unsigned(18643, LUT_AMPL_WIDTH - 1),
		6314 => to_unsigned(18646, LUT_AMPL_WIDTH - 1),
		6315 => to_unsigned(18649, LUT_AMPL_WIDTH - 1),
		6316 => to_unsigned(18651, LUT_AMPL_WIDTH - 1),
		6317 => to_unsigned(18654, LUT_AMPL_WIDTH - 1),
		6318 => to_unsigned(18656, LUT_AMPL_WIDTH - 1),
		6319 => to_unsigned(18659, LUT_AMPL_WIDTH - 1),
		6320 => to_unsigned(18661, LUT_AMPL_WIDTH - 1),
		6321 => to_unsigned(18664, LUT_AMPL_WIDTH - 1),
		6322 => to_unsigned(18667, LUT_AMPL_WIDTH - 1),
		6323 => to_unsigned(18669, LUT_AMPL_WIDTH - 1),
		6324 => to_unsigned(18672, LUT_AMPL_WIDTH - 1),
		6325 => to_unsigned(18674, LUT_AMPL_WIDTH - 1),
		6326 => to_unsigned(18677, LUT_AMPL_WIDTH - 1),
		6327 => to_unsigned(18680, LUT_AMPL_WIDTH - 1),
		6328 => to_unsigned(18682, LUT_AMPL_WIDTH - 1),
		6329 => to_unsigned(18685, LUT_AMPL_WIDTH - 1),
		6330 => to_unsigned(18687, LUT_AMPL_WIDTH - 1),
		6331 => to_unsigned(18690, LUT_AMPL_WIDTH - 1),
		6332 => to_unsigned(18692, LUT_AMPL_WIDTH - 1),
		6333 => to_unsigned(18695, LUT_AMPL_WIDTH - 1),
		6334 => to_unsigned(18698, LUT_AMPL_WIDTH - 1),
		6335 => to_unsigned(18700, LUT_AMPL_WIDTH - 1),
		6336 => to_unsigned(18703, LUT_AMPL_WIDTH - 1),
		6337 => to_unsigned(18705, LUT_AMPL_WIDTH - 1),
		6338 => to_unsigned(18708, LUT_AMPL_WIDTH - 1),
		6339 => to_unsigned(18711, LUT_AMPL_WIDTH - 1),
		6340 => to_unsigned(18713, LUT_AMPL_WIDTH - 1),
		6341 => to_unsigned(18716, LUT_AMPL_WIDTH - 1),
		6342 => to_unsigned(18718, LUT_AMPL_WIDTH - 1),
		6343 => to_unsigned(18721, LUT_AMPL_WIDTH - 1),
		6344 => to_unsigned(18723, LUT_AMPL_WIDTH - 1),
		6345 => to_unsigned(18726, LUT_AMPL_WIDTH - 1),
		6346 => to_unsigned(18729, LUT_AMPL_WIDTH - 1),
		6347 => to_unsigned(18731, LUT_AMPL_WIDTH - 1),
		6348 => to_unsigned(18734, LUT_AMPL_WIDTH - 1),
		6349 => to_unsigned(18736, LUT_AMPL_WIDTH - 1),
		6350 => to_unsigned(18739, LUT_AMPL_WIDTH - 1),
		6351 => to_unsigned(18741, LUT_AMPL_WIDTH - 1),
		6352 => to_unsigned(18744, LUT_AMPL_WIDTH - 1),
		6353 => to_unsigned(18747, LUT_AMPL_WIDTH - 1),
		6354 => to_unsigned(18749, LUT_AMPL_WIDTH - 1),
		6355 => to_unsigned(18752, LUT_AMPL_WIDTH - 1),
		6356 => to_unsigned(18754, LUT_AMPL_WIDTH - 1),
		6357 => to_unsigned(18757, LUT_AMPL_WIDTH - 1),
		6358 => to_unsigned(18759, LUT_AMPL_WIDTH - 1),
		6359 => to_unsigned(18762, LUT_AMPL_WIDTH - 1),
		6360 => to_unsigned(18765, LUT_AMPL_WIDTH - 1),
		6361 => to_unsigned(18767, LUT_AMPL_WIDTH - 1),
		6362 => to_unsigned(18770, LUT_AMPL_WIDTH - 1),
		6363 => to_unsigned(18772, LUT_AMPL_WIDTH - 1),
		6364 => to_unsigned(18775, LUT_AMPL_WIDTH - 1),
		6365 => to_unsigned(18778, LUT_AMPL_WIDTH - 1),
		6366 => to_unsigned(18780, LUT_AMPL_WIDTH - 1),
		6367 => to_unsigned(18783, LUT_AMPL_WIDTH - 1),
		6368 => to_unsigned(18785, LUT_AMPL_WIDTH - 1),
		6369 => to_unsigned(18788, LUT_AMPL_WIDTH - 1),
		6370 => to_unsigned(18790, LUT_AMPL_WIDTH - 1),
		6371 => to_unsigned(18793, LUT_AMPL_WIDTH - 1),
		6372 => to_unsigned(18796, LUT_AMPL_WIDTH - 1),
		6373 => to_unsigned(18798, LUT_AMPL_WIDTH - 1),
		6374 => to_unsigned(18801, LUT_AMPL_WIDTH - 1),
		6375 => to_unsigned(18803, LUT_AMPL_WIDTH - 1),
		6376 => to_unsigned(18806, LUT_AMPL_WIDTH - 1),
		6377 => to_unsigned(18808, LUT_AMPL_WIDTH - 1),
		6378 => to_unsigned(18811, LUT_AMPL_WIDTH - 1),
		6379 => to_unsigned(18814, LUT_AMPL_WIDTH - 1),
		6380 => to_unsigned(18816, LUT_AMPL_WIDTH - 1),
		6381 => to_unsigned(18819, LUT_AMPL_WIDTH - 1),
		6382 => to_unsigned(18821, LUT_AMPL_WIDTH - 1),
		6383 => to_unsigned(18824, LUT_AMPL_WIDTH - 1),
		6384 => to_unsigned(18826, LUT_AMPL_WIDTH - 1),
		6385 => to_unsigned(18829, LUT_AMPL_WIDTH - 1),
		6386 => to_unsigned(18832, LUT_AMPL_WIDTH - 1),
		6387 => to_unsigned(18834, LUT_AMPL_WIDTH - 1),
		6388 => to_unsigned(18837, LUT_AMPL_WIDTH - 1),
		6389 => to_unsigned(18839, LUT_AMPL_WIDTH - 1),
		6390 => to_unsigned(18842, LUT_AMPL_WIDTH - 1),
		6391 => to_unsigned(18844, LUT_AMPL_WIDTH - 1),
		6392 => to_unsigned(18847, LUT_AMPL_WIDTH - 1),
		6393 => to_unsigned(18850, LUT_AMPL_WIDTH - 1),
		6394 => to_unsigned(18852, LUT_AMPL_WIDTH - 1),
		6395 => to_unsigned(18855, LUT_AMPL_WIDTH - 1),
		6396 => to_unsigned(18857, LUT_AMPL_WIDTH - 1),
		6397 => to_unsigned(18860, LUT_AMPL_WIDTH - 1),
		6398 => to_unsigned(18862, LUT_AMPL_WIDTH - 1),
		6399 => to_unsigned(18865, LUT_AMPL_WIDTH - 1),
		6400 => to_unsigned(18868, LUT_AMPL_WIDTH - 1),
		6401 => to_unsigned(18870, LUT_AMPL_WIDTH - 1),
		6402 => to_unsigned(18873, LUT_AMPL_WIDTH - 1),
		6403 => to_unsigned(18875, LUT_AMPL_WIDTH - 1),
		6404 => to_unsigned(18878, LUT_AMPL_WIDTH - 1),
		6405 => to_unsigned(18880, LUT_AMPL_WIDTH - 1),
		6406 => to_unsigned(18883, LUT_AMPL_WIDTH - 1),
		6407 => to_unsigned(18885, LUT_AMPL_WIDTH - 1),
		6408 => to_unsigned(18888, LUT_AMPL_WIDTH - 1),
		6409 => to_unsigned(18891, LUT_AMPL_WIDTH - 1),
		6410 => to_unsigned(18893, LUT_AMPL_WIDTH - 1),
		6411 => to_unsigned(18896, LUT_AMPL_WIDTH - 1),
		6412 => to_unsigned(18898, LUT_AMPL_WIDTH - 1),
		6413 => to_unsigned(18901, LUT_AMPL_WIDTH - 1),
		6414 => to_unsigned(18903, LUT_AMPL_WIDTH - 1),
		6415 => to_unsigned(18906, LUT_AMPL_WIDTH - 1),
		6416 => to_unsigned(18909, LUT_AMPL_WIDTH - 1),
		6417 => to_unsigned(18911, LUT_AMPL_WIDTH - 1),
		6418 => to_unsigned(18914, LUT_AMPL_WIDTH - 1),
		6419 => to_unsigned(18916, LUT_AMPL_WIDTH - 1),
		6420 => to_unsigned(18919, LUT_AMPL_WIDTH - 1),
		6421 => to_unsigned(18921, LUT_AMPL_WIDTH - 1),
		6422 => to_unsigned(18924, LUT_AMPL_WIDTH - 1),
		6423 => to_unsigned(18927, LUT_AMPL_WIDTH - 1),
		6424 => to_unsigned(18929, LUT_AMPL_WIDTH - 1),
		6425 => to_unsigned(18932, LUT_AMPL_WIDTH - 1),
		6426 => to_unsigned(18934, LUT_AMPL_WIDTH - 1),
		6427 => to_unsigned(18937, LUT_AMPL_WIDTH - 1),
		6428 => to_unsigned(18939, LUT_AMPL_WIDTH - 1),
		6429 => to_unsigned(18942, LUT_AMPL_WIDTH - 1),
		6430 => to_unsigned(18944, LUT_AMPL_WIDTH - 1),
		6431 => to_unsigned(18947, LUT_AMPL_WIDTH - 1),
		6432 => to_unsigned(18950, LUT_AMPL_WIDTH - 1),
		6433 => to_unsigned(18952, LUT_AMPL_WIDTH - 1),
		6434 => to_unsigned(18955, LUT_AMPL_WIDTH - 1),
		6435 => to_unsigned(18957, LUT_AMPL_WIDTH - 1),
		6436 => to_unsigned(18960, LUT_AMPL_WIDTH - 1),
		6437 => to_unsigned(18962, LUT_AMPL_WIDTH - 1),
		6438 => to_unsigned(18965, LUT_AMPL_WIDTH - 1),
		6439 => to_unsigned(18968, LUT_AMPL_WIDTH - 1),
		6440 => to_unsigned(18970, LUT_AMPL_WIDTH - 1),
		6441 => to_unsigned(18973, LUT_AMPL_WIDTH - 1),
		6442 => to_unsigned(18975, LUT_AMPL_WIDTH - 1),
		6443 => to_unsigned(18978, LUT_AMPL_WIDTH - 1),
		6444 => to_unsigned(18980, LUT_AMPL_WIDTH - 1),
		6445 => to_unsigned(18983, LUT_AMPL_WIDTH - 1),
		6446 => to_unsigned(18985, LUT_AMPL_WIDTH - 1),
		6447 => to_unsigned(18988, LUT_AMPL_WIDTH - 1),
		6448 => to_unsigned(18991, LUT_AMPL_WIDTH - 1),
		6449 => to_unsigned(18993, LUT_AMPL_WIDTH - 1),
		6450 => to_unsigned(18996, LUT_AMPL_WIDTH - 1),
		6451 => to_unsigned(18998, LUT_AMPL_WIDTH - 1),
		6452 => to_unsigned(19001, LUT_AMPL_WIDTH - 1),
		6453 => to_unsigned(19003, LUT_AMPL_WIDTH - 1),
		6454 => to_unsigned(19006, LUT_AMPL_WIDTH - 1),
		6455 => to_unsigned(19009, LUT_AMPL_WIDTH - 1),
		6456 => to_unsigned(19011, LUT_AMPL_WIDTH - 1),
		6457 => to_unsigned(19014, LUT_AMPL_WIDTH - 1),
		6458 => to_unsigned(19016, LUT_AMPL_WIDTH - 1),
		6459 => to_unsigned(19019, LUT_AMPL_WIDTH - 1),
		6460 => to_unsigned(19021, LUT_AMPL_WIDTH - 1),
		6461 => to_unsigned(19024, LUT_AMPL_WIDTH - 1),
		6462 => to_unsigned(19026, LUT_AMPL_WIDTH - 1),
		6463 => to_unsigned(19029, LUT_AMPL_WIDTH - 1),
		6464 => to_unsigned(19032, LUT_AMPL_WIDTH - 1),
		6465 => to_unsigned(19034, LUT_AMPL_WIDTH - 1),
		6466 => to_unsigned(19037, LUT_AMPL_WIDTH - 1),
		6467 => to_unsigned(19039, LUT_AMPL_WIDTH - 1),
		6468 => to_unsigned(19042, LUT_AMPL_WIDTH - 1),
		6469 => to_unsigned(19044, LUT_AMPL_WIDTH - 1),
		6470 => to_unsigned(19047, LUT_AMPL_WIDTH - 1),
		6471 => to_unsigned(19049, LUT_AMPL_WIDTH - 1),
		6472 => to_unsigned(19052, LUT_AMPL_WIDTH - 1),
		6473 => to_unsigned(19055, LUT_AMPL_WIDTH - 1),
		6474 => to_unsigned(19057, LUT_AMPL_WIDTH - 1),
		6475 => to_unsigned(19060, LUT_AMPL_WIDTH - 1),
		6476 => to_unsigned(19062, LUT_AMPL_WIDTH - 1),
		6477 => to_unsigned(19065, LUT_AMPL_WIDTH - 1),
		6478 => to_unsigned(19067, LUT_AMPL_WIDTH - 1),
		6479 => to_unsigned(19070, LUT_AMPL_WIDTH - 1),
		6480 => to_unsigned(19072, LUT_AMPL_WIDTH - 1),
		6481 => to_unsigned(19075, LUT_AMPL_WIDTH - 1),
		6482 => to_unsigned(19078, LUT_AMPL_WIDTH - 1),
		6483 => to_unsigned(19080, LUT_AMPL_WIDTH - 1),
		6484 => to_unsigned(19083, LUT_AMPL_WIDTH - 1),
		6485 => to_unsigned(19085, LUT_AMPL_WIDTH - 1),
		6486 => to_unsigned(19088, LUT_AMPL_WIDTH - 1),
		6487 => to_unsigned(19090, LUT_AMPL_WIDTH - 1),
		6488 => to_unsigned(19093, LUT_AMPL_WIDTH - 1),
		6489 => to_unsigned(19095, LUT_AMPL_WIDTH - 1),
		6490 => to_unsigned(19098, LUT_AMPL_WIDTH - 1),
		6491 => to_unsigned(19101, LUT_AMPL_WIDTH - 1),
		6492 => to_unsigned(19103, LUT_AMPL_WIDTH - 1),
		6493 => to_unsigned(19106, LUT_AMPL_WIDTH - 1),
		6494 => to_unsigned(19108, LUT_AMPL_WIDTH - 1),
		6495 => to_unsigned(19111, LUT_AMPL_WIDTH - 1),
		6496 => to_unsigned(19113, LUT_AMPL_WIDTH - 1),
		6497 => to_unsigned(19116, LUT_AMPL_WIDTH - 1),
		6498 => to_unsigned(19118, LUT_AMPL_WIDTH - 1),
		6499 => to_unsigned(19121, LUT_AMPL_WIDTH - 1),
		6500 => to_unsigned(19123, LUT_AMPL_WIDTH - 1),
		6501 => to_unsigned(19126, LUT_AMPL_WIDTH - 1),
		6502 => to_unsigned(19129, LUT_AMPL_WIDTH - 1),
		6503 => to_unsigned(19131, LUT_AMPL_WIDTH - 1),
		6504 => to_unsigned(19134, LUT_AMPL_WIDTH - 1),
		6505 => to_unsigned(19136, LUT_AMPL_WIDTH - 1),
		6506 => to_unsigned(19139, LUT_AMPL_WIDTH - 1),
		6507 => to_unsigned(19141, LUT_AMPL_WIDTH - 1),
		6508 => to_unsigned(19144, LUT_AMPL_WIDTH - 1),
		6509 => to_unsigned(19146, LUT_AMPL_WIDTH - 1),
		6510 => to_unsigned(19149, LUT_AMPL_WIDTH - 1),
		6511 => to_unsigned(19152, LUT_AMPL_WIDTH - 1),
		6512 => to_unsigned(19154, LUT_AMPL_WIDTH - 1),
		6513 => to_unsigned(19157, LUT_AMPL_WIDTH - 1),
		6514 => to_unsigned(19159, LUT_AMPL_WIDTH - 1),
		6515 => to_unsigned(19162, LUT_AMPL_WIDTH - 1),
		6516 => to_unsigned(19164, LUT_AMPL_WIDTH - 1),
		6517 => to_unsigned(19167, LUT_AMPL_WIDTH - 1),
		6518 => to_unsigned(19169, LUT_AMPL_WIDTH - 1),
		6519 => to_unsigned(19172, LUT_AMPL_WIDTH - 1),
		6520 => to_unsigned(19174, LUT_AMPL_WIDTH - 1),
		6521 => to_unsigned(19177, LUT_AMPL_WIDTH - 1),
		6522 => to_unsigned(19180, LUT_AMPL_WIDTH - 1),
		6523 => to_unsigned(19182, LUT_AMPL_WIDTH - 1),
		6524 => to_unsigned(19185, LUT_AMPL_WIDTH - 1),
		6525 => to_unsigned(19187, LUT_AMPL_WIDTH - 1),
		6526 => to_unsigned(19190, LUT_AMPL_WIDTH - 1),
		6527 => to_unsigned(19192, LUT_AMPL_WIDTH - 1),
		6528 => to_unsigned(19195, LUT_AMPL_WIDTH - 1),
		6529 => to_unsigned(19197, LUT_AMPL_WIDTH - 1),
		6530 => to_unsigned(19200, LUT_AMPL_WIDTH - 1),
		6531 => to_unsigned(19202, LUT_AMPL_WIDTH - 1),
		6532 => to_unsigned(19205, LUT_AMPL_WIDTH - 1),
		6533 => to_unsigned(19208, LUT_AMPL_WIDTH - 1),
		6534 => to_unsigned(19210, LUT_AMPL_WIDTH - 1),
		6535 => to_unsigned(19213, LUT_AMPL_WIDTH - 1),
		6536 => to_unsigned(19215, LUT_AMPL_WIDTH - 1),
		6537 => to_unsigned(19218, LUT_AMPL_WIDTH - 1),
		6538 => to_unsigned(19220, LUT_AMPL_WIDTH - 1),
		6539 => to_unsigned(19223, LUT_AMPL_WIDTH - 1),
		6540 => to_unsigned(19225, LUT_AMPL_WIDTH - 1),
		6541 => to_unsigned(19228, LUT_AMPL_WIDTH - 1),
		6542 => to_unsigned(19230, LUT_AMPL_WIDTH - 1),
		6543 => to_unsigned(19233, LUT_AMPL_WIDTH - 1),
		6544 => to_unsigned(19236, LUT_AMPL_WIDTH - 1),
		6545 => to_unsigned(19238, LUT_AMPL_WIDTH - 1),
		6546 => to_unsigned(19241, LUT_AMPL_WIDTH - 1),
		6547 => to_unsigned(19243, LUT_AMPL_WIDTH - 1),
		6548 => to_unsigned(19246, LUT_AMPL_WIDTH - 1),
		6549 => to_unsigned(19248, LUT_AMPL_WIDTH - 1),
		6550 => to_unsigned(19251, LUT_AMPL_WIDTH - 1),
		6551 => to_unsigned(19253, LUT_AMPL_WIDTH - 1),
		6552 => to_unsigned(19256, LUT_AMPL_WIDTH - 1),
		6553 => to_unsigned(19258, LUT_AMPL_WIDTH - 1),
		6554 => to_unsigned(19261, LUT_AMPL_WIDTH - 1),
		6555 => to_unsigned(19264, LUT_AMPL_WIDTH - 1),
		6556 => to_unsigned(19266, LUT_AMPL_WIDTH - 1),
		6557 => to_unsigned(19269, LUT_AMPL_WIDTH - 1),
		6558 => to_unsigned(19271, LUT_AMPL_WIDTH - 1),
		6559 => to_unsigned(19274, LUT_AMPL_WIDTH - 1),
		6560 => to_unsigned(19276, LUT_AMPL_WIDTH - 1),
		6561 => to_unsigned(19279, LUT_AMPL_WIDTH - 1),
		6562 => to_unsigned(19281, LUT_AMPL_WIDTH - 1),
		6563 => to_unsigned(19284, LUT_AMPL_WIDTH - 1),
		6564 => to_unsigned(19286, LUT_AMPL_WIDTH - 1),
		6565 => to_unsigned(19289, LUT_AMPL_WIDTH - 1),
		6566 => to_unsigned(19291, LUT_AMPL_WIDTH - 1),
		6567 => to_unsigned(19294, LUT_AMPL_WIDTH - 1),
		6568 => to_unsigned(19297, LUT_AMPL_WIDTH - 1),
		6569 => to_unsigned(19299, LUT_AMPL_WIDTH - 1),
		6570 => to_unsigned(19302, LUT_AMPL_WIDTH - 1),
		6571 => to_unsigned(19304, LUT_AMPL_WIDTH - 1),
		6572 => to_unsigned(19307, LUT_AMPL_WIDTH - 1),
		6573 => to_unsigned(19309, LUT_AMPL_WIDTH - 1),
		6574 => to_unsigned(19312, LUT_AMPL_WIDTH - 1),
		6575 => to_unsigned(19314, LUT_AMPL_WIDTH - 1),
		6576 => to_unsigned(19317, LUT_AMPL_WIDTH - 1),
		6577 => to_unsigned(19319, LUT_AMPL_WIDTH - 1),
		6578 => to_unsigned(19322, LUT_AMPL_WIDTH - 1),
		6579 => to_unsigned(19324, LUT_AMPL_WIDTH - 1),
		6580 => to_unsigned(19327, LUT_AMPL_WIDTH - 1),
		6581 => to_unsigned(19330, LUT_AMPL_WIDTH - 1),
		6582 => to_unsigned(19332, LUT_AMPL_WIDTH - 1),
		6583 => to_unsigned(19335, LUT_AMPL_WIDTH - 1),
		6584 => to_unsigned(19337, LUT_AMPL_WIDTH - 1),
		6585 => to_unsigned(19340, LUT_AMPL_WIDTH - 1),
		6586 => to_unsigned(19342, LUT_AMPL_WIDTH - 1),
		6587 => to_unsigned(19345, LUT_AMPL_WIDTH - 1),
		6588 => to_unsigned(19347, LUT_AMPL_WIDTH - 1),
		6589 => to_unsigned(19350, LUT_AMPL_WIDTH - 1),
		6590 => to_unsigned(19352, LUT_AMPL_WIDTH - 1),
		6591 => to_unsigned(19355, LUT_AMPL_WIDTH - 1),
		6592 => to_unsigned(19357, LUT_AMPL_WIDTH - 1),
		6593 => to_unsigned(19360, LUT_AMPL_WIDTH - 1),
		6594 => to_unsigned(19362, LUT_AMPL_WIDTH - 1),
		6595 => to_unsigned(19365, LUT_AMPL_WIDTH - 1),
		6596 => to_unsigned(19368, LUT_AMPL_WIDTH - 1),
		6597 => to_unsigned(19370, LUT_AMPL_WIDTH - 1),
		6598 => to_unsigned(19373, LUT_AMPL_WIDTH - 1),
		6599 => to_unsigned(19375, LUT_AMPL_WIDTH - 1),
		6600 => to_unsigned(19378, LUT_AMPL_WIDTH - 1),
		6601 => to_unsigned(19380, LUT_AMPL_WIDTH - 1),
		6602 => to_unsigned(19383, LUT_AMPL_WIDTH - 1),
		6603 => to_unsigned(19385, LUT_AMPL_WIDTH - 1),
		6604 => to_unsigned(19388, LUT_AMPL_WIDTH - 1),
		6605 => to_unsigned(19390, LUT_AMPL_WIDTH - 1),
		6606 => to_unsigned(19393, LUT_AMPL_WIDTH - 1),
		6607 => to_unsigned(19395, LUT_AMPL_WIDTH - 1),
		6608 => to_unsigned(19398, LUT_AMPL_WIDTH - 1),
		6609 => to_unsigned(19400, LUT_AMPL_WIDTH - 1),
		6610 => to_unsigned(19403, LUT_AMPL_WIDTH - 1),
		6611 => to_unsigned(19406, LUT_AMPL_WIDTH - 1),
		6612 => to_unsigned(19408, LUT_AMPL_WIDTH - 1),
		6613 => to_unsigned(19411, LUT_AMPL_WIDTH - 1),
		6614 => to_unsigned(19413, LUT_AMPL_WIDTH - 1),
		6615 => to_unsigned(19416, LUT_AMPL_WIDTH - 1),
		6616 => to_unsigned(19418, LUT_AMPL_WIDTH - 1),
		6617 => to_unsigned(19421, LUT_AMPL_WIDTH - 1),
		6618 => to_unsigned(19423, LUT_AMPL_WIDTH - 1),
		6619 => to_unsigned(19426, LUT_AMPL_WIDTH - 1),
		6620 => to_unsigned(19428, LUT_AMPL_WIDTH - 1),
		6621 => to_unsigned(19431, LUT_AMPL_WIDTH - 1),
		6622 => to_unsigned(19433, LUT_AMPL_WIDTH - 1),
		6623 => to_unsigned(19436, LUT_AMPL_WIDTH - 1),
		6624 => to_unsigned(19438, LUT_AMPL_WIDTH - 1),
		6625 => to_unsigned(19441, LUT_AMPL_WIDTH - 1),
		6626 => to_unsigned(19444, LUT_AMPL_WIDTH - 1),
		6627 => to_unsigned(19446, LUT_AMPL_WIDTH - 1),
		6628 => to_unsigned(19449, LUT_AMPL_WIDTH - 1),
		6629 => to_unsigned(19451, LUT_AMPL_WIDTH - 1),
		6630 => to_unsigned(19454, LUT_AMPL_WIDTH - 1),
		6631 => to_unsigned(19456, LUT_AMPL_WIDTH - 1),
		6632 => to_unsigned(19459, LUT_AMPL_WIDTH - 1),
		6633 => to_unsigned(19461, LUT_AMPL_WIDTH - 1),
		6634 => to_unsigned(19464, LUT_AMPL_WIDTH - 1),
		6635 => to_unsigned(19466, LUT_AMPL_WIDTH - 1),
		6636 => to_unsigned(19469, LUT_AMPL_WIDTH - 1),
		6637 => to_unsigned(19471, LUT_AMPL_WIDTH - 1),
		6638 => to_unsigned(19474, LUT_AMPL_WIDTH - 1),
		6639 => to_unsigned(19476, LUT_AMPL_WIDTH - 1),
		6640 => to_unsigned(19479, LUT_AMPL_WIDTH - 1),
		6641 => to_unsigned(19481, LUT_AMPL_WIDTH - 1),
		6642 => to_unsigned(19484, LUT_AMPL_WIDTH - 1),
		6643 => to_unsigned(19486, LUT_AMPL_WIDTH - 1),
		6644 => to_unsigned(19489, LUT_AMPL_WIDTH - 1),
		6645 => to_unsigned(19492, LUT_AMPL_WIDTH - 1),
		6646 => to_unsigned(19494, LUT_AMPL_WIDTH - 1),
		6647 => to_unsigned(19497, LUT_AMPL_WIDTH - 1),
		6648 => to_unsigned(19499, LUT_AMPL_WIDTH - 1),
		6649 => to_unsigned(19502, LUT_AMPL_WIDTH - 1),
		6650 => to_unsigned(19504, LUT_AMPL_WIDTH - 1),
		6651 => to_unsigned(19507, LUT_AMPL_WIDTH - 1),
		6652 => to_unsigned(19509, LUT_AMPL_WIDTH - 1),
		6653 => to_unsigned(19512, LUT_AMPL_WIDTH - 1),
		6654 => to_unsigned(19514, LUT_AMPL_WIDTH - 1),
		6655 => to_unsigned(19517, LUT_AMPL_WIDTH - 1),
		6656 => to_unsigned(19519, LUT_AMPL_WIDTH - 1),
		6657 => to_unsigned(19522, LUT_AMPL_WIDTH - 1),
		6658 => to_unsigned(19524, LUT_AMPL_WIDTH - 1),
		6659 => to_unsigned(19527, LUT_AMPL_WIDTH - 1),
		6660 => to_unsigned(19529, LUT_AMPL_WIDTH - 1),
		6661 => to_unsigned(19532, LUT_AMPL_WIDTH - 1),
		6662 => to_unsigned(19534, LUT_AMPL_WIDTH - 1),
		6663 => to_unsigned(19537, LUT_AMPL_WIDTH - 1),
		6664 => to_unsigned(19539, LUT_AMPL_WIDTH - 1),
		6665 => to_unsigned(19542, LUT_AMPL_WIDTH - 1),
		6666 => to_unsigned(19545, LUT_AMPL_WIDTH - 1),
		6667 => to_unsigned(19547, LUT_AMPL_WIDTH - 1),
		6668 => to_unsigned(19550, LUT_AMPL_WIDTH - 1),
		6669 => to_unsigned(19552, LUT_AMPL_WIDTH - 1),
		6670 => to_unsigned(19555, LUT_AMPL_WIDTH - 1),
		6671 => to_unsigned(19557, LUT_AMPL_WIDTH - 1),
		6672 => to_unsigned(19560, LUT_AMPL_WIDTH - 1),
		6673 => to_unsigned(19562, LUT_AMPL_WIDTH - 1),
		6674 => to_unsigned(19565, LUT_AMPL_WIDTH - 1),
		6675 => to_unsigned(19567, LUT_AMPL_WIDTH - 1),
		6676 => to_unsigned(19570, LUT_AMPL_WIDTH - 1),
		6677 => to_unsigned(19572, LUT_AMPL_WIDTH - 1),
		6678 => to_unsigned(19575, LUT_AMPL_WIDTH - 1),
		6679 => to_unsigned(19577, LUT_AMPL_WIDTH - 1),
		6680 => to_unsigned(19580, LUT_AMPL_WIDTH - 1),
		6681 => to_unsigned(19582, LUT_AMPL_WIDTH - 1),
		6682 => to_unsigned(19585, LUT_AMPL_WIDTH - 1),
		6683 => to_unsigned(19587, LUT_AMPL_WIDTH - 1),
		6684 => to_unsigned(19590, LUT_AMPL_WIDTH - 1),
		6685 => to_unsigned(19592, LUT_AMPL_WIDTH - 1),
		6686 => to_unsigned(19595, LUT_AMPL_WIDTH - 1),
		6687 => to_unsigned(19597, LUT_AMPL_WIDTH - 1),
		6688 => to_unsigned(19600, LUT_AMPL_WIDTH - 1),
		6689 => to_unsigned(19602, LUT_AMPL_WIDTH - 1),
		6690 => to_unsigned(19605, LUT_AMPL_WIDTH - 1),
		6691 => to_unsigned(19607, LUT_AMPL_WIDTH - 1),
		6692 => to_unsigned(19610, LUT_AMPL_WIDTH - 1),
		6693 => to_unsigned(19613, LUT_AMPL_WIDTH - 1),
		6694 => to_unsigned(19615, LUT_AMPL_WIDTH - 1),
		6695 => to_unsigned(19618, LUT_AMPL_WIDTH - 1),
		6696 => to_unsigned(19620, LUT_AMPL_WIDTH - 1),
		6697 => to_unsigned(19623, LUT_AMPL_WIDTH - 1),
		6698 => to_unsigned(19625, LUT_AMPL_WIDTH - 1),
		6699 => to_unsigned(19628, LUT_AMPL_WIDTH - 1),
		6700 => to_unsigned(19630, LUT_AMPL_WIDTH - 1),
		6701 => to_unsigned(19633, LUT_AMPL_WIDTH - 1),
		6702 => to_unsigned(19635, LUT_AMPL_WIDTH - 1),
		6703 => to_unsigned(19638, LUT_AMPL_WIDTH - 1),
		6704 => to_unsigned(19640, LUT_AMPL_WIDTH - 1),
		6705 => to_unsigned(19643, LUT_AMPL_WIDTH - 1),
		6706 => to_unsigned(19645, LUT_AMPL_WIDTH - 1),
		6707 => to_unsigned(19648, LUT_AMPL_WIDTH - 1),
		6708 => to_unsigned(19650, LUT_AMPL_WIDTH - 1),
		6709 => to_unsigned(19653, LUT_AMPL_WIDTH - 1),
		6710 => to_unsigned(19655, LUT_AMPL_WIDTH - 1),
		6711 => to_unsigned(19658, LUT_AMPL_WIDTH - 1),
		6712 => to_unsigned(19660, LUT_AMPL_WIDTH - 1),
		6713 => to_unsigned(19663, LUT_AMPL_WIDTH - 1),
		6714 => to_unsigned(19665, LUT_AMPL_WIDTH - 1),
		6715 => to_unsigned(19668, LUT_AMPL_WIDTH - 1),
		6716 => to_unsigned(19670, LUT_AMPL_WIDTH - 1),
		6717 => to_unsigned(19673, LUT_AMPL_WIDTH - 1),
		6718 => to_unsigned(19675, LUT_AMPL_WIDTH - 1),
		6719 => to_unsigned(19678, LUT_AMPL_WIDTH - 1),
		6720 => to_unsigned(19680, LUT_AMPL_WIDTH - 1),
		6721 => to_unsigned(19683, LUT_AMPL_WIDTH - 1),
		6722 => to_unsigned(19685, LUT_AMPL_WIDTH - 1),
		6723 => to_unsigned(19688, LUT_AMPL_WIDTH - 1),
		6724 => to_unsigned(19690, LUT_AMPL_WIDTH - 1),
		6725 => to_unsigned(19693, LUT_AMPL_WIDTH - 1),
		6726 => to_unsigned(19695, LUT_AMPL_WIDTH - 1),
		6727 => to_unsigned(19698, LUT_AMPL_WIDTH - 1),
		6728 => to_unsigned(19700, LUT_AMPL_WIDTH - 1),
		6729 => to_unsigned(19703, LUT_AMPL_WIDTH - 1),
		6730 => to_unsigned(19706, LUT_AMPL_WIDTH - 1),
		6731 => to_unsigned(19708, LUT_AMPL_WIDTH - 1),
		6732 => to_unsigned(19711, LUT_AMPL_WIDTH - 1),
		6733 => to_unsigned(19713, LUT_AMPL_WIDTH - 1),
		6734 => to_unsigned(19716, LUT_AMPL_WIDTH - 1),
		6735 => to_unsigned(19718, LUT_AMPL_WIDTH - 1),
		6736 => to_unsigned(19721, LUT_AMPL_WIDTH - 1),
		6737 => to_unsigned(19723, LUT_AMPL_WIDTH - 1),
		6738 => to_unsigned(19726, LUT_AMPL_WIDTH - 1),
		6739 => to_unsigned(19728, LUT_AMPL_WIDTH - 1),
		6740 => to_unsigned(19731, LUT_AMPL_WIDTH - 1),
		6741 => to_unsigned(19733, LUT_AMPL_WIDTH - 1),
		6742 => to_unsigned(19736, LUT_AMPL_WIDTH - 1),
		6743 => to_unsigned(19738, LUT_AMPL_WIDTH - 1),
		6744 => to_unsigned(19741, LUT_AMPL_WIDTH - 1),
		6745 => to_unsigned(19743, LUT_AMPL_WIDTH - 1),
		6746 => to_unsigned(19746, LUT_AMPL_WIDTH - 1),
		6747 => to_unsigned(19748, LUT_AMPL_WIDTH - 1),
		6748 => to_unsigned(19751, LUT_AMPL_WIDTH - 1),
		6749 => to_unsigned(19753, LUT_AMPL_WIDTH - 1),
		6750 => to_unsigned(19756, LUT_AMPL_WIDTH - 1),
		6751 => to_unsigned(19758, LUT_AMPL_WIDTH - 1),
		6752 => to_unsigned(19761, LUT_AMPL_WIDTH - 1),
		6753 => to_unsigned(19763, LUT_AMPL_WIDTH - 1),
		6754 => to_unsigned(19766, LUT_AMPL_WIDTH - 1),
		6755 => to_unsigned(19768, LUT_AMPL_WIDTH - 1),
		6756 => to_unsigned(19771, LUT_AMPL_WIDTH - 1),
		6757 => to_unsigned(19773, LUT_AMPL_WIDTH - 1),
		6758 => to_unsigned(19776, LUT_AMPL_WIDTH - 1),
		6759 => to_unsigned(19778, LUT_AMPL_WIDTH - 1),
		6760 => to_unsigned(19781, LUT_AMPL_WIDTH - 1),
		6761 => to_unsigned(19783, LUT_AMPL_WIDTH - 1),
		6762 => to_unsigned(19786, LUT_AMPL_WIDTH - 1),
		6763 => to_unsigned(19788, LUT_AMPL_WIDTH - 1),
		6764 => to_unsigned(19791, LUT_AMPL_WIDTH - 1),
		6765 => to_unsigned(19793, LUT_AMPL_WIDTH - 1),
		6766 => to_unsigned(19796, LUT_AMPL_WIDTH - 1),
		6767 => to_unsigned(19798, LUT_AMPL_WIDTH - 1),
		6768 => to_unsigned(19801, LUT_AMPL_WIDTH - 1),
		6769 => to_unsigned(19803, LUT_AMPL_WIDTH - 1),
		6770 => to_unsigned(19806, LUT_AMPL_WIDTH - 1),
		6771 => to_unsigned(19808, LUT_AMPL_WIDTH - 1),
		6772 => to_unsigned(19811, LUT_AMPL_WIDTH - 1),
		6773 => to_unsigned(19813, LUT_AMPL_WIDTH - 1),
		6774 => to_unsigned(19816, LUT_AMPL_WIDTH - 1),
		6775 => to_unsigned(19818, LUT_AMPL_WIDTH - 1),
		6776 => to_unsigned(19821, LUT_AMPL_WIDTH - 1),
		6777 => to_unsigned(19823, LUT_AMPL_WIDTH - 1),
		6778 => to_unsigned(19826, LUT_AMPL_WIDTH - 1),
		6779 => to_unsigned(19828, LUT_AMPL_WIDTH - 1),
		6780 => to_unsigned(19831, LUT_AMPL_WIDTH - 1),
		6781 => to_unsigned(19833, LUT_AMPL_WIDTH - 1),
		6782 => to_unsigned(19836, LUT_AMPL_WIDTH - 1),
		6783 => to_unsigned(19838, LUT_AMPL_WIDTH - 1),
		6784 => to_unsigned(19841, LUT_AMPL_WIDTH - 1),
		6785 => to_unsigned(19843, LUT_AMPL_WIDTH - 1),
		6786 => to_unsigned(19846, LUT_AMPL_WIDTH - 1),
		6787 => to_unsigned(19848, LUT_AMPL_WIDTH - 1),
		6788 => to_unsigned(19851, LUT_AMPL_WIDTH - 1),
		6789 => to_unsigned(19853, LUT_AMPL_WIDTH - 1),
		6790 => to_unsigned(19856, LUT_AMPL_WIDTH - 1),
		6791 => to_unsigned(19858, LUT_AMPL_WIDTH - 1),
		6792 => to_unsigned(19861, LUT_AMPL_WIDTH - 1),
		6793 => to_unsigned(19863, LUT_AMPL_WIDTH - 1),
		6794 => to_unsigned(19866, LUT_AMPL_WIDTH - 1),
		6795 => to_unsigned(19868, LUT_AMPL_WIDTH - 1),
		6796 => to_unsigned(19871, LUT_AMPL_WIDTH - 1),
		6797 => to_unsigned(19873, LUT_AMPL_WIDTH - 1),
		6798 => to_unsigned(19876, LUT_AMPL_WIDTH - 1),
		6799 => to_unsigned(19878, LUT_AMPL_WIDTH - 1),
		6800 => to_unsigned(19881, LUT_AMPL_WIDTH - 1),
		6801 => to_unsigned(19883, LUT_AMPL_WIDTH - 1),
		6802 => to_unsigned(19886, LUT_AMPL_WIDTH - 1),
		6803 => to_unsigned(19888, LUT_AMPL_WIDTH - 1),
		6804 => to_unsigned(19891, LUT_AMPL_WIDTH - 1),
		6805 => to_unsigned(19893, LUT_AMPL_WIDTH - 1),
		6806 => to_unsigned(19896, LUT_AMPL_WIDTH - 1),
		6807 => to_unsigned(19898, LUT_AMPL_WIDTH - 1),
		6808 => to_unsigned(19901, LUT_AMPL_WIDTH - 1),
		6809 => to_unsigned(19903, LUT_AMPL_WIDTH - 1),
		6810 => to_unsigned(19906, LUT_AMPL_WIDTH - 1),
		6811 => to_unsigned(19908, LUT_AMPL_WIDTH - 1),
		6812 => to_unsigned(19911, LUT_AMPL_WIDTH - 1),
		6813 => to_unsigned(19913, LUT_AMPL_WIDTH - 1),
		6814 => to_unsigned(19916, LUT_AMPL_WIDTH - 1),
		6815 => to_unsigned(19918, LUT_AMPL_WIDTH - 1),
		6816 => to_unsigned(19921, LUT_AMPL_WIDTH - 1),
		6817 => to_unsigned(19923, LUT_AMPL_WIDTH - 1),
		6818 => to_unsigned(19926, LUT_AMPL_WIDTH - 1),
		6819 => to_unsigned(19928, LUT_AMPL_WIDTH - 1),
		6820 => to_unsigned(19931, LUT_AMPL_WIDTH - 1),
		6821 => to_unsigned(19933, LUT_AMPL_WIDTH - 1),
		6822 => to_unsigned(19936, LUT_AMPL_WIDTH - 1),
		6823 => to_unsigned(19938, LUT_AMPL_WIDTH - 1),
		6824 => to_unsigned(19941, LUT_AMPL_WIDTH - 1),
		6825 => to_unsigned(19943, LUT_AMPL_WIDTH - 1),
		6826 => to_unsigned(19946, LUT_AMPL_WIDTH - 1),
		6827 => to_unsigned(19948, LUT_AMPL_WIDTH - 1),
		6828 => to_unsigned(19951, LUT_AMPL_WIDTH - 1),
		6829 => to_unsigned(19953, LUT_AMPL_WIDTH - 1),
		6830 => to_unsigned(19956, LUT_AMPL_WIDTH - 1),
		6831 => to_unsigned(19958, LUT_AMPL_WIDTH - 1),
		6832 => to_unsigned(19961, LUT_AMPL_WIDTH - 1),
		6833 => to_unsigned(19963, LUT_AMPL_WIDTH - 1),
		6834 => to_unsigned(19966, LUT_AMPL_WIDTH - 1),
		6835 => to_unsigned(19968, LUT_AMPL_WIDTH - 1),
		6836 => to_unsigned(19971, LUT_AMPL_WIDTH - 1),
		6837 => to_unsigned(19973, LUT_AMPL_WIDTH - 1),
		6838 => to_unsigned(19976, LUT_AMPL_WIDTH - 1),
		6839 => to_unsigned(19978, LUT_AMPL_WIDTH - 1),
		6840 => to_unsigned(19981, LUT_AMPL_WIDTH - 1),
		6841 => to_unsigned(19983, LUT_AMPL_WIDTH - 1),
		6842 => to_unsigned(19985, LUT_AMPL_WIDTH - 1),
		6843 => to_unsigned(19988, LUT_AMPL_WIDTH - 1),
		6844 => to_unsigned(19990, LUT_AMPL_WIDTH - 1),
		6845 => to_unsigned(19993, LUT_AMPL_WIDTH - 1),
		6846 => to_unsigned(19995, LUT_AMPL_WIDTH - 1),
		6847 => to_unsigned(19998, LUT_AMPL_WIDTH - 1),
		6848 => to_unsigned(20000, LUT_AMPL_WIDTH - 1),
		6849 => to_unsigned(20003, LUT_AMPL_WIDTH - 1),
		6850 => to_unsigned(20005, LUT_AMPL_WIDTH - 1),
		6851 => to_unsigned(20008, LUT_AMPL_WIDTH - 1),
		6852 => to_unsigned(20010, LUT_AMPL_WIDTH - 1),
		6853 => to_unsigned(20013, LUT_AMPL_WIDTH - 1),
		6854 => to_unsigned(20015, LUT_AMPL_WIDTH - 1),
		6855 => to_unsigned(20018, LUT_AMPL_WIDTH - 1),
		6856 => to_unsigned(20020, LUT_AMPL_WIDTH - 1),
		6857 => to_unsigned(20023, LUT_AMPL_WIDTH - 1),
		6858 => to_unsigned(20025, LUT_AMPL_WIDTH - 1),
		6859 => to_unsigned(20028, LUT_AMPL_WIDTH - 1),
		6860 => to_unsigned(20030, LUT_AMPL_WIDTH - 1),
		6861 => to_unsigned(20033, LUT_AMPL_WIDTH - 1),
		6862 => to_unsigned(20035, LUT_AMPL_WIDTH - 1),
		6863 => to_unsigned(20038, LUT_AMPL_WIDTH - 1),
		6864 => to_unsigned(20040, LUT_AMPL_WIDTH - 1),
		6865 => to_unsigned(20043, LUT_AMPL_WIDTH - 1),
		6866 => to_unsigned(20045, LUT_AMPL_WIDTH - 1),
		6867 => to_unsigned(20048, LUT_AMPL_WIDTH - 1),
		6868 => to_unsigned(20050, LUT_AMPL_WIDTH - 1),
		6869 => to_unsigned(20053, LUT_AMPL_WIDTH - 1),
		6870 => to_unsigned(20055, LUT_AMPL_WIDTH - 1),
		6871 => to_unsigned(20058, LUT_AMPL_WIDTH - 1),
		6872 => to_unsigned(20060, LUT_AMPL_WIDTH - 1),
		6873 => to_unsigned(20063, LUT_AMPL_WIDTH - 1),
		6874 => to_unsigned(20065, LUT_AMPL_WIDTH - 1),
		6875 => to_unsigned(20068, LUT_AMPL_WIDTH - 1),
		6876 => to_unsigned(20070, LUT_AMPL_WIDTH - 1),
		6877 => to_unsigned(20072, LUT_AMPL_WIDTH - 1),
		6878 => to_unsigned(20075, LUT_AMPL_WIDTH - 1),
		6879 => to_unsigned(20077, LUT_AMPL_WIDTH - 1),
		6880 => to_unsigned(20080, LUT_AMPL_WIDTH - 1),
		6881 => to_unsigned(20082, LUT_AMPL_WIDTH - 1),
		6882 => to_unsigned(20085, LUT_AMPL_WIDTH - 1),
		6883 => to_unsigned(20087, LUT_AMPL_WIDTH - 1),
		6884 => to_unsigned(20090, LUT_AMPL_WIDTH - 1),
		6885 => to_unsigned(20092, LUT_AMPL_WIDTH - 1),
		6886 => to_unsigned(20095, LUT_AMPL_WIDTH - 1),
		6887 => to_unsigned(20097, LUT_AMPL_WIDTH - 1),
		6888 => to_unsigned(20100, LUT_AMPL_WIDTH - 1),
		6889 => to_unsigned(20102, LUT_AMPL_WIDTH - 1),
		6890 => to_unsigned(20105, LUT_AMPL_WIDTH - 1),
		6891 => to_unsigned(20107, LUT_AMPL_WIDTH - 1),
		6892 => to_unsigned(20110, LUT_AMPL_WIDTH - 1),
		6893 => to_unsigned(20112, LUT_AMPL_WIDTH - 1),
		6894 => to_unsigned(20115, LUT_AMPL_WIDTH - 1),
		6895 => to_unsigned(20117, LUT_AMPL_WIDTH - 1),
		6896 => to_unsigned(20120, LUT_AMPL_WIDTH - 1),
		6897 => to_unsigned(20122, LUT_AMPL_WIDTH - 1),
		6898 => to_unsigned(20125, LUT_AMPL_WIDTH - 1),
		6899 => to_unsigned(20127, LUT_AMPL_WIDTH - 1),
		6900 => to_unsigned(20130, LUT_AMPL_WIDTH - 1),
		6901 => to_unsigned(20132, LUT_AMPL_WIDTH - 1),
		6902 => to_unsigned(20135, LUT_AMPL_WIDTH - 1),
		6903 => to_unsigned(20137, LUT_AMPL_WIDTH - 1),
		6904 => to_unsigned(20139, LUT_AMPL_WIDTH - 1),
		6905 => to_unsigned(20142, LUT_AMPL_WIDTH - 1),
		6906 => to_unsigned(20144, LUT_AMPL_WIDTH - 1),
		6907 => to_unsigned(20147, LUT_AMPL_WIDTH - 1),
		6908 => to_unsigned(20149, LUT_AMPL_WIDTH - 1),
		6909 => to_unsigned(20152, LUT_AMPL_WIDTH - 1),
		6910 => to_unsigned(20154, LUT_AMPL_WIDTH - 1),
		6911 => to_unsigned(20157, LUT_AMPL_WIDTH - 1),
		6912 => to_unsigned(20159, LUT_AMPL_WIDTH - 1),
		6913 => to_unsigned(20162, LUT_AMPL_WIDTH - 1),
		6914 => to_unsigned(20164, LUT_AMPL_WIDTH - 1),
		6915 => to_unsigned(20167, LUT_AMPL_WIDTH - 1),
		6916 => to_unsigned(20169, LUT_AMPL_WIDTH - 1),
		6917 => to_unsigned(20172, LUT_AMPL_WIDTH - 1),
		6918 => to_unsigned(20174, LUT_AMPL_WIDTH - 1),
		6919 => to_unsigned(20177, LUT_AMPL_WIDTH - 1),
		6920 => to_unsigned(20179, LUT_AMPL_WIDTH - 1),
		6921 => to_unsigned(20182, LUT_AMPL_WIDTH - 1),
		6922 => to_unsigned(20184, LUT_AMPL_WIDTH - 1),
		6923 => to_unsigned(20187, LUT_AMPL_WIDTH - 1),
		6924 => to_unsigned(20189, LUT_AMPL_WIDTH - 1),
		6925 => to_unsigned(20191, LUT_AMPL_WIDTH - 1),
		6926 => to_unsigned(20194, LUT_AMPL_WIDTH - 1),
		6927 => to_unsigned(20196, LUT_AMPL_WIDTH - 1),
		6928 => to_unsigned(20199, LUT_AMPL_WIDTH - 1),
		6929 => to_unsigned(20201, LUT_AMPL_WIDTH - 1),
		6930 => to_unsigned(20204, LUT_AMPL_WIDTH - 1),
		6931 => to_unsigned(20206, LUT_AMPL_WIDTH - 1),
		6932 => to_unsigned(20209, LUT_AMPL_WIDTH - 1),
		6933 => to_unsigned(20211, LUT_AMPL_WIDTH - 1),
		6934 => to_unsigned(20214, LUT_AMPL_WIDTH - 1),
		6935 => to_unsigned(20216, LUT_AMPL_WIDTH - 1),
		6936 => to_unsigned(20219, LUT_AMPL_WIDTH - 1),
		6937 => to_unsigned(20221, LUT_AMPL_WIDTH - 1),
		6938 => to_unsigned(20224, LUT_AMPL_WIDTH - 1),
		6939 => to_unsigned(20226, LUT_AMPL_WIDTH - 1),
		6940 => to_unsigned(20229, LUT_AMPL_WIDTH - 1),
		6941 => to_unsigned(20231, LUT_AMPL_WIDTH - 1),
		6942 => to_unsigned(20234, LUT_AMPL_WIDTH - 1),
		6943 => to_unsigned(20236, LUT_AMPL_WIDTH - 1),
		6944 => to_unsigned(20238, LUT_AMPL_WIDTH - 1),
		6945 => to_unsigned(20241, LUT_AMPL_WIDTH - 1),
		6946 => to_unsigned(20243, LUT_AMPL_WIDTH - 1),
		6947 => to_unsigned(20246, LUT_AMPL_WIDTH - 1),
		6948 => to_unsigned(20248, LUT_AMPL_WIDTH - 1),
		6949 => to_unsigned(20251, LUT_AMPL_WIDTH - 1),
		6950 => to_unsigned(20253, LUT_AMPL_WIDTH - 1),
		6951 => to_unsigned(20256, LUT_AMPL_WIDTH - 1),
		6952 => to_unsigned(20258, LUT_AMPL_WIDTH - 1),
		6953 => to_unsigned(20261, LUT_AMPL_WIDTH - 1),
		6954 => to_unsigned(20263, LUT_AMPL_WIDTH - 1),
		6955 => to_unsigned(20266, LUT_AMPL_WIDTH - 1),
		6956 => to_unsigned(20268, LUT_AMPL_WIDTH - 1),
		6957 => to_unsigned(20271, LUT_AMPL_WIDTH - 1),
		6958 => to_unsigned(20273, LUT_AMPL_WIDTH - 1),
		6959 => to_unsigned(20275, LUT_AMPL_WIDTH - 1),
		6960 => to_unsigned(20278, LUT_AMPL_WIDTH - 1),
		6961 => to_unsigned(20280, LUT_AMPL_WIDTH - 1),
		6962 => to_unsigned(20283, LUT_AMPL_WIDTH - 1),
		6963 => to_unsigned(20285, LUT_AMPL_WIDTH - 1),
		6964 => to_unsigned(20288, LUT_AMPL_WIDTH - 1),
		6965 => to_unsigned(20290, LUT_AMPL_WIDTH - 1),
		6966 => to_unsigned(20293, LUT_AMPL_WIDTH - 1),
		6967 => to_unsigned(20295, LUT_AMPL_WIDTH - 1),
		6968 => to_unsigned(20298, LUT_AMPL_WIDTH - 1),
		6969 => to_unsigned(20300, LUT_AMPL_WIDTH - 1),
		6970 => to_unsigned(20303, LUT_AMPL_WIDTH - 1),
		6971 => to_unsigned(20305, LUT_AMPL_WIDTH - 1),
		6972 => to_unsigned(20308, LUT_AMPL_WIDTH - 1),
		6973 => to_unsigned(20310, LUT_AMPL_WIDTH - 1),
		6974 => to_unsigned(20312, LUT_AMPL_WIDTH - 1),
		6975 => to_unsigned(20315, LUT_AMPL_WIDTH - 1),
		6976 => to_unsigned(20317, LUT_AMPL_WIDTH - 1),
		6977 => to_unsigned(20320, LUT_AMPL_WIDTH - 1),
		6978 => to_unsigned(20322, LUT_AMPL_WIDTH - 1),
		6979 => to_unsigned(20325, LUT_AMPL_WIDTH - 1),
		6980 => to_unsigned(20327, LUT_AMPL_WIDTH - 1),
		6981 => to_unsigned(20330, LUT_AMPL_WIDTH - 1),
		6982 => to_unsigned(20332, LUT_AMPL_WIDTH - 1),
		6983 => to_unsigned(20335, LUT_AMPL_WIDTH - 1),
		6984 => to_unsigned(20337, LUT_AMPL_WIDTH - 1),
		6985 => to_unsigned(20340, LUT_AMPL_WIDTH - 1),
		6986 => to_unsigned(20342, LUT_AMPL_WIDTH - 1),
		6987 => to_unsigned(20345, LUT_AMPL_WIDTH - 1),
		6988 => to_unsigned(20347, LUT_AMPL_WIDTH - 1),
		6989 => to_unsigned(20349, LUT_AMPL_WIDTH - 1),
		6990 => to_unsigned(20352, LUT_AMPL_WIDTH - 1),
		6991 => to_unsigned(20354, LUT_AMPL_WIDTH - 1),
		6992 => to_unsigned(20357, LUT_AMPL_WIDTH - 1),
		6993 => to_unsigned(20359, LUT_AMPL_WIDTH - 1),
		6994 => to_unsigned(20362, LUT_AMPL_WIDTH - 1),
		6995 => to_unsigned(20364, LUT_AMPL_WIDTH - 1),
		6996 => to_unsigned(20367, LUT_AMPL_WIDTH - 1),
		6997 => to_unsigned(20369, LUT_AMPL_WIDTH - 1),
		6998 => to_unsigned(20372, LUT_AMPL_WIDTH - 1),
		6999 => to_unsigned(20374, LUT_AMPL_WIDTH - 1),
		7000 => to_unsigned(20377, LUT_AMPL_WIDTH - 1),
		7001 => to_unsigned(20379, LUT_AMPL_WIDTH - 1),
		7002 => to_unsigned(20381, LUT_AMPL_WIDTH - 1),
		7003 => to_unsigned(20384, LUT_AMPL_WIDTH - 1),
		7004 => to_unsigned(20386, LUT_AMPL_WIDTH - 1),
		7005 => to_unsigned(20389, LUT_AMPL_WIDTH - 1),
		7006 => to_unsigned(20391, LUT_AMPL_WIDTH - 1),
		7007 => to_unsigned(20394, LUT_AMPL_WIDTH - 1),
		7008 => to_unsigned(20396, LUT_AMPL_WIDTH - 1),
		7009 => to_unsigned(20399, LUT_AMPL_WIDTH - 1),
		7010 => to_unsigned(20401, LUT_AMPL_WIDTH - 1),
		7011 => to_unsigned(20404, LUT_AMPL_WIDTH - 1),
		7012 => to_unsigned(20406, LUT_AMPL_WIDTH - 1),
		7013 => to_unsigned(20408, LUT_AMPL_WIDTH - 1),
		7014 => to_unsigned(20411, LUT_AMPL_WIDTH - 1),
		7015 => to_unsigned(20413, LUT_AMPL_WIDTH - 1),
		7016 => to_unsigned(20416, LUT_AMPL_WIDTH - 1),
		7017 => to_unsigned(20418, LUT_AMPL_WIDTH - 1),
		7018 => to_unsigned(20421, LUT_AMPL_WIDTH - 1),
		7019 => to_unsigned(20423, LUT_AMPL_WIDTH - 1),
		7020 => to_unsigned(20426, LUT_AMPL_WIDTH - 1),
		7021 => to_unsigned(20428, LUT_AMPL_WIDTH - 1),
		7022 => to_unsigned(20431, LUT_AMPL_WIDTH - 1),
		7023 => to_unsigned(20433, LUT_AMPL_WIDTH - 1),
		7024 => to_unsigned(20436, LUT_AMPL_WIDTH - 1),
		7025 => to_unsigned(20438, LUT_AMPL_WIDTH - 1),
		7026 => to_unsigned(20440, LUT_AMPL_WIDTH - 1),
		7027 => to_unsigned(20443, LUT_AMPL_WIDTH - 1),
		7028 => to_unsigned(20445, LUT_AMPL_WIDTH - 1),
		7029 => to_unsigned(20448, LUT_AMPL_WIDTH - 1),
		7030 => to_unsigned(20450, LUT_AMPL_WIDTH - 1),
		7031 => to_unsigned(20453, LUT_AMPL_WIDTH - 1),
		7032 => to_unsigned(20455, LUT_AMPL_WIDTH - 1),
		7033 => to_unsigned(20458, LUT_AMPL_WIDTH - 1),
		7034 => to_unsigned(20460, LUT_AMPL_WIDTH - 1),
		7035 => to_unsigned(20463, LUT_AMPL_WIDTH - 1),
		7036 => to_unsigned(20465, LUT_AMPL_WIDTH - 1),
		7037 => to_unsigned(20467, LUT_AMPL_WIDTH - 1),
		7038 => to_unsigned(20470, LUT_AMPL_WIDTH - 1),
		7039 => to_unsigned(20472, LUT_AMPL_WIDTH - 1),
		7040 => to_unsigned(20475, LUT_AMPL_WIDTH - 1),
		7041 => to_unsigned(20477, LUT_AMPL_WIDTH - 1),
		7042 => to_unsigned(20480, LUT_AMPL_WIDTH - 1),
		7043 => to_unsigned(20482, LUT_AMPL_WIDTH - 1),
		7044 => to_unsigned(20485, LUT_AMPL_WIDTH - 1),
		7045 => to_unsigned(20487, LUT_AMPL_WIDTH - 1),
		7046 => to_unsigned(20489, LUT_AMPL_WIDTH - 1),
		7047 => to_unsigned(20492, LUT_AMPL_WIDTH - 1),
		7048 => to_unsigned(20494, LUT_AMPL_WIDTH - 1),
		7049 => to_unsigned(20497, LUT_AMPL_WIDTH - 1),
		7050 => to_unsigned(20499, LUT_AMPL_WIDTH - 1),
		7051 => to_unsigned(20502, LUT_AMPL_WIDTH - 1),
		7052 => to_unsigned(20504, LUT_AMPL_WIDTH - 1),
		7053 => to_unsigned(20507, LUT_AMPL_WIDTH - 1),
		7054 => to_unsigned(20509, LUT_AMPL_WIDTH - 1),
		7055 => to_unsigned(20512, LUT_AMPL_WIDTH - 1),
		7056 => to_unsigned(20514, LUT_AMPL_WIDTH - 1),
		7057 => to_unsigned(20516, LUT_AMPL_WIDTH - 1),
		7058 => to_unsigned(20519, LUT_AMPL_WIDTH - 1),
		7059 => to_unsigned(20521, LUT_AMPL_WIDTH - 1),
		7060 => to_unsigned(20524, LUT_AMPL_WIDTH - 1),
		7061 => to_unsigned(20526, LUT_AMPL_WIDTH - 1),
		7062 => to_unsigned(20529, LUT_AMPL_WIDTH - 1),
		7063 => to_unsigned(20531, LUT_AMPL_WIDTH - 1),
		7064 => to_unsigned(20534, LUT_AMPL_WIDTH - 1),
		7065 => to_unsigned(20536, LUT_AMPL_WIDTH - 1),
		7066 => to_unsigned(20538, LUT_AMPL_WIDTH - 1),
		7067 => to_unsigned(20541, LUT_AMPL_WIDTH - 1),
		7068 => to_unsigned(20543, LUT_AMPL_WIDTH - 1),
		7069 => to_unsigned(20546, LUT_AMPL_WIDTH - 1),
		7070 => to_unsigned(20548, LUT_AMPL_WIDTH - 1),
		7071 => to_unsigned(20551, LUT_AMPL_WIDTH - 1),
		7072 => to_unsigned(20553, LUT_AMPL_WIDTH - 1),
		7073 => to_unsigned(20556, LUT_AMPL_WIDTH - 1),
		7074 => to_unsigned(20558, LUT_AMPL_WIDTH - 1),
		7075 => to_unsigned(20560, LUT_AMPL_WIDTH - 1),
		7076 => to_unsigned(20563, LUT_AMPL_WIDTH - 1),
		7077 => to_unsigned(20565, LUT_AMPL_WIDTH - 1),
		7078 => to_unsigned(20568, LUT_AMPL_WIDTH - 1),
		7079 => to_unsigned(20570, LUT_AMPL_WIDTH - 1),
		7080 => to_unsigned(20573, LUT_AMPL_WIDTH - 1),
		7081 => to_unsigned(20575, LUT_AMPL_WIDTH - 1),
		7082 => to_unsigned(20578, LUT_AMPL_WIDTH - 1),
		7083 => to_unsigned(20580, LUT_AMPL_WIDTH - 1),
		7084 => to_unsigned(20583, LUT_AMPL_WIDTH - 1),
		7085 => to_unsigned(20585, LUT_AMPL_WIDTH - 1),
		7086 => to_unsigned(20587, LUT_AMPL_WIDTH - 1),
		7087 => to_unsigned(20590, LUT_AMPL_WIDTH - 1),
		7088 => to_unsigned(20592, LUT_AMPL_WIDTH - 1),
		7089 => to_unsigned(20595, LUT_AMPL_WIDTH - 1),
		7090 => to_unsigned(20597, LUT_AMPL_WIDTH - 1),
		7091 => to_unsigned(20600, LUT_AMPL_WIDTH - 1),
		7092 => to_unsigned(20602, LUT_AMPL_WIDTH - 1),
		7093 => to_unsigned(20604, LUT_AMPL_WIDTH - 1),
		7094 => to_unsigned(20607, LUT_AMPL_WIDTH - 1),
		7095 => to_unsigned(20609, LUT_AMPL_WIDTH - 1),
		7096 => to_unsigned(20612, LUT_AMPL_WIDTH - 1),
		7097 => to_unsigned(20614, LUT_AMPL_WIDTH - 1),
		7098 => to_unsigned(20617, LUT_AMPL_WIDTH - 1),
		7099 => to_unsigned(20619, LUT_AMPL_WIDTH - 1),
		7100 => to_unsigned(20622, LUT_AMPL_WIDTH - 1),
		7101 => to_unsigned(20624, LUT_AMPL_WIDTH - 1),
		7102 => to_unsigned(20626, LUT_AMPL_WIDTH - 1),
		7103 => to_unsigned(20629, LUT_AMPL_WIDTH - 1),
		7104 => to_unsigned(20631, LUT_AMPL_WIDTH - 1),
		7105 => to_unsigned(20634, LUT_AMPL_WIDTH - 1),
		7106 => to_unsigned(20636, LUT_AMPL_WIDTH - 1),
		7107 => to_unsigned(20639, LUT_AMPL_WIDTH - 1),
		7108 => to_unsigned(20641, LUT_AMPL_WIDTH - 1),
		7109 => to_unsigned(20644, LUT_AMPL_WIDTH - 1),
		7110 => to_unsigned(20646, LUT_AMPL_WIDTH - 1),
		7111 => to_unsigned(20648, LUT_AMPL_WIDTH - 1),
		7112 => to_unsigned(20651, LUT_AMPL_WIDTH - 1),
		7113 => to_unsigned(20653, LUT_AMPL_WIDTH - 1),
		7114 => to_unsigned(20656, LUT_AMPL_WIDTH - 1),
		7115 => to_unsigned(20658, LUT_AMPL_WIDTH - 1),
		7116 => to_unsigned(20661, LUT_AMPL_WIDTH - 1),
		7117 => to_unsigned(20663, LUT_AMPL_WIDTH - 1),
		7118 => to_unsigned(20666, LUT_AMPL_WIDTH - 1),
		7119 => to_unsigned(20668, LUT_AMPL_WIDTH - 1),
		7120 => to_unsigned(20670, LUT_AMPL_WIDTH - 1),
		7121 => to_unsigned(20673, LUT_AMPL_WIDTH - 1),
		7122 => to_unsigned(20675, LUT_AMPL_WIDTH - 1),
		7123 => to_unsigned(20678, LUT_AMPL_WIDTH - 1),
		7124 => to_unsigned(20680, LUT_AMPL_WIDTH - 1),
		7125 => to_unsigned(20683, LUT_AMPL_WIDTH - 1),
		7126 => to_unsigned(20685, LUT_AMPL_WIDTH - 1),
		7127 => to_unsigned(20687, LUT_AMPL_WIDTH - 1),
		7128 => to_unsigned(20690, LUT_AMPL_WIDTH - 1),
		7129 => to_unsigned(20692, LUT_AMPL_WIDTH - 1),
		7130 => to_unsigned(20695, LUT_AMPL_WIDTH - 1),
		7131 => to_unsigned(20697, LUT_AMPL_WIDTH - 1),
		7132 => to_unsigned(20700, LUT_AMPL_WIDTH - 1),
		7133 => to_unsigned(20702, LUT_AMPL_WIDTH - 1),
		7134 => to_unsigned(20704, LUT_AMPL_WIDTH - 1),
		7135 => to_unsigned(20707, LUT_AMPL_WIDTH - 1),
		7136 => to_unsigned(20709, LUT_AMPL_WIDTH - 1),
		7137 => to_unsigned(20712, LUT_AMPL_WIDTH - 1),
		7138 => to_unsigned(20714, LUT_AMPL_WIDTH - 1),
		7139 => to_unsigned(20717, LUT_AMPL_WIDTH - 1),
		7140 => to_unsigned(20719, LUT_AMPL_WIDTH - 1),
		7141 => to_unsigned(20722, LUT_AMPL_WIDTH - 1),
		7142 => to_unsigned(20724, LUT_AMPL_WIDTH - 1),
		7143 => to_unsigned(20726, LUT_AMPL_WIDTH - 1),
		7144 => to_unsigned(20729, LUT_AMPL_WIDTH - 1),
		7145 => to_unsigned(20731, LUT_AMPL_WIDTH - 1),
		7146 => to_unsigned(20734, LUT_AMPL_WIDTH - 1),
		7147 => to_unsigned(20736, LUT_AMPL_WIDTH - 1),
		7148 => to_unsigned(20739, LUT_AMPL_WIDTH - 1),
		7149 => to_unsigned(20741, LUT_AMPL_WIDTH - 1),
		7150 => to_unsigned(20743, LUT_AMPL_WIDTH - 1),
		7151 => to_unsigned(20746, LUT_AMPL_WIDTH - 1),
		7152 => to_unsigned(20748, LUT_AMPL_WIDTH - 1),
		7153 => to_unsigned(20751, LUT_AMPL_WIDTH - 1),
		7154 => to_unsigned(20753, LUT_AMPL_WIDTH - 1),
		7155 => to_unsigned(20756, LUT_AMPL_WIDTH - 1),
		7156 => to_unsigned(20758, LUT_AMPL_WIDTH - 1),
		7157 => to_unsigned(20760, LUT_AMPL_WIDTH - 1),
		7158 => to_unsigned(20763, LUT_AMPL_WIDTH - 1),
		7159 => to_unsigned(20765, LUT_AMPL_WIDTH - 1),
		7160 => to_unsigned(20768, LUT_AMPL_WIDTH - 1),
		7161 => to_unsigned(20770, LUT_AMPL_WIDTH - 1),
		7162 => to_unsigned(20773, LUT_AMPL_WIDTH - 1),
		7163 => to_unsigned(20775, LUT_AMPL_WIDTH - 1),
		7164 => to_unsigned(20777, LUT_AMPL_WIDTH - 1),
		7165 => to_unsigned(20780, LUT_AMPL_WIDTH - 1),
		7166 => to_unsigned(20782, LUT_AMPL_WIDTH - 1),
		7167 => to_unsigned(20785, LUT_AMPL_WIDTH - 1),
		7168 => to_unsigned(20787, LUT_AMPL_WIDTH - 1),
		7169 => to_unsigned(20790, LUT_AMPL_WIDTH - 1),
		7170 => to_unsigned(20792, LUT_AMPL_WIDTH - 1),
		7171 => to_unsigned(20794, LUT_AMPL_WIDTH - 1),
		7172 => to_unsigned(20797, LUT_AMPL_WIDTH - 1),
		7173 => to_unsigned(20799, LUT_AMPL_WIDTH - 1),
		7174 => to_unsigned(20802, LUT_AMPL_WIDTH - 1),
		7175 => to_unsigned(20804, LUT_AMPL_WIDTH - 1),
		7176 => to_unsigned(20807, LUT_AMPL_WIDTH - 1),
		7177 => to_unsigned(20809, LUT_AMPL_WIDTH - 1),
		7178 => to_unsigned(20811, LUT_AMPL_WIDTH - 1),
		7179 => to_unsigned(20814, LUT_AMPL_WIDTH - 1),
		7180 => to_unsigned(20816, LUT_AMPL_WIDTH - 1),
		7181 => to_unsigned(20819, LUT_AMPL_WIDTH - 1),
		7182 => to_unsigned(20821, LUT_AMPL_WIDTH - 1),
		7183 => to_unsigned(20824, LUT_AMPL_WIDTH - 1),
		7184 => to_unsigned(20826, LUT_AMPL_WIDTH - 1),
		7185 => to_unsigned(20828, LUT_AMPL_WIDTH - 1),
		7186 => to_unsigned(20831, LUT_AMPL_WIDTH - 1),
		7187 => to_unsigned(20833, LUT_AMPL_WIDTH - 1),
		7188 => to_unsigned(20836, LUT_AMPL_WIDTH - 1),
		7189 => to_unsigned(20838, LUT_AMPL_WIDTH - 1),
		7190 => to_unsigned(20841, LUT_AMPL_WIDTH - 1),
		7191 => to_unsigned(20843, LUT_AMPL_WIDTH - 1),
		7192 => to_unsigned(20845, LUT_AMPL_WIDTH - 1),
		7193 => to_unsigned(20848, LUT_AMPL_WIDTH - 1),
		7194 => to_unsigned(20850, LUT_AMPL_WIDTH - 1),
		7195 => to_unsigned(20853, LUT_AMPL_WIDTH - 1),
		7196 => to_unsigned(20855, LUT_AMPL_WIDTH - 1),
		7197 => to_unsigned(20858, LUT_AMPL_WIDTH - 1),
		7198 => to_unsigned(20860, LUT_AMPL_WIDTH - 1),
		7199 => to_unsigned(20862, LUT_AMPL_WIDTH - 1),
		7200 => to_unsigned(20865, LUT_AMPL_WIDTH - 1),
		7201 => to_unsigned(20867, LUT_AMPL_WIDTH - 1),
		7202 => to_unsigned(20870, LUT_AMPL_WIDTH - 1),
		7203 => to_unsigned(20872, LUT_AMPL_WIDTH - 1),
		7204 => to_unsigned(20874, LUT_AMPL_WIDTH - 1),
		7205 => to_unsigned(20877, LUT_AMPL_WIDTH - 1),
		7206 => to_unsigned(20879, LUT_AMPL_WIDTH - 1),
		7207 => to_unsigned(20882, LUT_AMPL_WIDTH - 1),
		7208 => to_unsigned(20884, LUT_AMPL_WIDTH - 1),
		7209 => to_unsigned(20887, LUT_AMPL_WIDTH - 1),
		7210 => to_unsigned(20889, LUT_AMPL_WIDTH - 1),
		7211 => to_unsigned(20891, LUT_AMPL_WIDTH - 1),
		7212 => to_unsigned(20894, LUT_AMPL_WIDTH - 1),
		7213 => to_unsigned(20896, LUT_AMPL_WIDTH - 1),
		7214 => to_unsigned(20899, LUT_AMPL_WIDTH - 1),
		7215 => to_unsigned(20901, LUT_AMPL_WIDTH - 1),
		7216 => to_unsigned(20904, LUT_AMPL_WIDTH - 1),
		7217 => to_unsigned(20906, LUT_AMPL_WIDTH - 1),
		7218 => to_unsigned(20908, LUT_AMPL_WIDTH - 1),
		7219 => to_unsigned(20911, LUT_AMPL_WIDTH - 1),
		7220 => to_unsigned(20913, LUT_AMPL_WIDTH - 1),
		7221 => to_unsigned(20916, LUT_AMPL_WIDTH - 1),
		7222 => to_unsigned(20918, LUT_AMPL_WIDTH - 1),
		7223 => to_unsigned(20920, LUT_AMPL_WIDTH - 1),
		7224 => to_unsigned(20923, LUT_AMPL_WIDTH - 1),
		7225 => to_unsigned(20925, LUT_AMPL_WIDTH - 1),
		7226 => to_unsigned(20928, LUT_AMPL_WIDTH - 1),
		7227 => to_unsigned(20930, LUT_AMPL_WIDTH - 1),
		7228 => to_unsigned(20933, LUT_AMPL_WIDTH - 1),
		7229 => to_unsigned(20935, LUT_AMPL_WIDTH - 1),
		7230 => to_unsigned(20937, LUT_AMPL_WIDTH - 1),
		7231 => to_unsigned(20940, LUT_AMPL_WIDTH - 1),
		7232 => to_unsigned(20942, LUT_AMPL_WIDTH - 1),
		7233 => to_unsigned(20945, LUT_AMPL_WIDTH - 1),
		7234 => to_unsigned(20947, LUT_AMPL_WIDTH - 1),
		7235 => to_unsigned(20949, LUT_AMPL_WIDTH - 1),
		7236 => to_unsigned(20952, LUT_AMPL_WIDTH - 1),
		7237 => to_unsigned(20954, LUT_AMPL_WIDTH - 1),
		7238 => to_unsigned(20957, LUT_AMPL_WIDTH - 1),
		7239 => to_unsigned(20959, LUT_AMPL_WIDTH - 1),
		7240 => to_unsigned(20962, LUT_AMPL_WIDTH - 1),
		7241 => to_unsigned(20964, LUT_AMPL_WIDTH - 1),
		7242 => to_unsigned(20966, LUT_AMPL_WIDTH - 1),
		7243 => to_unsigned(20969, LUT_AMPL_WIDTH - 1),
		7244 => to_unsigned(20971, LUT_AMPL_WIDTH - 1),
		7245 => to_unsigned(20974, LUT_AMPL_WIDTH - 1),
		7246 => to_unsigned(20976, LUT_AMPL_WIDTH - 1),
		7247 => to_unsigned(20978, LUT_AMPL_WIDTH - 1),
		7248 => to_unsigned(20981, LUT_AMPL_WIDTH - 1),
		7249 => to_unsigned(20983, LUT_AMPL_WIDTH - 1),
		7250 => to_unsigned(20986, LUT_AMPL_WIDTH - 1),
		7251 => to_unsigned(20988, LUT_AMPL_WIDTH - 1),
		7252 => to_unsigned(20990, LUT_AMPL_WIDTH - 1),
		7253 => to_unsigned(20993, LUT_AMPL_WIDTH - 1),
		7254 => to_unsigned(20995, LUT_AMPL_WIDTH - 1),
		7255 => to_unsigned(20998, LUT_AMPL_WIDTH - 1),
		7256 => to_unsigned(21000, LUT_AMPL_WIDTH - 1),
		7257 => to_unsigned(21003, LUT_AMPL_WIDTH - 1),
		7258 => to_unsigned(21005, LUT_AMPL_WIDTH - 1),
		7259 => to_unsigned(21007, LUT_AMPL_WIDTH - 1),
		7260 => to_unsigned(21010, LUT_AMPL_WIDTH - 1),
		7261 => to_unsigned(21012, LUT_AMPL_WIDTH - 1),
		7262 => to_unsigned(21015, LUT_AMPL_WIDTH - 1),
		7263 => to_unsigned(21017, LUT_AMPL_WIDTH - 1),
		7264 => to_unsigned(21019, LUT_AMPL_WIDTH - 1),
		7265 => to_unsigned(21022, LUT_AMPL_WIDTH - 1),
		7266 => to_unsigned(21024, LUT_AMPL_WIDTH - 1),
		7267 => to_unsigned(21027, LUT_AMPL_WIDTH - 1),
		7268 => to_unsigned(21029, LUT_AMPL_WIDTH - 1),
		7269 => to_unsigned(21031, LUT_AMPL_WIDTH - 1),
		7270 => to_unsigned(21034, LUT_AMPL_WIDTH - 1),
		7271 => to_unsigned(21036, LUT_AMPL_WIDTH - 1),
		7272 => to_unsigned(21039, LUT_AMPL_WIDTH - 1),
		7273 => to_unsigned(21041, LUT_AMPL_WIDTH - 1),
		7274 => to_unsigned(21043, LUT_AMPL_WIDTH - 1),
		7275 => to_unsigned(21046, LUT_AMPL_WIDTH - 1),
		7276 => to_unsigned(21048, LUT_AMPL_WIDTH - 1),
		7277 => to_unsigned(21051, LUT_AMPL_WIDTH - 1),
		7278 => to_unsigned(21053, LUT_AMPL_WIDTH - 1),
		7279 => to_unsigned(21056, LUT_AMPL_WIDTH - 1),
		7280 => to_unsigned(21058, LUT_AMPL_WIDTH - 1),
		7281 => to_unsigned(21060, LUT_AMPL_WIDTH - 1),
		7282 => to_unsigned(21063, LUT_AMPL_WIDTH - 1),
		7283 => to_unsigned(21065, LUT_AMPL_WIDTH - 1),
		7284 => to_unsigned(21068, LUT_AMPL_WIDTH - 1),
		7285 => to_unsigned(21070, LUT_AMPL_WIDTH - 1),
		7286 => to_unsigned(21072, LUT_AMPL_WIDTH - 1),
		7287 => to_unsigned(21075, LUT_AMPL_WIDTH - 1),
		7288 => to_unsigned(21077, LUT_AMPL_WIDTH - 1),
		7289 => to_unsigned(21080, LUT_AMPL_WIDTH - 1),
		7290 => to_unsigned(21082, LUT_AMPL_WIDTH - 1),
		7291 => to_unsigned(21084, LUT_AMPL_WIDTH - 1),
		7292 => to_unsigned(21087, LUT_AMPL_WIDTH - 1),
		7293 => to_unsigned(21089, LUT_AMPL_WIDTH - 1),
		7294 => to_unsigned(21092, LUT_AMPL_WIDTH - 1),
		7295 => to_unsigned(21094, LUT_AMPL_WIDTH - 1),
		7296 => to_unsigned(21096, LUT_AMPL_WIDTH - 1),
		7297 => to_unsigned(21099, LUT_AMPL_WIDTH - 1),
		7298 => to_unsigned(21101, LUT_AMPL_WIDTH - 1),
		7299 => to_unsigned(21104, LUT_AMPL_WIDTH - 1),
		7300 => to_unsigned(21106, LUT_AMPL_WIDTH - 1),
		7301 => to_unsigned(21108, LUT_AMPL_WIDTH - 1),
		7302 => to_unsigned(21111, LUT_AMPL_WIDTH - 1),
		7303 => to_unsigned(21113, LUT_AMPL_WIDTH - 1),
		7304 => to_unsigned(21116, LUT_AMPL_WIDTH - 1),
		7305 => to_unsigned(21118, LUT_AMPL_WIDTH - 1),
		7306 => to_unsigned(21120, LUT_AMPL_WIDTH - 1),
		7307 => to_unsigned(21123, LUT_AMPL_WIDTH - 1),
		7308 => to_unsigned(21125, LUT_AMPL_WIDTH - 1),
		7309 => to_unsigned(21128, LUT_AMPL_WIDTH - 1),
		7310 => to_unsigned(21130, LUT_AMPL_WIDTH - 1),
		7311 => to_unsigned(21132, LUT_AMPL_WIDTH - 1),
		7312 => to_unsigned(21135, LUT_AMPL_WIDTH - 1),
		7313 => to_unsigned(21137, LUT_AMPL_WIDTH - 1),
		7314 => to_unsigned(21140, LUT_AMPL_WIDTH - 1),
		7315 => to_unsigned(21142, LUT_AMPL_WIDTH - 1),
		7316 => to_unsigned(21144, LUT_AMPL_WIDTH - 1),
		7317 => to_unsigned(21147, LUT_AMPL_WIDTH - 1),
		7318 => to_unsigned(21149, LUT_AMPL_WIDTH - 1),
		7319 => to_unsigned(21152, LUT_AMPL_WIDTH - 1),
		7320 => to_unsigned(21154, LUT_AMPL_WIDTH - 1),
		7321 => to_unsigned(21156, LUT_AMPL_WIDTH - 1),
		7322 => to_unsigned(21159, LUT_AMPL_WIDTH - 1),
		7323 => to_unsigned(21161, LUT_AMPL_WIDTH - 1),
		7324 => to_unsigned(21164, LUT_AMPL_WIDTH - 1),
		7325 => to_unsigned(21166, LUT_AMPL_WIDTH - 1),
		7326 => to_unsigned(21168, LUT_AMPL_WIDTH - 1),
		7327 => to_unsigned(21171, LUT_AMPL_WIDTH - 1),
		7328 => to_unsigned(21173, LUT_AMPL_WIDTH - 1),
		7329 => to_unsigned(21176, LUT_AMPL_WIDTH - 1),
		7330 => to_unsigned(21178, LUT_AMPL_WIDTH - 1),
		7331 => to_unsigned(21180, LUT_AMPL_WIDTH - 1),
		7332 => to_unsigned(21183, LUT_AMPL_WIDTH - 1),
		7333 => to_unsigned(21185, LUT_AMPL_WIDTH - 1),
		7334 => to_unsigned(21188, LUT_AMPL_WIDTH - 1),
		7335 => to_unsigned(21190, LUT_AMPL_WIDTH - 1),
		7336 => to_unsigned(21192, LUT_AMPL_WIDTH - 1),
		7337 => to_unsigned(21195, LUT_AMPL_WIDTH - 1),
		7338 => to_unsigned(21197, LUT_AMPL_WIDTH - 1),
		7339 => to_unsigned(21200, LUT_AMPL_WIDTH - 1),
		7340 => to_unsigned(21202, LUT_AMPL_WIDTH - 1),
		7341 => to_unsigned(21204, LUT_AMPL_WIDTH - 1),
		7342 => to_unsigned(21207, LUT_AMPL_WIDTH - 1),
		7343 => to_unsigned(21209, LUT_AMPL_WIDTH - 1),
		7344 => to_unsigned(21212, LUT_AMPL_WIDTH - 1),
		7345 => to_unsigned(21214, LUT_AMPL_WIDTH - 1),
		7346 => to_unsigned(21216, LUT_AMPL_WIDTH - 1),
		7347 => to_unsigned(21219, LUT_AMPL_WIDTH - 1),
		7348 => to_unsigned(21221, LUT_AMPL_WIDTH - 1),
		7349 => to_unsigned(21224, LUT_AMPL_WIDTH - 1),
		7350 => to_unsigned(21226, LUT_AMPL_WIDTH - 1),
		7351 => to_unsigned(21228, LUT_AMPL_WIDTH - 1),
		7352 => to_unsigned(21231, LUT_AMPL_WIDTH - 1),
		7353 => to_unsigned(21233, LUT_AMPL_WIDTH - 1),
		7354 => to_unsigned(21236, LUT_AMPL_WIDTH - 1),
		7355 => to_unsigned(21238, LUT_AMPL_WIDTH - 1),
		7356 => to_unsigned(21240, LUT_AMPL_WIDTH - 1),
		7357 => to_unsigned(21243, LUT_AMPL_WIDTH - 1),
		7358 => to_unsigned(21245, LUT_AMPL_WIDTH - 1),
		7359 => to_unsigned(21247, LUT_AMPL_WIDTH - 1),
		7360 => to_unsigned(21250, LUT_AMPL_WIDTH - 1),
		7361 => to_unsigned(21252, LUT_AMPL_WIDTH - 1),
		7362 => to_unsigned(21255, LUT_AMPL_WIDTH - 1),
		7363 => to_unsigned(21257, LUT_AMPL_WIDTH - 1),
		7364 => to_unsigned(21259, LUT_AMPL_WIDTH - 1),
		7365 => to_unsigned(21262, LUT_AMPL_WIDTH - 1),
		7366 => to_unsigned(21264, LUT_AMPL_WIDTH - 1),
		7367 => to_unsigned(21267, LUT_AMPL_WIDTH - 1),
		7368 => to_unsigned(21269, LUT_AMPL_WIDTH - 1),
		7369 => to_unsigned(21271, LUT_AMPL_WIDTH - 1),
		7370 => to_unsigned(21274, LUT_AMPL_WIDTH - 1),
		7371 => to_unsigned(21276, LUT_AMPL_WIDTH - 1),
		7372 => to_unsigned(21279, LUT_AMPL_WIDTH - 1),
		7373 => to_unsigned(21281, LUT_AMPL_WIDTH - 1),
		7374 => to_unsigned(21283, LUT_AMPL_WIDTH - 1),
		7375 => to_unsigned(21286, LUT_AMPL_WIDTH - 1),
		7376 => to_unsigned(21288, LUT_AMPL_WIDTH - 1),
		7377 => to_unsigned(21290, LUT_AMPL_WIDTH - 1),
		7378 => to_unsigned(21293, LUT_AMPL_WIDTH - 1),
		7379 => to_unsigned(21295, LUT_AMPL_WIDTH - 1),
		7380 => to_unsigned(21298, LUT_AMPL_WIDTH - 1),
		7381 => to_unsigned(21300, LUT_AMPL_WIDTH - 1),
		7382 => to_unsigned(21302, LUT_AMPL_WIDTH - 1),
		7383 => to_unsigned(21305, LUT_AMPL_WIDTH - 1),
		7384 => to_unsigned(21307, LUT_AMPL_WIDTH - 1),
		7385 => to_unsigned(21310, LUT_AMPL_WIDTH - 1),
		7386 => to_unsigned(21312, LUT_AMPL_WIDTH - 1),
		7387 => to_unsigned(21314, LUT_AMPL_WIDTH - 1),
		7388 => to_unsigned(21317, LUT_AMPL_WIDTH - 1),
		7389 => to_unsigned(21319, LUT_AMPL_WIDTH - 1),
		7390 => to_unsigned(21322, LUT_AMPL_WIDTH - 1),
		7391 => to_unsigned(21324, LUT_AMPL_WIDTH - 1),
		7392 => to_unsigned(21326, LUT_AMPL_WIDTH - 1),
		7393 => to_unsigned(21329, LUT_AMPL_WIDTH - 1),
		7394 => to_unsigned(21331, LUT_AMPL_WIDTH - 1),
		7395 => to_unsigned(21333, LUT_AMPL_WIDTH - 1),
		7396 => to_unsigned(21336, LUT_AMPL_WIDTH - 1),
		7397 => to_unsigned(21338, LUT_AMPL_WIDTH - 1),
		7398 => to_unsigned(21341, LUT_AMPL_WIDTH - 1),
		7399 => to_unsigned(21343, LUT_AMPL_WIDTH - 1),
		7400 => to_unsigned(21345, LUT_AMPL_WIDTH - 1),
		7401 => to_unsigned(21348, LUT_AMPL_WIDTH - 1),
		7402 => to_unsigned(21350, LUT_AMPL_WIDTH - 1),
		7403 => to_unsigned(21353, LUT_AMPL_WIDTH - 1),
		7404 => to_unsigned(21355, LUT_AMPL_WIDTH - 1),
		7405 => to_unsigned(21357, LUT_AMPL_WIDTH - 1),
		7406 => to_unsigned(21360, LUT_AMPL_WIDTH - 1),
		7407 => to_unsigned(21362, LUT_AMPL_WIDTH - 1),
		7408 => to_unsigned(21364, LUT_AMPL_WIDTH - 1),
		7409 => to_unsigned(21367, LUT_AMPL_WIDTH - 1),
		7410 => to_unsigned(21369, LUT_AMPL_WIDTH - 1),
		7411 => to_unsigned(21372, LUT_AMPL_WIDTH - 1),
		7412 => to_unsigned(21374, LUT_AMPL_WIDTH - 1),
		7413 => to_unsigned(21376, LUT_AMPL_WIDTH - 1),
		7414 => to_unsigned(21379, LUT_AMPL_WIDTH - 1),
		7415 => to_unsigned(21381, LUT_AMPL_WIDTH - 1),
		7416 => to_unsigned(21383, LUT_AMPL_WIDTH - 1),
		7417 => to_unsigned(21386, LUT_AMPL_WIDTH - 1),
		7418 => to_unsigned(21388, LUT_AMPL_WIDTH - 1),
		7419 => to_unsigned(21391, LUT_AMPL_WIDTH - 1),
		7420 => to_unsigned(21393, LUT_AMPL_WIDTH - 1),
		7421 => to_unsigned(21395, LUT_AMPL_WIDTH - 1),
		7422 => to_unsigned(21398, LUT_AMPL_WIDTH - 1),
		7423 => to_unsigned(21400, LUT_AMPL_WIDTH - 1),
		7424 => to_unsigned(21403, LUT_AMPL_WIDTH - 1),
		7425 => to_unsigned(21405, LUT_AMPL_WIDTH - 1),
		7426 => to_unsigned(21407, LUT_AMPL_WIDTH - 1),
		7427 => to_unsigned(21410, LUT_AMPL_WIDTH - 1),
		7428 => to_unsigned(21412, LUT_AMPL_WIDTH - 1),
		7429 => to_unsigned(21414, LUT_AMPL_WIDTH - 1),
		7430 => to_unsigned(21417, LUT_AMPL_WIDTH - 1),
		7431 => to_unsigned(21419, LUT_AMPL_WIDTH - 1),
		7432 => to_unsigned(21422, LUT_AMPL_WIDTH - 1),
		7433 => to_unsigned(21424, LUT_AMPL_WIDTH - 1),
		7434 => to_unsigned(21426, LUT_AMPL_WIDTH - 1),
		7435 => to_unsigned(21429, LUT_AMPL_WIDTH - 1),
		7436 => to_unsigned(21431, LUT_AMPL_WIDTH - 1),
		7437 => to_unsigned(21433, LUT_AMPL_WIDTH - 1),
		7438 => to_unsigned(21436, LUT_AMPL_WIDTH - 1),
		7439 => to_unsigned(21438, LUT_AMPL_WIDTH - 1),
		7440 => to_unsigned(21441, LUT_AMPL_WIDTH - 1),
		7441 => to_unsigned(21443, LUT_AMPL_WIDTH - 1),
		7442 => to_unsigned(21445, LUT_AMPL_WIDTH - 1),
		7443 => to_unsigned(21448, LUT_AMPL_WIDTH - 1),
		7444 => to_unsigned(21450, LUT_AMPL_WIDTH - 1),
		7445 => to_unsigned(21452, LUT_AMPL_WIDTH - 1),
		7446 => to_unsigned(21455, LUT_AMPL_WIDTH - 1),
		7447 => to_unsigned(21457, LUT_AMPL_WIDTH - 1),
		7448 => to_unsigned(21460, LUT_AMPL_WIDTH - 1),
		7449 => to_unsigned(21462, LUT_AMPL_WIDTH - 1),
		7450 => to_unsigned(21464, LUT_AMPL_WIDTH - 1),
		7451 => to_unsigned(21467, LUT_AMPL_WIDTH - 1),
		7452 => to_unsigned(21469, LUT_AMPL_WIDTH - 1),
		7453 => to_unsigned(21471, LUT_AMPL_WIDTH - 1),
		7454 => to_unsigned(21474, LUT_AMPL_WIDTH - 1),
		7455 => to_unsigned(21476, LUT_AMPL_WIDTH - 1),
		7456 => to_unsigned(21479, LUT_AMPL_WIDTH - 1),
		7457 => to_unsigned(21481, LUT_AMPL_WIDTH - 1),
		7458 => to_unsigned(21483, LUT_AMPL_WIDTH - 1),
		7459 => to_unsigned(21486, LUT_AMPL_WIDTH - 1),
		7460 => to_unsigned(21488, LUT_AMPL_WIDTH - 1),
		7461 => to_unsigned(21490, LUT_AMPL_WIDTH - 1),
		7462 => to_unsigned(21493, LUT_AMPL_WIDTH - 1),
		7463 => to_unsigned(21495, LUT_AMPL_WIDTH - 1),
		7464 => to_unsigned(21498, LUT_AMPL_WIDTH - 1),
		7465 => to_unsigned(21500, LUT_AMPL_WIDTH - 1),
		7466 => to_unsigned(21502, LUT_AMPL_WIDTH - 1),
		7467 => to_unsigned(21505, LUT_AMPL_WIDTH - 1),
		7468 => to_unsigned(21507, LUT_AMPL_WIDTH - 1),
		7469 => to_unsigned(21509, LUT_AMPL_WIDTH - 1),
		7470 => to_unsigned(21512, LUT_AMPL_WIDTH - 1),
		7471 => to_unsigned(21514, LUT_AMPL_WIDTH - 1),
		7472 => to_unsigned(21516, LUT_AMPL_WIDTH - 1),
		7473 => to_unsigned(21519, LUT_AMPL_WIDTH - 1),
		7474 => to_unsigned(21521, LUT_AMPL_WIDTH - 1),
		7475 => to_unsigned(21524, LUT_AMPL_WIDTH - 1),
		7476 => to_unsigned(21526, LUT_AMPL_WIDTH - 1),
		7477 => to_unsigned(21528, LUT_AMPL_WIDTH - 1),
		7478 => to_unsigned(21531, LUT_AMPL_WIDTH - 1),
		7479 => to_unsigned(21533, LUT_AMPL_WIDTH - 1),
		7480 => to_unsigned(21535, LUT_AMPL_WIDTH - 1),
		7481 => to_unsigned(21538, LUT_AMPL_WIDTH - 1),
		7482 => to_unsigned(21540, LUT_AMPL_WIDTH - 1),
		7483 => to_unsigned(21543, LUT_AMPL_WIDTH - 1),
		7484 => to_unsigned(21545, LUT_AMPL_WIDTH - 1),
		7485 => to_unsigned(21547, LUT_AMPL_WIDTH - 1),
		7486 => to_unsigned(21550, LUT_AMPL_WIDTH - 1),
		7487 => to_unsigned(21552, LUT_AMPL_WIDTH - 1),
		7488 => to_unsigned(21554, LUT_AMPL_WIDTH - 1),
		7489 => to_unsigned(21557, LUT_AMPL_WIDTH - 1),
		7490 => to_unsigned(21559, LUT_AMPL_WIDTH - 1),
		7491 => to_unsigned(21561, LUT_AMPL_WIDTH - 1),
		7492 => to_unsigned(21564, LUT_AMPL_WIDTH - 1),
		7493 => to_unsigned(21566, LUT_AMPL_WIDTH - 1),
		7494 => to_unsigned(21569, LUT_AMPL_WIDTH - 1),
		7495 => to_unsigned(21571, LUT_AMPL_WIDTH - 1),
		7496 => to_unsigned(21573, LUT_AMPL_WIDTH - 1),
		7497 => to_unsigned(21576, LUT_AMPL_WIDTH - 1),
		7498 => to_unsigned(21578, LUT_AMPL_WIDTH - 1),
		7499 => to_unsigned(21580, LUT_AMPL_WIDTH - 1),
		7500 => to_unsigned(21583, LUT_AMPL_WIDTH - 1),
		7501 => to_unsigned(21585, LUT_AMPL_WIDTH - 1),
		7502 => to_unsigned(21587, LUT_AMPL_WIDTH - 1),
		7503 => to_unsigned(21590, LUT_AMPL_WIDTH - 1),
		7504 => to_unsigned(21592, LUT_AMPL_WIDTH - 1),
		7505 => to_unsigned(21595, LUT_AMPL_WIDTH - 1),
		7506 => to_unsigned(21597, LUT_AMPL_WIDTH - 1),
		7507 => to_unsigned(21599, LUT_AMPL_WIDTH - 1),
		7508 => to_unsigned(21602, LUT_AMPL_WIDTH - 1),
		7509 => to_unsigned(21604, LUT_AMPL_WIDTH - 1),
		7510 => to_unsigned(21606, LUT_AMPL_WIDTH - 1),
		7511 => to_unsigned(21609, LUT_AMPL_WIDTH - 1),
		7512 => to_unsigned(21611, LUT_AMPL_WIDTH - 1),
		7513 => to_unsigned(21613, LUT_AMPL_WIDTH - 1),
		7514 => to_unsigned(21616, LUT_AMPL_WIDTH - 1),
		7515 => to_unsigned(21618, LUT_AMPL_WIDTH - 1),
		7516 => to_unsigned(21621, LUT_AMPL_WIDTH - 1),
		7517 => to_unsigned(21623, LUT_AMPL_WIDTH - 1),
		7518 => to_unsigned(21625, LUT_AMPL_WIDTH - 1),
		7519 => to_unsigned(21628, LUT_AMPL_WIDTH - 1),
		7520 => to_unsigned(21630, LUT_AMPL_WIDTH - 1),
		7521 => to_unsigned(21632, LUT_AMPL_WIDTH - 1),
		7522 => to_unsigned(21635, LUT_AMPL_WIDTH - 1),
		7523 => to_unsigned(21637, LUT_AMPL_WIDTH - 1),
		7524 => to_unsigned(21639, LUT_AMPL_WIDTH - 1),
		7525 => to_unsigned(21642, LUT_AMPL_WIDTH - 1),
		7526 => to_unsigned(21644, LUT_AMPL_WIDTH - 1),
		7527 => to_unsigned(21646, LUT_AMPL_WIDTH - 1),
		7528 => to_unsigned(21649, LUT_AMPL_WIDTH - 1),
		7529 => to_unsigned(21651, LUT_AMPL_WIDTH - 1),
		7530 => to_unsigned(21654, LUT_AMPL_WIDTH - 1),
		7531 => to_unsigned(21656, LUT_AMPL_WIDTH - 1),
		7532 => to_unsigned(21658, LUT_AMPL_WIDTH - 1),
		7533 => to_unsigned(21661, LUT_AMPL_WIDTH - 1),
		7534 => to_unsigned(21663, LUT_AMPL_WIDTH - 1),
		7535 => to_unsigned(21665, LUT_AMPL_WIDTH - 1),
		7536 => to_unsigned(21668, LUT_AMPL_WIDTH - 1),
		7537 => to_unsigned(21670, LUT_AMPL_WIDTH - 1),
		7538 => to_unsigned(21672, LUT_AMPL_WIDTH - 1),
		7539 => to_unsigned(21675, LUT_AMPL_WIDTH - 1),
		7540 => to_unsigned(21677, LUT_AMPL_WIDTH - 1),
		7541 => to_unsigned(21679, LUT_AMPL_WIDTH - 1),
		7542 => to_unsigned(21682, LUT_AMPL_WIDTH - 1),
		7543 => to_unsigned(21684, LUT_AMPL_WIDTH - 1),
		7544 => to_unsigned(21687, LUT_AMPL_WIDTH - 1),
		7545 => to_unsigned(21689, LUT_AMPL_WIDTH - 1),
		7546 => to_unsigned(21691, LUT_AMPL_WIDTH - 1),
		7547 => to_unsigned(21694, LUT_AMPL_WIDTH - 1),
		7548 => to_unsigned(21696, LUT_AMPL_WIDTH - 1),
		7549 => to_unsigned(21698, LUT_AMPL_WIDTH - 1),
		7550 => to_unsigned(21701, LUT_AMPL_WIDTH - 1),
		7551 => to_unsigned(21703, LUT_AMPL_WIDTH - 1),
		7552 => to_unsigned(21705, LUT_AMPL_WIDTH - 1),
		7553 => to_unsigned(21708, LUT_AMPL_WIDTH - 1),
		7554 => to_unsigned(21710, LUT_AMPL_WIDTH - 1),
		7555 => to_unsigned(21712, LUT_AMPL_WIDTH - 1),
		7556 => to_unsigned(21715, LUT_AMPL_WIDTH - 1),
		7557 => to_unsigned(21717, LUT_AMPL_WIDTH - 1),
		7558 => to_unsigned(21719, LUT_AMPL_WIDTH - 1),
		7559 => to_unsigned(21722, LUT_AMPL_WIDTH - 1),
		7560 => to_unsigned(21724, LUT_AMPL_WIDTH - 1),
		7561 => to_unsigned(21727, LUT_AMPL_WIDTH - 1),
		7562 => to_unsigned(21729, LUT_AMPL_WIDTH - 1),
		7563 => to_unsigned(21731, LUT_AMPL_WIDTH - 1),
		7564 => to_unsigned(21734, LUT_AMPL_WIDTH - 1),
		7565 => to_unsigned(21736, LUT_AMPL_WIDTH - 1),
		7566 => to_unsigned(21738, LUT_AMPL_WIDTH - 1),
		7567 => to_unsigned(21741, LUT_AMPL_WIDTH - 1),
		7568 => to_unsigned(21743, LUT_AMPL_WIDTH - 1),
		7569 => to_unsigned(21745, LUT_AMPL_WIDTH - 1),
		7570 => to_unsigned(21748, LUT_AMPL_WIDTH - 1),
		7571 => to_unsigned(21750, LUT_AMPL_WIDTH - 1),
		7572 => to_unsigned(21752, LUT_AMPL_WIDTH - 1),
		7573 => to_unsigned(21755, LUT_AMPL_WIDTH - 1),
		7574 => to_unsigned(21757, LUT_AMPL_WIDTH - 1),
		7575 => to_unsigned(21759, LUT_AMPL_WIDTH - 1),
		7576 => to_unsigned(21762, LUT_AMPL_WIDTH - 1),
		7577 => to_unsigned(21764, LUT_AMPL_WIDTH - 1),
		7578 => to_unsigned(21766, LUT_AMPL_WIDTH - 1),
		7579 => to_unsigned(21769, LUT_AMPL_WIDTH - 1),
		7580 => to_unsigned(21771, LUT_AMPL_WIDTH - 1),
		7581 => to_unsigned(21774, LUT_AMPL_WIDTH - 1),
		7582 => to_unsigned(21776, LUT_AMPL_WIDTH - 1),
		7583 => to_unsigned(21778, LUT_AMPL_WIDTH - 1),
		7584 => to_unsigned(21781, LUT_AMPL_WIDTH - 1),
		7585 => to_unsigned(21783, LUT_AMPL_WIDTH - 1),
		7586 => to_unsigned(21785, LUT_AMPL_WIDTH - 1),
		7587 => to_unsigned(21788, LUT_AMPL_WIDTH - 1),
		7588 => to_unsigned(21790, LUT_AMPL_WIDTH - 1),
		7589 => to_unsigned(21792, LUT_AMPL_WIDTH - 1),
		7590 => to_unsigned(21795, LUT_AMPL_WIDTH - 1),
		7591 => to_unsigned(21797, LUT_AMPL_WIDTH - 1),
		7592 => to_unsigned(21799, LUT_AMPL_WIDTH - 1),
		7593 => to_unsigned(21802, LUT_AMPL_WIDTH - 1),
		7594 => to_unsigned(21804, LUT_AMPL_WIDTH - 1),
		7595 => to_unsigned(21806, LUT_AMPL_WIDTH - 1),
		7596 => to_unsigned(21809, LUT_AMPL_WIDTH - 1),
		7597 => to_unsigned(21811, LUT_AMPL_WIDTH - 1),
		7598 => to_unsigned(21813, LUT_AMPL_WIDTH - 1),
		7599 => to_unsigned(21816, LUT_AMPL_WIDTH - 1),
		7600 => to_unsigned(21818, LUT_AMPL_WIDTH - 1),
		7601 => to_unsigned(21820, LUT_AMPL_WIDTH - 1),
		7602 => to_unsigned(21823, LUT_AMPL_WIDTH - 1),
		7603 => to_unsigned(21825, LUT_AMPL_WIDTH - 1),
		7604 => to_unsigned(21827, LUT_AMPL_WIDTH - 1),
		7605 => to_unsigned(21830, LUT_AMPL_WIDTH - 1),
		7606 => to_unsigned(21832, LUT_AMPL_WIDTH - 1),
		7607 => to_unsigned(21835, LUT_AMPL_WIDTH - 1),
		7608 => to_unsigned(21837, LUT_AMPL_WIDTH - 1),
		7609 => to_unsigned(21839, LUT_AMPL_WIDTH - 1),
		7610 => to_unsigned(21842, LUT_AMPL_WIDTH - 1),
		7611 => to_unsigned(21844, LUT_AMPL_WIDTH - 1),
		7612 => to_unsigned(21846, LUT_AMPL_WIDTH - 1),
		7613 => to_unsigned(21849, LUT_AMPL_WIDTH - 1),
		7614 => to_unsigned(21851, LUT_AMPL_WIDTH - 1),
		7615 => to_unsigned(21853, LUT_AMPL_WIDTH - 1),
		7616 => to_unsigned(21856, LUT_AMPL_WIDTH - 1),
		7617 => to_unsigned(21858, LUT_AMPL_WIDTH - 1),
		7618 => to_unsigned(21860, LUT_AMPL_WIDTH - 1),
		7619 => to_unsigned(21863, LUT_AMPL_WIDTH - 1),
		7620 => to_unsigned(21865, LUT_AMPL_WIDTH - 1),
		7621 => to_unsigned(21867, LUT_AMPL_WIDTH - 1),
		7622 => to_unsigned(21870, LUT_AMPL_WIDTH - 1),
		7623 => to_unsigned(21872, LUT_AMPL_WIDTH - 1),
		7624 => to_unsigned(21874, LUT_AMPL_WIDTH - 1),
		7625 => to_unsigned(21877, LUT_AMPL_WIDTH - 1),
		7626 => to_unsigned(21879, LUT_AMPL_WIDTH - 1),
		7627 => to_unsigned(21881, LUT_AMPL_WIDTH - 1),
		7628 => to_unsigned(21884, LUT_AMPL_WIDTH - 1),
		7629 => to_unsigned(21886, LUT_AMPL_WIDTH - 1),
		7630 => to_unsigned(21888, LUT_AMPL_WIDTH - 1),
		7631 => to_unsigned(21891, LUT_AMPL_WIDTH - 1),
		7632 => to_unsigned(21893, LUT_AMPL_WIDTH - 1),
		7633 => to_unsigned(21895, LUT_AMPL_WIDTH - 1),
		7634 => to_unsigned(21898, LUT_AMPL_WIDTH - 1),
		7635 => to_unsigned(21900, LUT_AMPL_WIDTH - 1),
		7636 => to_unsigned(21902, LUT_AMPL_WIDTH - 1),
		7637 => to_unsigned(21905, LUT_AMPL_WIDTH - 1),
		7638 => to_unsigned(21907, LUT_AMPL_WIDTH - 1),
		7639 => to_unsigned(21909, LUT_AMPL_WIDTH - 1),
		7640 => to_unsigned(21912, LUT_AMPL_WIDTH - 1),
		7641 => to_unsigned(21914, LUT_AMPL_WIDTH - 1),
		7642 => to_unsigned(21916, LUT_AMPL_WIDTH - 1),
		7643 => to_unsigned(21919, LUT_AMPL_WIDTH - 1),
		7644 => to_unsigned(21921, LUT_AMPL_WIDTH - 1),
		7645 => to_unsigned(21923, LUT_AMPL_WIDTH - 1),
		7646 => to_unsigned(21926, LUT_AMPL_WIDTH - 1),
		7647 => to_unsigned(21928, LUT_AMPL_WIDTH - 1),
		7648 => to_unsigned(21930, LUT_AMPL_WIDTH - 1),
		7649 => to_unsigned(21933, LUT_AMPL_WIDTH - 1),
		7650 => to_unsigned(21935, LUT_AMPL_WIDTH - 1),
		7651 => to_unsigned(21937, LUT_AMPL_WIDTH - 1),
		7652 => to_unsigned(21940, LUT_AMPL_WIDTH - 1),
		7653 => to_unsigned(21942, LUT_AMPL_WIDTH - 1),
		7654 => to_unsigned(21944, LUT_AMPL_WIDTH - 1),
		7655 => to_unsigned(21947, LUT_AMPL_WIDTH - 1),
		7656 => to_unsigned(21949, LUT_AMPL_WIDTH - 1),
		7657 => to_unsigned(21951, LUT_AMPL_WIDTH - 1),
		7658 => to_unsigned(21954, LUT_AMPL_WIDTH - 1),
		7659 => to_unsigned(21956, LUT_AMPL_WIDTH - 1),
		7660 => to_unsigned(21958, LUT_AMPL_WIDTH - 1),
		7661 => to_unsigned(21961, LUT_AMPL_WIDTH - 1),
		7662 => to_unsigned(21963, LUT_AMPL_WIDTH - 1),
		7663 => to_unsigned(21965, LUT_AMPL_WIDTH - 1),
		7664 => to_unsigned(21968, LUT_AMPL_WIDTH - 1),
		7665 => to_unsigned(21970, LUT_AMPL_WIDTH - 1),
		7666 => to_unsigned(21972, LUT_AMPL_WIDTH - 1),
		7667 => to_unsigned(21975, LUT_AMPL_WIDTH - 1),
		7668 => to_unsigned(21977, LUT_AMPL_WIDTH - 1),
		7669 => to_unsigned(21979, LUT_AMPL_WIDTH - 1),
		7670 => to_unsigned(21982, LUT_AMPL_WIDTH - 1),
		7671 => to_unsigned(21984, LUT_AMPL_WIDTH - 1),
		7672 => to_unsigned(21986, LUT_AMPL_WIDTH - 1),
		7673 => to_unsigned(21989, LUT_AMPL_WIDTH - 1),
		7674 => to_unsigned(21991, LUT_AMPL_WIDTH - 1),
		7675 => to_unsigned(21993, LUT_AMPL_WIDTH - 1),
		7676 => to_unsigned(21996, LUT_AMPL_WIDTH - 1),
		7677 => to_unsigned(21998, LUT_AMPL_WIDTH - 1),
		7678 => to_unsigned(22000, LUT_AMPL_WIDTH - 1),
		7679 => to_unsigned(22003, LUT_AMPL_WIDTH - 1),
		7680 => to_unsigned(22005, LUT_AMPL_WIDTH - 1),
		7681 => to_unsigned(22007, LUT_AMPL_WIDTH - 1),
		7682 => to_unsigned(22010, LUT_AMPL_WIDTH - 1),
		7683 => to_unsigned(22012, LUT_AMPL_WIDTH - 1),
		7684 => to_unsigned(22014, LUT_AMPL_WIDTH - 1),
		7685 => to_unsigned(22017, LUT_AMPL_WIDTH - 1),
		7686 => to_unsigned(22019, LUT_AMPL_WIDTH - 1),
		7687 => to_unsigned(22021, LUT_AMPL_WIDTH - 1),
		7688 => to_unsigned(22024, LUT_AMPL_WIDTH - 1),
		7689 => to_unsigned(22026, LUT_AMPL_WIDTH - 1),
		7690 => to_unsigned(22028, LUT_AMPL_WIDTH - 1),
		7691 => to_unsigned(22031, LUT_AMPL_WIDTH - 1),
		7692 => to_unsigned(22033, LUT_AMPL_WIDTH - 1),
		7693 => to_unsigned(22035, LUT_AMPL_WIDTH - 1),
		7694 => to_unsigned(22038, LUT_AMPL_WIDTH - 1),
		7695 => to_unsigned(22040, LUT_AMPL_WIDTH - 1),
		7696 => to_unsigned(22042, LUT_AMPL_WIDTH - 1),
		7697 => to_unsigned(22045, LUT_AMPL_WIDTH - 1),
		7698 => to_unsigned(22047, LUT_AMPL_WIDTH - 1),
		7699 => to_unsigned(22049, LUT_AMPL_WIDTH - 1),
		7700 => to_unsigned(22051, LUT_AMPL_WIDTH - 1),
		7701 => to_unsigned(22054, LUT_AMPL_WIDTH - 1),
		7702 => to_unsigned(22056, LUT_AMPL_WIDTH - 1),
		7703 => to_unsigned(22058, LUT_AMPL_WIDTH - 1),
		7704 => to_unsigned(22061, LUT_AMPL_WIDTH - 1),
		7705 => to_unsigned(22063, LUT_AMPL_WIDTH - 1),
		7706 => to_unsigned(22065, LUT_AMPL_WIDTH - 1),
		7707 => to_unsigned(22068, LUT_AMPL_WIDTH - 1),
		7708 => to_unsigned(22070, LUT_AMPL_WIDTH - 1),
		7709 => to_unsigned(22072, LUT_AMPL_WIDTH - 1),
		7710 => to_unsigned(22075, LUT_AMPL_WIDTH - 1),
		7711 => to_unsigned(22077, LUT_AMPL_WIDTH - 1),
		7712 => to_unsigned(22079, LUT_AMPL_WIDTH - 1),
		7713 => to_unsigned(22082, LUT_AMPL_WIDTH - 1),
		7714 => to_unsigned(22084, LUT_AMPL_WIDTH - 1),
		7715 => to_unsigned(22086, LUT_AMPL_WIDTH - 1),
		7716 => to_unsigned(22089, LUT_AMPL_WIDTH - 1),
		7717 => to_unsigned(22091, LUT_AMPL_WIDTH - 1),
		7718 => to_unsigned(22093, LUT_AMPL_WIDTH - 1),
		7719 => to_unsigned(22096, LUT_AMPL_WIDTH - 1),
		7720 => to_unsigned(22098, LUT_AMPL_WIDTH - 1),
		7721 => to_unsigned(22100, LUT_AMPL_WIDTH - 1),
		7722 => to_unsigned(22103, LUT_AMPL_WIDTH - 1),
		7723 => to_unsigned(22105, LUT_AMPL_WIDTH - 1),
		7724 => to_unsigned(22107, LUT_AMPL_WIDTH - 1),
		7725 => to_unsigned(22110, LUT_AMPL_WIDTH - 1),
		7726 => to_unsigned(22112, LUT_AMPL_WIDTH - 1),
		7727 => to_unsigned(22114, LUT_AMPL_WIDTH - 1),
		7728 => to_unsigned(22116, LUT_AMPL_WIDTH - 1),
		7729 => to_unsigned(22119, LUT_AMPL_WIDTH - 1),
		7730 => to_unsigned(22121, LUT_AMPL_WIDTH - 1),
		7731 => to_unsigned(22123, LUT_AMPL_WIDTH - 1),
		7732 => to_unsigned(22126, LUT_AMPL_WIDTH - 1),
		7733 => to_unsigned(22128, LUT_AMPL_WIDTH - 1),
		7734 => to_unsigned(22130, LUT_AMPL_WIDTH - 1),
		7735 => to_unsigned(22133, LUT_AMPL_WIDTH - 1),
		7736 => to_unsigned(22135, LUT_AMPL_WIDTH - 1),
		7737 => to_unsigned(22137, LUT_AMPL_WIDTH - 1),
		7738 => to_unsigned(22140, LUT_AMPL_WIDTH - 1),
		7739 => to_unsigned(22142, LUT_AMPL_WIDTH - 1),
		7740 => to_unsigned(22144, LUT_AMPL_WIDTH - 1),
		7741 => to_unsigned(22147, LUT_AMPL_WIDTH - 1),
		7742 => to_unsigned(22149, LUT_AMPL_WIDTH - 1),
		7743 => to_unsigned(22151, LUT_AMPL_WIDTH - 1),
		7744 => to_unsigned(22154, LUT_AMPL_WIDTH - 1),
		7745 => to_unsigned(22156, LUT_AMPL_WIDTH - 1),
		7746 => to_unsigned(22158, LUT_AMPL_WIDTH - 1),
		7747 => to_unsigned(22160, LUT_AMPL_WIDTH - 1),
		7748 => to_unsigned(22163, LUT_AMPL_WIDTH - 1),
		7749 => to_unsigned(22165, LUT_AMPL_WIDTH - 1),
		7750 => to_unsigned(22167, LUT_AMPL_WIDTH - 1),
		7751 => to_unsigned(22170, LUT_AMPL_WIDTH - 1),
		7752 => to_unsigned(22172, LUT_AMPL_WIDTH - 1),
		7753 => to_unsigned(22174, LUT_AMPL_WIDTH - 1),
		7754 => to_unsigned(22177, LUT_AMPL_WIDTH - 1),
		7755 => to_unsigned(22179, LUT_AMPL_WIDTH - 1),
		7756 => to_unsigned(22181, LUT_AMPL_WIDTH - 1),
		7757 => to_unsigned(22184, LUT_AMPL_WIDTH - 1),
		7758 => to_unsigned(22186, LUT_AMPL_WIDTH - 1),
		7759 => to_unsigned(22188, LUT_AMPL_WIDTH - 1),
		7760 => to_unsigned(22191, LUT_AMPL_WIDTH - 1),
		7761 => to_unsigned(22193, LUT_AMPL_WIDTH - 1),
		7762 => to_unsigned(22195, LUT_AMPL_WIDTH - 1),
		7763 => to_unsigned(22197, LUT_AMPL_WIDTH - 1),
		7764 => to_unsigned(22200, LUT_AMPL_WIDTH - 1),
		7765 => to_unsigned(22202, LUT_AMPL_WIDTH - 1),
		7766 => to_unsigned(22204, LUT_AMPL_WIDTH - 1),
		7767 => to_unsigned(22207, LUT_AMPL_WIDTH - 1),
		7768 => to_unsigned(22209, LUT_AMPL_WIDTH - 1),
		7769 => to_unsigned(22211, LUT_AMPL_WIDTH - 1),
		7770 => to_unsigned(22214, LUT_AMPL_WIDTH - 1),
		7771 => to_unsigned(22216, LUT_AMPL_WIDTH - 1),
		7772 => to_unsigned(22218, LUT_AMPL_WIDTH - 1),
		7773 => to_unsigned(22221, LUT_AMPL_WIDTH - 1),
		7774 => to_unsigned(22223, LUT_AMPL_WIDTH - 1),
		7775 => to_unsigned(22225, LUT_AMPL_WIDTH - 1),
		7776 => to_unsigned(22227, LUT_AMPL_WIDTH - 1),
		7777 => to_unsigned(22230, LUT_AMPL_WIDTH - 1),
		7778 => to_unsigned(22232, LUT_AMPL_WIDTH - 1),
		7779 => to_unsigned(22234, LUT_AMPL_WIDTH - 1),
		7780 => to_unsigned(22237, LUT_AMPL_WIDTH - 1),
		7781 => to_unsigned(22239, LUT_AMPL_WIDTH - 1),
		7782 => to_unsigned(22241, LUT_AMPL_WIDTH - 1),
		7783 => to_unsigned(22244, LUT_AMPL_WIDTH - 1),
		7784 => to_unsigned(22246, LUT_AMPL_WIDTH - 1),
		7785 => to_unsigned(22248, LUT_AMPL_WIDTH - 1),
		7786 => to_unsigned(22251, LUT_AMPL_WIDTH - 1),
		7787 => to_unsigned(22253, LUT_AMPL_WIDTH - 1),
		7788 => to_unsigned(22255, LUT_AMPL_WIDTH - 1),
		7789 => to_unsigned(22257, LUT_AMPL_WIDTH - 1),
		7790 => to_unsigned(22260, LUT_AMPL_WIDTH - 1),
		7791 => to_unsigned(22262, LUT_AMPL_WIDTH - 1),
		7792 => to_unsigned(22264, LUT_AMPL_WIDTH - 1),
		7793 => to_unsigned(22267, LUT_AMPL_WIDTH - 1),
		7794 => to_unsigned(22269, LUT_AMPL_WIDTH - 1),
		7795 => to_unsigned(22271, LUT_AMPL_WIDTH - 1),
		7796 => to_unsigned(22274, LUT_AMPL_WIDTH - 1),
		7797 => to_unsigned(22276, LUT_AMPL_WIDTH - 1),
		7798 => to_unsigned(22278, LUT_AMPL_WIDTH - 1),
		7799 => to_unsigned(22281, LUT_AMPL_WIDTH - 1),
		7800 => to_unsigned(22283, LUT_AMPL_WIDTH - 1),
		7801 => to_unsigned(22285, LUT_AMPL_WIDTH - 1),
		7802 => to_unsigned(22287, LUT_AMPL_WIDTH - 1),
		7803 => to_unsigned(22290, LUT_AMPL_WIDTH - 1),
		7804 => to_unsigned(22292, LUT_AMPL_WIDTH - 1),
		7805 => to_unsigned(22294, LUT_AMPL_WIDTH - 1),
		7806 => to_unsigned(22297, LUT_AMPL_WIDTH - 1),
		7807 => to_unsigned(22299, LUT_AMPL_WIDTH - 1),
		7808 => to_unsigned(22301, LUT_AMPL_WIDTH - 1),
		7809 => to_unsigned(22304, LUT_AMPL_WIDTH - 1),
		7810 => to_unsigned(22306, LUT_AMPL_WIDTH - 1),
		7811 => to_unsigned(22308, LUT_AMPL_WIDTH - 1),
		7812 => to_unsigned(22310, LUT_AMPL_WIDTH - 1),
		7813 => to_unsigned(22313, LUT_AMPL_WIDTH - 1),
		7814 => to_unsigned(22315, LUT_AMPL_WIDTH - 1),
		7815 => to_unsigned(22317, LUT_AMPL_WIDTH - 1),
		7816 => to_unsigned(22320, LUT_AMPL_WIDTH - 1),
		7817 => to_unsigned(22322, LUT_AMPL_WIDTH - 1),
		7818 => to_unsigned(22324, LUT_AMPL_WIDTH - 1),
		7819 => to_unsigned(22327, LUT_AMPL_WIDTH - 1),
		7820 => to_unsigned(22329, LUT_AMPL_WIDTH - 1),
		7821 => to_unsigned(22331, LUT_AMPL_WIDTH - 1),
		7822 => to_unsigned(22333, LUT_AMPL_WIDTH - 1),
		7823 => to_unsigned(22336, LUT_AMPL_WIDTH - 1),
		7824 => to_unsigned(22338, LUT_AMPL_WIDTH - 1),
		7825 => to_unsigned(22340, LUT_AMPL_WIDTH - 1),
		7826 => to_unsigned(22343, LUT_AMPL_WIDTH - 1),
		7827 => to_unsigned(22345, LUT_AMPL_WIDTH - 1),
		7828 => to_unsigned(22347, LUT_AMPL_WIDTH - 1),
		7829 => to_unsigned(22350, LUT_AMPL_WIDTH - 1),
		7830 => to_unsigned(22352, LUT_AMPL_WIDTH - 1),
		7831 => to_unsigned(22354, LUT_AMPL_WIDTH - 1),
		7832 => to_unsigned(22356, LUT_AMPL_WIDTH - 1),
		7833 => to_unsigned(22359, LUT_AMPL_WIDTH - 1),
		7834 => to_unsigned(22361, LUT_AMPL_WIDTH - 1),
		7835 => to_unsigned(22363, LUT_AMPL_WIDTH - 1),
		7836 => to_unsigned(22366, LUT_AMPL_WIDTH - 1),
		7837 => to_unsigned(22368, LUT_AMPL_WIDTH - 1),
		7838 => to_unsigned(22370, LUT_AMPL_WIDTH - 1),
		7839 => to_unsigned(22373, LUT_AMPL_WIDTH - 1),
		7840 => to_unsigned(22375, LUT_AMPL_WIDTH - 1),
		7841 => to_unsigned(22377, LUT_AMPL_WIDTH - 1),
		7842 => to_unsigned(22379, LUT_AMPL_WIDTH - 1),
		7843 => to_unsigned(22382, LUT_AMPL_WIDTH - 1),
		7844 => to_unsigned(22384, LUT_AMPL_WIDTH - 1),
		7845 => to_unsigned(22386, LUT_AMPL_WIDTH - 1),
		7846 => to_unsigned(22389, LUT_AMPL_WIDTH - 1),
		7847 => to_unsigned(22391, LUT_AMPL_WIDTH - 1),
		7848 => to_unsigned(22393, LUT_AMPL_WIDTH - 1),
		7849 => to_unsigned(22395, LUT_AMPL_WIDTH - 1),
		7850 => to_unsigned(22398, LUT_AMPL_WIDTH - 1),
		7851 => to_unsigned(22400, LUT_AMPL_WIDTH - 1),
		7852 => to_unsigned(22402, LUT_AMPL_WIDTH - 1),
		7853 => to_unsigned(22405, LUT_AMPL_WIDTH - 1),
		7854 => to_unsigned(22407, LUT_AMPL_WIDTH - 1),
		7855 => to_unsigned(22409, LUT_AMPL_WIDTH - 1),
		7856 => to_unsigned(22411, LUT_AMPL_WIDTH - 1),
		7857 => to_unsigned(22414, LUT_AMPL_WIDTH - 1),
		7858 => to_unsigned(22416, LUT_AMPL_WIDTH - 1),
		7859 => to_unsigned(22418, LUT_AMPL_WIDTH - 1),
		7860 => to_unsigned(22421, LUT_AMPL_WIDTH - 1),
		7861 => to_unsigned(22423, LUT_AMPL_WIDTH - 1),
		7862 => to_unsigned(22425, LUT_AMPL_WIDTH - 1),
		7863 => to_unsigned(22428, LUT_AMPL_WIDTH - 1),
		7864 => to_unsigned(22430, LUT_AMPL_WIDTH - 1),
		7865 => to_unsigned(22432, LUT_AMPL_WIDTH - 1),
		7866 => to_unsigned(22434, LUT_AMPL_WIDTH - 1),
		7867 => to_unsigned(22437, LUT_AMPL_WIDTH - 1),
		7868 => to_unsigned(22439, LUT_AMPL_WIDTH - 1),
		7869 => to_unsigned(22441, LUT_AMPL_WIDTH - 1),
		7870 => to_unsigned(22444, LUT_AMPL_WIDTH - 1),
		7871 => to_unsigned(22446, LUT_AMPL_WIDTH - 1),
		7872 => to_unsigned(22448, LUT_AMPL_WIDTH - 1),
		7873 => to_unsigned(22450, LUT_AMPL_WIDTH - 1),
		7874 => to_unsigned(22453, LUT_AMPL_WIDTH - 1),
		7875 => to_unsigned(22455, LUT_AMPL_WIDTH - 1),
		7876 => to_unsigned(22457, LUT_AMPL_WIDTH - 1),
		7877 => to_unsigned(22460, LUT_AMPL_WIDTH - 1),
		7878 => to_unsigned(22462, LUT_AMPL_WIDTH - 1),
		7879 => to_unsigned(22464, LUT_AMPL_WIDTH - 1),
		7880 => to_unsigned(22466, LUT_AMPL_WIDTH - 1),
		7881 => to_unsigned(22469, LUT_AMPL_WIDTH - 1),
		7882 => to_unsigned(22471, LUT_AMPL_WIDTH - 1),
		7883 => to_unsigned(22473, LUT_AMPL_WIDTH - 1),
		7884 => to_unsigned(22476, LUT_AMPL_WIDTH - 1),
		7885 => to_unsigned(22478, LUT_AMPL_WIDTH - 1),
		7886 => to_unsigned(22480, LUT_AMPL_WIDTH - 1),
		7887 => to_unsigned(22482, LUT_AMPL_WIDTH - 1),
		7888 => to_unsigned(22485, LUT_AMPL_WIDTH - 1),
		7889 => to_unsigned(22487, LUT_AMPL_WIDTH - 1),
		7890 => to_unsigned(22489, LUT_AMPL_WIDTH - 1),
		7891 => to_unsigned(22492, LUT_AMPL_WIDTH - 1),
		7892 => to_unsigned(22494, LUT_AMPL_WIDTH - 1),
		7893 => to_unsigned(22496, LUT_AMPL_WIDTH - 1),
		7894 => to_unsigned(22498, LUT_AMPL_WIDTH - 1),
		7895 => to_unsigned(22501, LUT_AMPL_WIDTH - 1),
		7896 => to_unsigned(22503, LUT_AMPL_WIDTH - 1),
		7897 => to_unsigned(22505, LUT_AMPL_WIDTH - 1),
		7898 => to_unsigned(22508, LUT_AMPL_WIDTH - 1),
		7899 => to_unsigned(22510, LUT_AMPL_WIDTH - 1),
		7900 => to_unsigned(22512, LUT_AMPL_WIDTH - 1),
		7901 => to_unsigned(22514, LUT_AMPL_WIDTH - 1),
		7902 => to_unsigned(22517, LUT_AMPL_WIDTH - 1),
		7903 => to_unsigned(22519, LUT_AMPL_WIDTH - 1),
		7904 => to_unsigned(22521, LUT_AMPL_WIDTH - 1),
		7905 => to_unsigned(22524, LUT_AMPL_WIDTH - 1),
		7906 => to_unsigned(22526, LUT_AMPL_WIDTH - 1),
		7907 => to_unsigned(22528, LUT_AMPL_WIDTH - 1),
		7908 => to_unsigned(22530, LUT_AMPL_WIDTH - 1),
		7909 => to_unsigned(22533, LUT_AMPL_WIDTH - 1),
		7910 => to_unsigned(22535, LUT_AMPL_WIDTH - 1),
		7911 => to_unsigned(22537, LUT_AMPL_WIDTH - 1),
		7912 => to_unsigned(22540, LUT_AMPL_WIDTH - 1),
		7913 => to_unsigned(22542, LUT_AMPL_WIDTH - 1),
		7914 => to_unsigned(22544, LUT_AMPL_WIDTH - 1),
		7915 => to_unsigned(22546, LUT_AMPL_WIDTH - 1),
		7916 => to_unsigned(22549, LUT_AMPL_WIDTH - 1),
		7917 => to_unsigned(22551, LUT_AMPL_WIDTH - 1),
		7918 => to_unsigned(22553, LUT_AMPL_WIDTH - 1),
		7919 => to_unsigned(22555, LUT_AMPL_WIDTH - 1),
		7920 => to_unsigned(22558, LUT_AMPL_WIDTH - 1),
		7921 => to_unsigned(22560, LUT_AMPL_WIDTH - 1),
		7922 => to_unsigned(22562, LUT_AMPL_WIDTH - 1),
		7923 => to_unsigned(22565, LUT_AMPL_WIDTH - 1),
		7924 => to_unsigned(22567, LUT_AMPL_WIDTH - 1),
		7925 => to_unsigned(22569, LUT_AMPL_WIDTH - 1),
		7926 => to_unsigned(22571, LUT_AMPL_WIDTH - 1),
		7927 => to_unsigned(22574, LUT_AMPL_WIDTH - 1),
		7928 => to_unsigned(22576, LUT_AMPL_WIDTH - 1),
		7929 => to_unsigned(22578, LUT_AMPL_WIDTH - 1),
		7930 => to_unsigned(22581, LUT_AMPL_WIDTH - 1),
		7931 => to_unsigned(22583, LUT_AMPL_WIDTH - 1),
		7932 => to_unsigned(22585, LUT_AMPL_WIDTH - 1),
		7933 => to_unsigned(22587, LUT_AMPL_WIDTH - 1),
		7934 => to_unsigned(22590, LUT_AMPL_WIDTH - 1),
		7935 => to_unsigned(22592, LUT_AMPL_WIDTH - 1),
		7936 => to_unsigned(22594, LUT_AMPL_WIDTH - 1),
		7937 => to_unsigned(22596, LUT_AMPL_WIDTH - 1),
		7938 => to_unsigned(22599, LUT_AMPL_WIDTH - 1),
		7939 => to_unsigned(22601, LUT_AMPL_WIDTH - 1),
		7940 => to_unsigned(22603, LUT_AMPL_WIDTH - 1),
		7941 => to_unsigned(22606, LUT_AMPL_WIDTH - 1),
		7942 => to_unsigned(22608, LUT_AMPL_WIDTH - 1),
		7943 => to_unsigned(22610, LUT_AMPL_WIDTH - 1),
		7944 => to_unsigned(22612, LUT_AMPL_WIDTH - 1),
		7945 => to_unsigned(22615, LUT_AMPL_WIDTH - 1),
		7946 => to_unsigned(22617, LUT_AMPL_WIDTH - 1),
		7947 => to_unsigned(22619, LUT_AMPL_WIDTH - 1),
		7948 => to_unsigned(22621, LUT_AMPL_WIDTH - 1),
		7949 => to_unsigned(22624, LUT_AMPL_WIDTH - 1),
		7950 => to_unsigned(22626, LUT_AMPL_WIDTH - 1),
		7951 => to_unsigned(22628, LUT_AMPL_WIDTH - 1),
		7952 => to_unsigned(22631, LUT_AMPL_WIDTH - 1),
		7953 => to_unsigned(22633, LUT_AMPL_WIDTH - 1),
		7954 => to_unsigned(22635, LUT_AMPL_WIDTH - 1),
		7955 => to_unsigned(22637, LUT_AMPL_WIDTH - 1),
		7956 => to_unsigned(22640, LUT_AMPL_WIDTH - 1),
		7957 => to_unsigned(22642, LUT_AMPL_WIDTH - 1),
		7958 => to_unsigned(22644, LUT_AMPL_WIDTH - 1),
		7959 => to_unsigned(22646, LUT_AMPL_WIDTH - 1),
		7960 => to_unsigned(22649, LUT_AMPL_WIDTH - 1),
		7961 => to_unsigned(22651, LUT_AMPL_WIDTH - 1),
		7962 => to_unsigned(22653, LUT_AMPL_WIDTH - 1),
		7963 => to_unsigned(22656, LUT_AMPL_WIDTH - 1),
		7964 => to_unsigned(22658, LUT_AMPL_WIDTH - 1),
		7965 => to_unsigned(22660, LUT_AMPL_WIDTH - 1),
		7966 => to_unsigned(22662, LUT_AMPL_WIDTH - 1),
		7967 => to_unsigned(22665, LUT_AMPL_WIDTH - 1),
		7968 => to_unsigned(22667, LUT_AMPL_WIDTH - 1),
		7969 => to_unsigned(22669, LUT_AMPL_WIDTH - 1),
		7970 => to_unsigned(22671, LUT_AMPL_WIDTH - 1),
		7971 => to_unsigned(22674, LUT_AMPL_WIDTH - 1),
		7972 => to_unsigned(22676, LUT_AMPL_WIDTH - 1),
		7973 => to_unsigned(22678, LUT_AMPL_WIDTH - 1),
		7974 => to_unsigned(22680, LUT_AMPL_WIDTH - 1),
		7975 => to_unsigned(22683, LUT_AMPL_WIDTH - 1),
		7976 => to_unsigned(22685, LUT_AMPL_WIDTH - 1),
		7977 => to_unsigned(22687, LUT_AMPL_WIDTH - 1),
		7978 => to_unsigned(22690, LUT_AMPL_WIDTH - 1),
		7979 => to_unsigned(22692, LUT_AMPL_WIDTH - 1),
		7980 => to_unsigned(22694, LUT_AMPL_WIDTH - 1),
		7981 => to_unsigned(22696, LUT_AMPL_WIDTH - 1),
		7982 => to_unsigned(22699, LUT_AMPL_WIDTH - 1),
		7983 => to_unsigned(22701, LUT_AMPL_WIDTH - 1),
		7984 => to_unsigned(22703, LUT_AMPL_WIDTH - 1),
		7985 => to_unsigned(22705, LUT_AMPL_WIDTH - 1),
		7986 => to_unsigned(22708, LUT_AMPL_WIDTH - 1),
		7987 => to_unsigned(22710, LUT_AMPL_WIDTH - 1),
		7988 => to_unsigned(22712, LUT_AMPL_WIDTH - 1),
		7989 => to_unsigned(22714, LUT_AMPL_WIDTH - 1),
		7990 => to_unsigned(22717, LUT_AMPL_WIDTH - 1),
		7991 => to_unsigned(22719, LUT_AMPL_WIDTH - 1),
		7992 => to_unsigned(22721, LUT_AMPL_WIDTH - 1),
		7993 => to_unsigned(22724, LUT_AMPL_WIDTH - 1),
		7994 => to_unsigned(22726, LUT_AMPL_WIDTH - 1),
		7995 => to_unsigned(22728, LUT_AMPL_WIDTH - 1),
		7996 => to_unsigned(22730, LUT_AMPL_WIDTH - 1),
		7997 => to_unsigned(22733, LUT_AMPL_WIDTH - 1),
		7998 => to_unsigned(22735, LUT_AMPL_WIDTH - 1),
		7999 => to_unsigned(22737, LUT_AMPL_WIDTH - 1),
		8000 => to_unsigned(22739, LUT_AMPL_WIDTH - 1),
		8001 => to_unsigned(22742, LUT_AMPL_WIDTH - 1),
		8002 => to_unsigned(22744, LUT_AMPL_WIDTH - 1),
		8003 => to_unsigned(22746, LUT_AMPL_WIDTH - 1),
		8004 => to_unsigned(22748, LUT_AMPL_WIDTH - 1),
		8005 => to_unsigned(22751, LUT_AMPL_WIDTH - 1),
		8006 => to_unsigned(22753, LUT_AMPL_WIDTH - 1),
		8007 => to_unsigned(22755, LUT_AMPL_WIDTH - 1),
		8008 => to_unsigned(22757, LUT_AMPL_WIDTH - 1),
		8009 => to_unsigned(22760, LUT_AMPL_WIDTH - 1),
		8010 => to_unsigned(22762, LUT_AMPL_WIDTH - 1),
		8011 => to_unsigned(22764, LUT_AMPL_WIDTH - 1),
		8012 => to_unsigned(22766, LUT_AMPL_WIDTH - 1),
		8013 => to_unsigned(22769, LUT_AMPL_WIDTH - 1),
		8014 => to_unsigned(22771, LUT_AMPL_WIDTH - 1),
		8015 => to_unsigned(22773, LUT_AMPL_WIDTH - 1),
		8016 => to_unsigned(22776, LUT_AMPL_WIDTH - 1),
		8017 => to_unsigned(22778, LUT_AMPL_WIDTH - 1),
		8018 => to_unsigned(22780, LUT_AMPL_WIDTH - 1),
		8019 => to_unsigned(22782, LUT_AMPL_WIDTH - 1),
		8020 => to_unsigned(22785, LUT_AMPL_WIDTH - 1),
		8021 => to_unsigned(22787, LUT_AMPL_WIDTH - 1),
		8022 => to_unsigned(22789, LUT_AMPL_WIDTH - 1),
		8023 => to_unsigned(22791, LUT_AMPL_WIDTH - 1),
		8024 => to_unsigned(22794, LUT_AMPL_WIDTH - 1),
		8025 => to_unsigned(22796, LUT_AMPL_WIDTH - 1),
		8026 => to_unsigned(22798, LUT_AMPL_WIDTH - 1),
		8027 => to_unsigned(22800, LUT_AMPL_WIDTH - 1),
		8028 => to_unsigned(22803, LUT_AMPL_WIDTH - 1),
		8029 => to_unsigned(22805, LUT_AMPL_WIDTH - 1),
		8030 => to_unsigned(22807, LUT_AMPL_WIDTH - 1),
		8031 => to_unsigned(22809, LUT_AMPL_WIDTH - 1),
		8032 => to_unsigned(22812, LUT_AMPL_WIDTH - 1),
		8033 => to_unsigned(22814, LUT_AMPL_WIDTH - 1),
		8034 => to_unsigned(22816, LUT_AMPL_WIDTH - 1),
		8035 => to_unsigned(22818, LUT_AMPL_WIDTH - 1),
		8036 => to_unsigned(22821, LUT_AMPL_WIDTH - 1),
		8037 => to_unsigned(22823, LUT_AMPL_WIDTH - 1),
		8038 => to_unsigned(22825, LUT_AMPL_WIDTH - 1),
		8039 => to_unsigned(22827, LUT_AMPL_WIDTH - 1),
		8040 => to_unsigned(22830, LUT_AMPL_WIDTH - 1),
		8041 => to_unsigned(22832, LUT_AMPL_WIDTH - 1),
		8042 => to_unsigned(22834, LUT_AMPL_WIDTH - 1),
		8043 => to_unsigned(22836, LUT_AMPL_WIDTH - 1),
		8044 => to_unsigned(22839, LUT_AMPL_WIDTH - 1),
		8045 => to_unsigned(22841, LUT_AMPL_WIDTH - 1),
		8046 => to_unsigned(22843, LUT_AMPL_WIDTH - 1),
		8047 => to_unsigned(22845, LUT_AMPL_WIDTH - 1),
		8048 => to_unsigned(22848, LUT_AMPL_WIDTH - 1),
		8049 => to_unsigned(22850, LUT_AMPL_WIDTH - 1),
		8050 => to_unsigned(22852, LUT_AMPL_WIDTH - 1),
		8051 => to_unsigned(22854, LUT_AMPL_WIDTH - 1),
		8052 => to_unsigned(22857, LUT_AMPL_WIDTH - 1),
		8053 => to_unsigned(22859, LUT_AMPL_WIDTH - 1),
		8054 => to_unsigned(22861, LUT_AMPL_WIDTH - 1),
		8055 => to_unsigned(22863, LUT_AMPL_WIDTH - 1),
		8056 => to_unsigned(22866, LUT_AMPL_WIDTH - 1),
		8057 => to_unsigned(22868, LUT_AMPL_WIDTH - 1),
		8058 => to_unsigned(22870, LUT_AMPL_WIDTH - 1),
		8059 => to_unsigned(22872, LUT_AMPL_WIDTH - 1),
		8060 => to_unsigned(22875, LUT_AMPL_WIDTH - 1),
		8061 => to_unsigned(22877, LUT_AMPL_WIDTH - 1),
		8062 => to_unsigned(22879, LUT_AMPL_WIDTH - 1),
		8063 => to_unsigned(22881, LUT_AMPL_WIDTH - 1),
		8064 => to_unsigned(22884, LUT_AMPL_WIDTH - 1),
		8065 => to_unsigned(22886, LUT_AMPL_WIDTH - 1),
		8066 => to_unsigned(22888, LUT_AMPL_WIDTH - 1),
		8067 => to_unsigned(22890, LUT_AMPL_WIDTH - 1),
		8068 => to_unsigned(22893, LUT_AMPL_WIDTH - 1),
		8069 => to_unsigned(22895, LUT_AMPL_WIDTH - 1),
		8070 => to_unsigned(22897, LUT_AMPL_WIDTH - 1),
		8071 => to_unsigned(22899, LUT_AMPL_WIDTH - 1),
		8072 => to_unsigned(22902, LUT_AMPL_WIDTH - 1),
		8073 => to_unsigned(22904, LUT_AMPL_WIDTH - 1),
		8074 => to_unsigned(22906, LUT_AMPL_WIDTH - 1),
		8075 => to_unsigned(22908, LUT_AMPL_WIDTH - 1),
		8076 => to_unsigned(22911, LUT_AMPL_WIDTH - 1),
		8077 => to_unsigned(22913, LUT_AMPL_WIDTH - 1),
		8078 => to_unsigned(22915, LUT_AMPL_WIDTH - 1),
		8079 => to_unsigned(22917, LUT_AMPL_WIDTH - 1),
		8080 => to_unsigned(22920, LUT_AMPL_WIDTH - 1),
		8081 => to_unsigned(22922, LUT_AMPL_WIDTH - 1),
		8082 => to_unsigned(22924, LUT_AMPL_WIDTH - 1),
		8083 => to_unsigned(22926, LUT_AMPL_WIDTH - 1),
		8084 => to_unsigned(22929, LUT_AMPL_WIDTH - 1),
		8085 => to_unsigned(22931, LUT_AMPL_WIDTH - 1),
		8086 => to_unsigned(22933, LUT_AMPL_WIDTH - 1),
		8087 => to_unsigned(22935, LUT_AMPL_WIDTH - 1),
		8088 => to_unsigned(22938, LUT_AMPL_WIDTH - 1),
		8089 => to_unsigned(22940, LUT_AMPL_WIDTH - 1),
		8090 => to_unsigned(22942, LUT_AMPL_WIDTH - 1),
		8091 => to_unsigned(22944, LUT_AMPL_WIDTH - 1),
		8092 => to_unsigned(22947, LUT_AMPL_WIDTH - 1),
		8093 => to_unsigned(22949, LUT_AMPL_WIDTH - 1),
		8094 => to_unsigned(22951, LUT_AMPL_WIDTH - 1),
		8095 => to_unsigned(22953, LUT_AMPL_WIDTH - 1),
		8096 => to_unsigned(22956, LUT_AMPL_WIDTH - 1),
		8097 => to_unsigned(22958, LUT_AMPL_WIDTH - 1),
		8098 => to_unsigned(22960, LUT_AMPL_WIDTH - 1),
		8099 => to_unsigned(22962, LUT_AMPL_WIDTH - 1),
		8100 => to_unsigned(22965, LUT_AMPL_WIDTH - 1),
		8101 => to_unsigned(22967, LUT_AMPL_WIDTH - 1),
		8102 => to_unsigned(22969, LUT_AMPL_WIDTH - 1),
		8103 => to_unsigned(22971, LUT_AMPL_WIDTH - 1),
		8104 => to_unsigned(22973, LUT_AMPL_WIDTH - 1),
		8105 => to_unsigned(22976, LUT_AMPL_WIDTH - 1),
		8106 => to_unsigned(22978, LUT_AMPL_WIDTH - 1),
		8107 => to_unsigned(22980, LUT_AMPL_WIDTH - 1),
		8108 => to_unsigned(22982, LUT_AMPL_WIDTH - 1),
		8109 => to_unsigned(22985, LUT_AMPL_WIDTH - 1),
		8110 => to_unsigned(22987, LUT_AMPL_WIDTH - 1),
		8111 => to_unsigned(22989, LUT_AMPL_WIDTH - 1),
		8112 => to_unsigned(22991, LUT_AMPL_WIDTH - 1),
		8113 => to_unsigned(22994, LUT_AMPL_WIDTH - 1),
		8114 => to_unsigned(22996, LUT_AMPL_WIDTH - 1),
		8115 => to_unsigned(22998, LUT_AMPL_WIDTH - 1),
		8116 => to_unsigned(23000, LUT_AMPL_WIDTH - 1),
		8117 => to_unsigned(23003, LUT_AMPL_WIDTH - 1),
		8118 => to_unsigned(23005, LUT_AMPL_WIDTH - 1),
		8119 => to_unsigned(23007, LUT_AMPL_WIDTH - 1),
		8120 => to_unsigned(23009, LUT_AMPL_WIDTH - 1),
		8121 => to_unsigned(23012, LUT_AMPL_WIDTH - 1),
		8122 => to_unsigned(23014, LUT_AMPL_WIDTH - 1),
		8123 => to_unsigned(23016, LUT_AMPL_WIDTH - 1),
		8124 => to_unsigned(23018, LUT_AMPL_WIDTH - 1),
		8125 => to_unsigned(23020, LUT_AMPL_WIDTH - 1),
		8126 => to_unsigned(23023, LUT_AMPL_WIDTH - 1),
		8127 => to_unsigned(23025, LUT_AMPL_WIDTH - 1),
		8128 => to_unsigned(23027, LUT_AMPL_WIDTH - 1),
		8129 => to_unsigned(23029, LUT_AMPL_WIDTH - 1),
		8130 => to_unsigned(23032, LUT_AMPL_WIDTH - 1),
		8131 => to_unsigned(23034, LUT_AMPL_WIDTH - 1),
		8132 => to_unsigned(23036, LUT_AMPL_WIDTH - 1),
		8133 => to_unsigned(23038, LUT_AMPL_WIDTH - 1),
		8134 => to_unsigned(23041, LUT_AMPL_WIDTH - 1),
		8135 => to_unsigned(23043, LUT_AMPL_WIDTH - 1),
		8136 => to_unsigned(23045, LUT_AMPL_WIDTH - 1),
		8137 => to_unsigned(23047, LUT_AMPL_WIDTH - 1),
		8138 => to_unsigned(23050, LUT_AMPL_WIDTH - 1),
		8139 => to_unsigned(23052, LUT_AMPL_WIDTH - 1),
		8140 => to_unsigned(23054, LUT_AMPL_WIDTH - 1),
		8141 => to_unsigned(23056, LUT_AMPL_WIDTH - 1),
		8142 => to_unsigned(23058, LUT_AMPL_WIDTH - 1),
		8143 => to_unsigned(23061, LUT_AMPL_WIDTH - 1),
		8144 => to_unsigned(23063, LUT_AMPL_WIDTH - 1),
		8145 => to_unsigned(23065, LUT_AMPL_WIDTH - 1),
		8146 => to_unsigned(23067, LUT_AMPL_WIDTH - 1),
		8147 => to_unsigned(23070, LUT_AMPL_WIDTH - 1),
		8148 => to_unsigned(23072, LUT_AMPL_WIDTH - 1),
		8149 => to_unsigned(23074, LUT_AMPL_WIDTH - 1),
		8150 => to_unsigned(23076, LUT_AMPL_WIDTH - 1),
		8151 => to_unsigned(23079, LUT_AMPL_WIDTH - 1),
		8152 => to_unsigned(23081, LUT_AMPL_WIDTH - 1),
		8153 => to_unsigned(23083, LUT_AMPL_WIDTH - 1),
		8154 => to_unsigned(23085, LUT_AMPL_WIDTH - 1),
		8155 => to_unsigned(23087, LUT_AMPL_WIDTH - 1),
		8156 => to_unsigned(23090, LUT_AMPL_WIDTH - 1),
		8157 => to_unsigned(23092, LUT_AMPL_WIDTH - 1),
		8158 => to_unsigned(23094, LUT_AMPL_WIDTH - 1),
		8159 => to_unsigned(23096, LUT_AMPL_WIDTH - 1),
		8160 => to_unsigned(23099, LUT_AMPL_WIDTH - 1),
		8161 => to_unsigned(23101, LUT_AMPL_WIDTH - 1),
		8162 => to_unsigned(23103, LUT_AMPL_WIDTH - 1),
		8163 => to_unsigned(23105, LUT_AMPL_WIDTH - 1),
		8164 => to_unsigned(23107, LUT_AMPL_WIDTH - 1),
		8165 => to_unsigned(23110, LUT_AMPL_WIDTH - 1),
		8166 => to_unsigned(23112, LUT_AMPL_WIDTH - 1),
		8167 => to_unsigned(23114, LUT_AMPL_WIDTH - 1),
		8168 => to_unsigned(23116, LUT_AMPL_WIDTH - 1),
		8169 => to_unsigned(23119, LUT_AMPL_WIDTH - 1),
		8170 => to_unsigned(23121, LUT_AMPL_WIDTH - 1),
		8171 => to_unsigned(23123, LUT_AMPL_WIDTH - 1),
		8172 => to_unsigned(23125, LUT_AMPL_WIDTH - 1),
		8173 => to_unsigned(23128, LUT_AMPL_WIDTH - 1),
		8174 => to_unsigned(23130, LUT_AMPL_WIDTH - 1),
		8175 => to_unsigned(23132, LUT_AMPL_WIDTH - 1),
		8176 => to_unsigned(23134, LUT_AMPL_WIDTH - 1),
		8177 => to_unsigned(23136, LUT_AMPL_WIDTH - 1),
		8178 => to_unsigned(23139, LUT_AMPL_WIDTH - 1),
		8179 => to_unsigned(23141, LUT_AMPL_WIDTH - 1),
		8180 => to_unsigned(23143, LUT_AMPL_WIDTH - 1),
		8181 => to_unsigned(23145, LUT_AMPL_WIDTH - 1),
		8182 => to_unsigned(23148, LUT_AMPL_WIDTH - 1),
		8183 => to_unsigned(23150, LUT_AMPL_WIDTH - 1),
		8184 => to_unsigned(23152, LUT_AMPL_WIDTH - 1),
		8185 => to_unsigned(23154, LUT_AMPL_WIDTH - 1),
		8186 => to_unsigned(23156, LUT_AMPL_WIDTH - 1),
		8187 => to_unsigned(23159, LUT_AMPL_WIDTH - 1),
		8188 => to_unsigned(23161, LUT_AMPL_WIDTH - 1),
		8189 => to_unsigned(23163, LUT_AMPL_WIDTH - 1),
		8190 => to_unsigned(23165, LUT_AMPL_WIDTH - 1),
		8191 => to_unsigned(23168, LUT_AMPL_WIDTH - 1),
		8192 => to_unsigned(23170, LUT_AMPL_WIDTH - 1),
		8193 => to_unsigned(23172, LUT_AMPL_WIDTH - 1),
		8194 => to_unsigned(23174, LUT_AMPL_WIDTH - 1),
		8195 => to_unsigned(23176, LUT_AMPL_WIDTH - 1),
		8196 => to_unsigned(23179, LUT_AMPL_WIDTH - 1),
		8197 => to_unsigned(23181, LUT_AMPL_WIDTH - 1),
		8198 => to_unsigned(23183, LUT_AMPL_WIDTH - 1),
		8199 => to_unsigned(23185, LUT_AMPL_WIDTH - 1),
		8200 => to_unsigned(23188, LUT_AMPL_WIDTH - 1),
		8201 => to_unsigned(23190, LUT_AMPL_WIDTH - 1),
		8202 => to_unsigned(23192, LUT_AMPL_WIDTH - 1),
		8203 => to_unsigned(23194, LUT_AMPL_WIDTH - 1),
		8204 => to_unsigned(23196, LUT_AMPL_WIDTH - 1),
		8205 => to_unsigned(23199, LUT_AMPL_WIDTH - 1),
		8206 => to_unsigned(23201, LUT_AMPL_WIDTH - 1),
		8207 => to_unsigned(23203, LUT_AMPL_WIDTH - 1),
		8208 => to_unsigned(23205, LUT_AMPL_WIDTH - 1),
		8209 => to_unsigned(23208, LUT_AMPL_WIDTH - 1),
		8210 => to_unsigned(23210, LUT_AMPL_WIDTH - 1),
		8211 => to_unsigned(23212, LUT_AMPL_WIDTH - 1),
		8212 => to_unsigned(23214, LUT_AMPL_WIDTH - 1),
		8213 => to_unsigned(23216, LUT_AMPL_WIDTH - 1),
		8214 => to_unsigned(23219, LUT_AMPL_WIDTH - 1),
		8215 => to_unsigned(23221, LUT_AMPL_WIDTH - 1),
		8216 => to_unsigned(23223, LUT_AMPL_WIDTH - 1),
		8217 => to_unsigned(23225, LUT_AMPL_WIDTH - 1),
		8218 => to_unsigned(23227, LUT_AMPL_WIDTH - 1),
		8219 => to_unsigned(23230, LUT_AMPL_WIDTH - 1),
		8220 => to_unsigned(23232, LUT_AMPL_WIDTH - 1),
		8221 => to_unsigned(23234, LUT_AMPL_WIDTH - 1),
		8222 => to_unsigned(23236, LUT_AMPL_WIDTH - 1),
		8223 => to_unsigned(23239, LUT_AMPL_WIDTH - 1),
		8224 => to_unsigned(23241, LUT_AMPL_WIDTH - 1),
		8225 => to_unsigned(23243, LUT_AMPL_WIDTH - 1),
		8226 => to_unsigned(23245, LUT_AMPL_WIDTH - 1),
		8227 => to_unsigned(23247, LUT_AMPL_WIDTH - 1),
		8228 => to_unsigned(23250, LUT_AMPL_WIDTH - 1),
		8229 => to_unsigned(23252, LUT_AMPL_WIDTH - 1),
		8230 => to_unsigned(23254, LUT_AMPL_WIDTH - 1),
		8231 => to_unsigned(23256, LUT_AMPL_WIDTH - 1),
		8232 => to_unsigned(23258, LUT_AMPL_WIDTH - 1),
		8233 => to_unsigned(23261, LUT_AMPL_WIDTH - 1),
		8234 => to_unsigned(23263, LUT_AMPL_WIDTH - 1),
		8235 => to_unsigned(23265, LUT_AMPL_WIDTH - 1),
		8236 => to_unsigned(23267, LUT_AMPL_WIDTH - 1),
		8237 => to_unsigned(23270, LUT_AMPL_WIDTH - 1),
		8238 => to_unsigned(23272, LUT_AMPL_WIDTH - 1),
		8239 => to_unsigned(23274, LUT_AMPL_WIDTH - 1),
		8240 => to_unsigned(23276, LUT_AMPL_WIDTH - 1),
		8241 => to_unsigned(23278, LUT_AMPL_WIDTH - 1),
		8242 => to_unsigned(23281, LUT_AMPL_WIDTH - 1),
		8243 => to_unsigned(23283, LUT_AMPL_WIDTH - 1),
		8244 => to_unsigned(23285, LUT_AMPL_WIDTH - 1),
		8245 => to_unsigned(23287, LUT_AMPL_WIDTH - 1),
		8246 => to_unsigned(23289, LUT_AMPL_WIDTH - 1),
		8247 => to_unsigned(23292, LUT_AMPL_WIDTH - 1),
		8248 => to_unsigned(23294, LUT_AMPL_WIDTH - 1),
		8249 => to_unsigned(23296, LUT_AMPL_WIDTH - 1),
		8250 => to_unsigned(23298, LUT_AMPL_WIDTH - 1),
		8251 => to_unsigned(23300, LUT_AMPL_WIDTH - 1),
		8252 => to_unsigned(23303, LUT_AMPL_WIDTH - 1),
		8253 => to_unsigned(23305, LUT_AMPL_WIDTH - 1),
		8254 => to_unsigned(23307, LUT_AMPL_WIDTH - 1),
		8255 => to_unsigned(23309, LUT_AMPL_WIDTH - 1),
		8256 => to_unsigned(23311, LUT_AMPL_WIDTH - 1),
		8257 => to_unsigned(23314, LUT_AMPL_WIDTH - 1),
		8258 => to_unsigned(23316, LUT_AMPL_WIDTH - 1),
		8259 => to_unsigned(23318, LUT_AMPL_WIDTH - 1),
		8260 => to_unsigned(23320, LUT_AMPL_WIDTH - 1),
		8261 => to_unsigned(23323, LUT_AMPL_WIDTH - 1),
		8262 => to_unsigned(23325, LUT_AMPL_WIDTH - 1),
		8263 => to_unsigned(23327, LUT_AMPL_WIDTH - 1),
		8264 => to_unsigned(23329, LUT_AMPL_WIDTH - 1),
		8265 => to_unsigned(23331, LUT_AMPL_WIDTH - 1),
		8266 => to_unsigned(23334, LUT_AMPL_WIDTH - 1),
		8267 => to_unsigned(23336, LUT_AMPL_WIDTH - 1),
		8268 => to_unsigned(23338, LUT_AMPL_WIDTH - 1),
		8269 => to_unsigned(23340, LUT_AMPL_WIDTH - 1),
		8270 => to_unsigned(23342, LUT_AMPL_WIDTH - 1),
		8271 => to_unsigned(23345, LUT_AMPL_WIDTH - 1),
		8272 => to_unsigned(23347, LUT_AMPL_WIDTH - 1),
		8273 => to_unsigned(23349, LUT_AMPL_WIDTH - 1),
		8274 => to_unsigned(23351, LUT_AMPL_WIDTH - 1),
		8275 => to_unsigned(23353, LUT_AMPL_WIDTH - 1),
		8276 => to_unsigned(23356, LUT_AMPL_WIDTH - 1),
		8277 => to_unsigned(23358, LUT_AMPL_WIDTH - 1),
		8278 => to_unsigned(23360, LUT_AMPL_WIDTH - 1),
		8279 => to_unsigned(23362, LUT_AMPL_WIDTH - 1),
		8280 => to_unsigned(23364, LUT_AMPL_WIDTH - 1),
		8281 => to_unsigned(23367, LUT_AMPL_WIDTH - 1),
		8282 => to_unsigned(23369, LUT_AMPL_WIDTH - 1),
		8283 => to_unsigned(23371, LUT_AMPL_WIDTH - 1),
		8284 => to_unsigned(23373, LUT_AMPL_WIDTH - 1),
		8285 => to_unsigned(23375, LUT_AMPL_WIDTH - 1),
		8286 => to_unsigned(23378, LUT_AMPL_WIDTH - 1),
		8287 => to_unsigned(23380, LUT_AMPL_WIDTH - 1),
		8288 => to_unsigned(23382, LUT_AMPL_WIDTH - 1),
		8289 => to_unsigned(23384, LUT_AMPL_WIDTH - 1),
		8290 => to_unsigned(23386, LUT_AMPL_WIDTH - 1),
		8291 => to_unsigned(23389, LUT_AMPL_WIDTH - 1),
		8292 => to_unsigned(23391, LUT_AMPL_WIDTH - 1),
		8293 => to_unsigned(23393, LUT_AMPL_WIDTH - 1),
		8294 => to_unsigned(23395, LUT_AMPL_WIDTH - 1),
		8295 => to_unsigned(23397, LUT_AMPL_WIDTH - 1),
		8296 => to_unsigned(23400, LUT_AMPL_WIDTH - 1),
		8297 => to_unsigned(23402, LUT_AMPL_WIDTH - 1),
		8298 => to_unsigned(23404, LUT_AMPL_WIDTH - 1),
		8299 => to_unsigned(23406, LUT_AMPL_WIDTH - 1),
		8300 => to_unsigned(23408, LUT_AMPL_WIDTH - 1),
		8301 => to_unsigned(23411, LUT_AMPL_WIDTH - 1),
		8302 => to_unsigned(23413, LUT_AMPL_WIDTH - 1),
		8303 => to_unsigned(23415, LUT_AMPL_WIDTH - 1),
		8304 => to_unsigned(23417, LUT_AMPL_WIDTH - 1),
		8305 => to_unsigned(23419, LUT_AMPL_WIDTH - 1),
		8306 => to_unsigned(23422, LUT_AMPL_WIDTH - 1),
		8307 => to_unsigned(23424, LUT_AMPL_WIDTH - 1),
		8308 => to_unsigned(23426, LUT_AMPL_WIDTH - 1),
		8309 => to_unsigned(23428, LUT_AMPL_WIDTH - 1),
		8310 => to_unsigned(23430, LUT_AMPL_WIDTH - 1),
		8311 => to_unsigned(23433, LUT_AMPL_WIDTH - 1),
		8312 => to_unsigned(23435, LUT_AMPL_WIDTH - 1),
		8313 => to_unsigned(23437, LUT_AMPL_WIDTH - 1),
		8314 => to_unsigned(23439, LUT_AMPL_WIDTH - 1),
		8315 => to_unsigned(23441, LUT_AMPL_WIDTH - 1),
		8316 => to_unsigned(23444, LUT_AMPL_WIDTH - 1),
		8317 => to_unsigned(23446, LUT_AMPL_WIDTH - 1),
		8318 => to_unsigned(23448, LUT_AMPL_WIDTH - 1),
		8319 => to_unsigned(23450, LUT_AMPL_WIDTH - 1),
		8320 => to_unsigned(23452, LUT_AMPL_WIDTH - 1),
		8321 => to_unsigned(23455, LUT_AMPL_WIDTH - 1),
		8322 => to_unsigned(23457, LUT_AMPL_WIDTH - 1),
		8323 => to_unsigned(23459, LUT_AMPL_WIDTH - 1),
		8324 => to_unsigned(23461, LUT_AMPL_WIDTH - 1),
		8325 => to_unsigned(23463, LUT_AMPL_WIDTH - 1),
		8326 => to_unsigned(23466, LUT_AMPL_WIDTH - 1),
		8327 => to_unsigned(23468, LUT_AMPL_WIDTH - 1),
		8328 => to_unsigned(23470, LUT_AMPL_WIDTH - 1),
		8329 => to_unsigned(23472, LUT_AMPL_WIDTH - 1),
		8330 => to_unsigned(23474, LUT_AMPL_WIDTH - 1),
		8331 => to_unsigned(23476, LUT_AMPL_WIDTH - 1),
		8332 => to_unsigned(23479, LUT_AMPL_WIDTH - 1),
		8333 => to_unsigned(23481, LUT_AMPL_WIDTH - 1),
		8334 => to_unsigned(23483, LUT_AMPL_WIDTH - 1),
		8335 => to_unsigned(23485, LUT_AMPL_WIDTH - 1),
		8336 => to_unsigned(23487, LUT_AMPL_WIDTH - 1),
		8337 => to_unsigned(23490, LUT_AMPL_WIDTH - 1),
		8338 => to_unsigned(23492, LUT_AMPL_WIDTH - 1),
		8339 => to_unsigned(23494, LUT_AMPL_WIDTH - 1),
		8340 => to_unsigned(23496, LUT_AMPL_WIDTH - 1),
		8341 => to_unsigned(23498, LUT_AMPL_WIDTH - 1),
		8342 => to_unsigned(23501, LUT_AMPL_WIDTH - 1),
		8343 => to_unsigned(23503, LUT_AMPL_WIDTH - 1),
		8344 => to_unsigned(23505, LUT_AMPL_WIDTH - 1),
		8345 => to_unsigned(23507, LUT_AMPL_WIDTH - 1),
		8346 => to_unsigned(23509, LUT_AMPL_WIDTH - 1),
		8347 => to_unsigned(23512, LUT_AMPL_WIDTH - 1),
		8348 => to_unsigned(23514, LUT_AMPL_WIDTH - 1),
		8349 => to_unsigned(23516, LUT_AMPL_WIDTH - 1),
		8350 => to_unsigned(23518, LUT_AMPL_WIDTH - 1),
		8351 => to_unsigned(23520, LUT_AMPL_WIDTH - 1),
		8352 => to_unsigned(23522, LUT_AMPL_WIDTH - 1),
		8353 => to_unsigned(23525, LUT_AMPL_WIDTH - 1),
		8354 => to_unsigned(23527, LUT_AMPL_WIDTH - 1),
		8355 => to_unsigned(23529, LUT_AMPL_WIDTH - 1),
		8356 => to_unsigned(23531, LUT_AMPL_WIDTH - 1),
		8357 => to_unsigned(23533, LUT_AMPL_WIDTH - 1),
		8358 => to_unsigned(23536, LUT_AMPL_WIDTH - 1),
		8359 => to_unsigned(23538, LUT_AMPL_WIDTH - 1),
		8360 => to_unsigned(23540, LUT_AMPL_WIDTH - 1),
		8361 => to_unsigned(23542, LUT_AMPL_WIDTH - 1),
		8362 => to_unsigned(23544, LUT_AMPL_WIDTH - 1),
		8363 => to_unsigned(23546, LUT_AMPL_WIDTH - 1),
		8364 => to_unsigned(23549, LUT_AMPL_WIDTH - 1),
		8365 => to_unsigned(23551, LUT_AMPL_WIDTH - 1),
		8366 => to_unsigned(23553, LUT_AMPL_WIDTH - 1),
		8367 => to_unsigned(23555, LUT_AMPL_WIDTH - 1),
		8368 => to_unsigned(23557, LUT_AMPL_WIDTH - 1),
		8369 => to_unsigned(23560, LUT_AMPL_WIDTH - 1),
		8370 => to_unsigned(23562, LUT_AMPL_WIDTH - 1),
		8371 => to_unsigned(23564, LUT_AMPL_WIDTH - 1),
		8372 => to_unsigned(23566, LUT_AMPL_WIDTH - 1),
		8373 => to_unsigned(23568, LUT_AMPL_WIDTH - 1),
		8374 => to_unsigned(23571, LUT_AMPL_WIDTH - 1),
		8375 => to_unsigned(23573, LUT_AMPL_WIDTH - 1),
		8376 => to_unsigned(23575, LUT_AMPL_WIDTH - 1),
		8377 => to_unsigned(23577, LUT_AMPL_WIDTH - 1),
		8378 => to_unsigned(23579, LUT_AMPL_WIDTH - 1),
		8379 => to_unsigned(23581, LUT_AMPL_WIDTH - 1),
		8380 => to_unsigned(23584, LUT_AMPL_WIDTH - 1),
		8381 => to_unsigned(23586, LUT_AMPL_WIDTH - 1),
		8382 => to_unsigned(23588, LUT_AMPL_WIDTH - 1),
		8383 => to_unsigned(23590, LUT_AMPL_WIDTH - 1),
		8384 => to_unsigned(23592, LUT_AMPL_WIDTH - 1),
		8385 => to_unsigned(23595, LUT_AMPL_WIDTH - 1),
		8386 => to_unsigned(23597, LUT_AMPL_WIDTH - 1),
		8387 => to_unsigned(23599, LUT_AMPL_WIDTH - 1),
		8388 => to_unsigned(23601, LUT_AMPL_WIDTH - 1),
		8389 => to_unsigned(23603, LUT_AMPL_WIDTH - 1),
		8390 => to_unsigned(23605, LUT_AMPL_WIDTH - 1),
		8391 => to_unsigned(23608, LUT_AMPL_WIDTH - 1),
		8392 => to_unsigned(23610, LUT_AMPL_WIDTH - 1),
		8393 => to_unsigned(23612, LUT_AMPL_WIDTH - 1),
		8394 => to_unsigned(23614, LUT_AMPL_WIDTH - 1),
		8395 => to_unsigned(23616, LUT_AMPL_WIDTH - 1),
		8396 => to_unsigned(23618, LUT_AMPL_WIDTH - 1),
		8397 => to_unsigned(23621, LUT_AMPL_WIDTH - 1),
		8398 => to_unsigned(23623, LUT_AMPL_WIDTH - 1),
		8399 => to_unsigned(23625, LUT_AMPL_WIDTH - 1),
		8400 => to_unsigned(23627, LUT_AMPL_WIDTH - 1),
		8401 => to_unsigned(23629, LUT_AMPL_WIDTH - 1),
		8402 => to_unsigned(23632, LUT_AMPL_WIDTH - 1),
		8403 => to_unsigned(23634, LUT_AMPL_WIDTH - 1),
		8404 => to_unsigned(23636, LUT_AMPL_WIDTH - 1),
		8405 => to_unsigned(23638, LUT_AMPL_WIDTH - 1),
		8406 => to_unsigned(23640, LUT_AMPL_WIDTH - 1),
		8407 => to_unsigned(23642, LUT_AMPL_WIDTH - 1),
		8408 => to_unsigned(23645, LUT_AMPL_WIDTH - 1),
		8409 => to_unsigned(23647, LUT_AMPL_WIDTH - 1),
		8410 => to_unsigned(23649, LUT_AMPL_WIDTH - 1),
		8411 => to_unsigned(23651, LUT_AMPL_WIDTH - 1),
		8412 => to_unsigned(23653, LUT_AMPL_WIDTH - 1),
		8413 => to_unsigned(23655, LUT_AMPL_WIDTH - 1),
		8414 => to_unsigned(23658, LUT_AMPL_WIDTH - 1),
		8415 => to_unsigned(23660, LUT_AMPL_WIDTH - 1),
		8416 => to_unsigned(23662, LUT_AMPL_WIDTH - 1),
		8417 => to_unsigned(23664, LUT_AMPL_WIDTH - 1),
		8418 => to_unsigned(23666, LUT_AMPL_WIDTH - 1),
		8419 => to_unsigned(23668, LUT_AMPL_WIDTH - 1),
		8420 => to_unsigned(23671, LUT_AMPL_WIDTH - 1),
		8421 => to_unsigned(23673, LUT_AMPL_WIDTH - 1),
		8422 => to_unsigned(23675, LUT_AMPL_WIDTH - 1),
		8423 => to_unsigned(23677, LUT_AMPL_WIDTH - 1),
		8424 => to_unsigned(23679, LUT_AMPL_WIDTH - 1),
		8425 => to_unsigned(23682, LUT_AMPL_WIDTH - 1),
		8426 => to_unsigned(23684, LUT_AMPL_WIDTH - 1),
		8427 => to_unsigned(23686, LUT_AMPL_WIDTH - 1),
		8428 => to_unsigned(23688, LUT_AMPL_WIDTH - 1),
		8429 => to_unsigned(23690, LUT_AMPL_WIDTH - 1),
		8430 => to_unsigned(23692, LUT_AMPL_WIDTH - 1),
		8431 => to_unsigned(23695, LUT_AMPL_WIDTH - 1),
		8432 => to_unsigned(23697, LUT_AMPL_WIDTH - 1),
		8433 => to_unsigned(23699, LUT_AMPL_WIDTH - 1),
		8434 => to_unsigned(23701, LUT_AMPL_WIDTH - 1),
		8435 => to_unsigned(23703, LUT_AMPL_WIDTH - 1),
		8436 => to_unsigned(23705, LUT_AMPL_WIDTH - 1),
		8437 => to_unsigned(23708, LUT_AMPL_WIDTH - 1),
		8438 => to_unsigned(23710, LUT_AMPL_WIDTH - 1),
		8439 => to_unsigned(23712, LUT_AMPL_WIDTH - 1),
		8440 => to_unsigned(23714, LUT_AMPL_WIDTH - 1),
		8441 => to_unsigned(23716, LUT_AMPL_WIDTH - 1),
		8442 => to_unsigned(23718, LUT_AMPL_WIDTH - 1),
		8443 => to_unsigned(23721, LUT_AMPL_WIDTH - 1),
		8444 => to_unsigned(23723, LUT_AMPL_WIDTH - 1),
		8445 => to_unsigned(23725, LUT_AMPL_WIDTH - 1),
		8446 => to_unsigned(23727, LUT_AMPL_WIDTH - 1),
		8447 => to_unsigned(23729, LUT_AMPL_WIDTH - 1),
		8448 => to_unsigned(23731, LUT_AMPL_WIDTH - 1),
		8449 => to_unsigned(23734, LUT_AMPL_WIDTH - 1),
		8450 => to_unsigned(23736, LUT_AMPL_WIDTH - 1),
		8451 => to_unsigned(23738, LUT_AMPL_WIDTH - 1),
		8452 => to_unsigned(23740, LUT_AMPL_WIDTH - 1),
		8453 => to_unsigned(23742, LUT_AMPL_WIDTH - 1),
		8454 => to_unsigned(23744, LUT_AMPL_WIDTH - 1),
		8455 => to_unsigned(23747, LUT_AMPL_WIDTH - 1),
		8456 => to_unsigned(23749, LUT_AMPL_WIDTH - 1),
		8457 => to_unsigned(23751, LUT_AMPL_WIDTH - 1),
		8458 => to_unsigned(23753, LUT_AMPL_WIDTH - 1),
		8459 => to_unsigned(23755, LUT_AMPL_WIDTH - 1),
		8460 => to_unsigned(23757, LUT_AMPL_WIDTH - 1),
		8461 => to_unsigned(23760, LUT_AMPL_WIDTH - 1),
		8462 => to_unsigned(23762, LUT_AMPL_WIDTH - 1),
		8463 => to_unsigned(23764, LUT_AMPL_WIDTH - 1),
		8464 => to_unsigned(23766, LUT_AMPL_WIDTH - 1),
		8465 => to_unsigned(23768, LUT_AMPL_WIDTH - 1),
		8466 => to_unsigned(23770, LUT_AMPL_WIDTH - 1),
		8467 => to_unsigned(23773, LUT_AMPL_WIDTH - 1),
		8468 => to_unsigned(23775, LUT_AMPL_WIDTH - 1),
		8469 => to_unsigned(23777, LUT_AMPL_WIDTH - 1),
		8470 => to_unsigned(23779, LUT_AMPL_WIDTH - 1),
		8471 => to_unsigned(23781, LUT_AMPL_WIDTH - 1),
		8472 => to_unsigned(23783, LUT_AMPL_WIDTH - 1),
		8473 => to_unsigned(23785, LUT_AMPL_WIDTH - 1),
		8474 => to_unsigned(23788, LUT_AMPL_WIDTH - 1),
		8475 => to_unsigned(23790, LUT_AMPL_WIDTH - 1),
		8476 => to_unsigned(23792, LUT_AMPL_WIDTH - 1),
		8477 => to_unsigned(23794, LUT_AMPL_WIDTH - 1),
		8478 => to_unsigned(23796, LUT_AMPL_WIDTH - 1),
		8479 => to_unsigned(23798, LUT_AMPL_WIDTH - 1),
		8480 => to_unsigned(23801, LUT_AMPL_WIDTH - 1),
		8481 => to_unsigned(23803, LUT_AMPL_WIDTH - 1),
		8482 => to_unsigned(23805, LUT_AMPL_WIDTH - 1),
		8483 => to_unsigned(23807, LUT_AMPL_WIDTH - 1),
		8484 => to_unsigned(23809, LUT_AMPL_WIDTH - 1),
		8485 => to_unsigned(23811, LUT_AMPL_WIDTH - 1),
		8486 => to_unsigned(23814, LUT_AMPL_WIDTH - 1),
		8487 => to_unsigned(23816, LUT_AMPL_WIDTH - 1),
		8488 => to_unsigned(23818, LUT_AMPL_WIDTH - 1),
		8489 => to_unsigned(23820, LUT_AMPL_WIDTH - 1),
		8490 => to_unsigned(23822, LUT_AMPL_WIDTH - 1),
		8491 => to_unsigned(23824, LUT_AMPL_WIDTH - 1),
		8492 => to_unsigned(23827, LUT_AMPL_WIDTH - 1),
		8493 => to_unsigned(23829, LUT_AMPL_WIDTH - 1),
		8494 => to_unsigned(23831, LUT_AMPL_WIDTH - 1),
		8495 => to_unsigned(23833, LUT_AMPL_WIDTH - 1),
		8496 => to_unsigned(23835, LUT_AMPL_WIDTH - 1),
		8497 => to_unsigned(23837, LUT_AMPL_WIDTH - 1),
		8498 => to_unsigned(23839, LUT_AMPL_WIDTH - 1),
		8499 => to_unsigned(23842, LUT_AMPL_WIDTH - 1),
		8500 => to_unsigned(23844, LUT_AMPL_WIDTH - 1),
		8501 => to_unsigned(23846, LUT_AMPL_WIDTH - 1),
		8502 => to_unsigned(23848, LUT_AMPL_WIDTH - 1),
		8503 => to_unsigned(23850, LUT_AMPL_WIDTH - 1),
		8504 => to_unsigned(23852, LUT_AMPL_WIDTH - 1),
		8505 => to_unsigned(23855, LUT_AMPL_WIDTH - 1),
		8506 => to_unsigned(23857, LUT_AMPL_WIDTH - 1),
		8507 => to_unsigned(23859, LUT_AMPL_WIDTH - 1),
		8508 => to_unsigned(23861, LUT_AMPL_WIDTH - 1),
		8509 => to_unsigned(23863, LUT_AMPL_WIDTH - 1),
		8510 => to_unsigned(23865, LUT_AMPL_WIDTH - 1),
		8511 => to_unsigned(23867, LUT_AMPL_WIDTH - 1),
		8512 => to_unsigned(23870, LUT_AMPL_WIDTH - 1),
		8513 => to_unsigned(23872, LUT_AMPL_WIDTH - 1),
		8514 => to_unsigned(23874, LUT_AMPL_WIDTH - 1),
		8515 => to_unsigned(23876, LUT_AMPL_WIDTH - 1),
		8516 => to_unsigned(23878, LUT_AMPL_WIDTH - 1),
		8517 => to_unsigned(23880, LUT_AMPL_WIDTH - 1),
		8518 => to_unsigned(23883, LUT_AMPL_WIDTH - 1),
		8519 => to_unsigned(23885, LUT_AMPL_WIDTH - 1),
		8520 => to_unsigned(23887, LUT_AMPL_WIDTH - 1),
		8521 => to_unsigned(23889, LUT_AMPL_WIDTH - 1),
		8522 => to_unsigned(23891, LUT_AMPL_WIDTH - 1),
		8523 => to_unsigned(23893, LUT_AMPL_WIDTH - 1),
		8524 => to_unsigned(23895, LUT_AMPL_WIDTH - 1),
		8525 => to_unsigned(23898, LUT_AMPL_WIDTH - 1),
		8526 => to_unsigned(23900, LUT_AMPL_WIDTH - 1),
		8527 => to_unsigned(23902, LUT_AMPL_WIDTH - 1),
		8528 => to_unsigned(23904, LUT_AMPL_WIDTH - 1),
		8529 => to_unsigned(23906, LUT_AMPL_WIDTH - 1),
		8530 => to_unsigned(23908, LUT_AMPL_WIDTH - 1),
		8531 => to_unsigned(23910, LUT_AMPL_WIDTH - 1),
		8532 => to_unsigned(23913, LUT_AMPL_WIDTH - 1),
		8533 => to_unsigned(23915, LUT_AMPL_WIDTH - 1),
		8534 => to_unsigned(23917, LUT_AMPL_WIDTH - 1),
		8535 => to_unsigned(23919, LUT_AMPL_WIDTH - 1),
		8536 => to_unsigned(23921, LUT_AMPL_WIDTH - 1),
		8537 => to_unsigned(23923, LUT_AMPL_WIDTH - 1),
		8538 => to_unsigned(23925, LUT_AMPL_WIDTH - 1),
		8539 => to_unsigned(23928, LUT_AMPL_WIDTH - 1),
		8540 => to_unsigned(23930, LUT_AMPL_WIDTH - 1),
		8541 => to_unsigned(23932, LUT_AMPL_WIDTH - 1),
		8542 => to_unsigned(23934, LUT_AMPL_WIDTH - 1),
		8543 => to_unsigned(23936, LUT_AMPL_WIDTH - 1),
		8544 => to_unsigned(23938, LUT_AMPL_WIDTH - 1),
		8545 => to_unsigned(23940, LUT_AMPL_WIDTH - 1),
		8546 => to_unsigned(23943, LUT_AMPL_WIDTH - 1),
		8547 => to_unsigned(23945, LUT_AMPL_WIDTH - 1),
		8548 => to_unsigned(23947, LUT_AMPL_WIDTH - 1),
		8549 => to_unsigned(23949, LUT_AMPL_WIDTH - 1),
		8550 => to_unsigned(23951, LUT_AMPL_WIDTH - 1),
		8551 => to_unsigned(23953, LUT_AMPL_WIDTH - 1),
		8552 => to_unsigned(23956, LUT_AMPL_WIDTH - 1),
		8553 => to_unsigned(23958, LUT_AMPL_WIDTH - 1),
		8554 => to_unsigned(23960, LUT_AMPL_WIDTH - 1),
		8555 => to_unsigned(23962, LUT_AMPL_WIDTH - 1),
		8556 => to_unsigned(23964, LUT_AMPL_WIDTH - 1),
		8557 => to_unsigned(23966, LUT_AMPL_WIDTH - 1),
		8558 => to_unsigned(23968, LUT_AMPL_WIDTH - 1),
		8559 => to_unsigned(23971, LUT_AMPL_WIDTH - 1),
		8560 => to_unsigned(23973, LUT_AMPL_WIDTH - 1),
		8561 => to_unsigned(23975, LUT_AMPL_WIDTH - 1),
		8562 => to_unsigned(23977, LUT_AMPL_WIDTH - 1),
		8563 => to_unsigned(23979, LUT_AMPL_WIDTH - 1),
		8564 => to_unsigned(23981, LUT_AMPL_WIDTH - 1),
		8565 => to_unsigned(23983, LUT_AMPL_WIDTH - 1),
		8566 => to_unsigned(23985, LUT_AMPL_WIDTH - 1),
		8567 => to_unsigned(23988, LUT_AMPL_WIDTH - 1),
		8568 => to_unsigned(23990, LUT_AMPL_WIDTH - 1),
		8569 => to_unsigned(23992, LUT_AMPL_WIDTH - 1),
		8570 => to_unsigned(23994, LUT_AMPL_WIDTH - 1),
		8571 => to_unsigned(23996, LUT_AMPL_WIDTH - 1),
		8572 => to_unsigned(23998, LUT_AMPL_WIDTH - 1),
		8573 => to_unsigned(24000, LUT_AMPL_WIDTH - 1),
		8574 => to_unsigned(24003, LUT_AMPL_WIDTH - 1),
		8575 => to_unsigned(24005, LUT_AMPL_WIDTH - 1),
		8576 => to_unsigned(24007, LUT_AMPL_WIDTH - 1),
		8577 => to_unsigned(24009, LUT_AMPL_WIDTH - 1),
		8578 => to_unsigned(24011, LUT_AMPL_WIDTH - 1),
		8579 => to_unsigned(24013, LUT_AMPL_WIDTH - 1),
		8580 => to_unsigned(24015, LUT_AMPL_WIDTH - 1),
		8581 => to_unsigned(24018, LUT_AMPL_WIDTH - 1),
		8582 => to_unsigned(24020, LUT_AMPL_WIDTH - 1),
		8583 => to_unsigned(24022, LUT_AMPL_WIDTH - 1),
		8584 => to_unsigned(24024, LUT_AMPL_WIDTH - 1),
		8585 => to_unsigned(24026, LUT_AMPL_WIDTH - 1),
		8586 => to_unsigned(24028, LUT_AMPL_WIDTH - 1),
		8587 => to_unsigned(24030, LUT_AMPL_WIDTH - 1),
		8588 => to_unsigned(24033, LUT_AMPL_WIDTH - 1),
		8589 => to_unsigned(24035, LUT_AMPL_WIDTH - 1),
		8590 => to_unsigned(24037, LUT_AMPL_WIDTH - 1),
		8591 => to_unsigned(24039, LUT_AMPL_WIDTH - 1),
		8592 => to_unsigned(24041, LUT_AMPL_WIDTH - 1),
		8593 => to_unsigned(24043, LUT_AMPL_WIDTH - 1),
		8594 => to_unsigned(24045, LUT_AMPL_WIDTH - 1),
		8595 => to_unsigned(24047, LUT_AMPL_WIDTH - 1),
		8596 => to_unsigned(24050, LUT_AMPL_WIDTH - 1),
		8597 => to_unsigned(24052, LUT_AMPL_WIDTH - 1),
		8598 => to_unsigned(24054, LUT_AMPL_WIDTH - 1),
		8599 => to_unsigned(24056, LUT_AMPL_WIDTH - 1),
		8600 => to_unsigned(24058, LUT_AMPL_WIDTH - 1),
		8601 => to_unsigned(24060, LUT_AMPL_WIDTH - 1),
		8602 => to_unsigned(24062, LUT_AMPL_WIDTH - 1),
		8603 => to_unsigned(24065, LUT_AMPL_WIDTH - 1),
		8604 => to_unsigned(24067, LUT_AMPL_WIDTH - 1),
		8605 => to_unsigned(24069, LUT_AMPL_WIDTH - 1),
		8606 => to_unsigned(24071, LUT_AMPL_WIDTH - 1),
		8607 => to_unsigned(24073, LUT_AMPL_WIDTH - 1),
		8608 => to_unsigned(24075, LUT_AMPL_WIDTH - 1),
		8609 => to_unsigned(24077, LUT_AMPL_WIDTH - 1),
		8610 => to_unsigned(24079, LUT_AMPL_WIDTH - 1),
		8611 => to_unsigned(24082, LUT_AMPL_WIDTH - 1),
		8612 => to_unsigned(24084, LUT_AMPL_WIDTH - 1),
		8613 => to_unsigned(24086, LUT_AMPL_WIDTH - 1),
		8614 => to_unsigned(24088, LUT_AMPL_WIDTH - 1),
		8615 => to_unsigned(24090, LUT_AMPL_WIDTH - 1),
		8616 => to_unsigned(24092, LUT_AMPL_WIDTH - 1),
		8617 => to_unsigned(24094, LUT_AMPL_WIDTH - 1),
		8618 => to_unsigned(24096, LUT_AMPL_WIDTH - 1),
		8619 => to_unsigned(24099, LUT_AMPL_WIDTH - 1),
		8620 => to_unsigned(24101, LUT_AMPL_WIDTH - 1),
		8621 => to_unsigned(24103, LUT_AMPL_WIDTH - 1),
		8622 => to_unsigned(24105, LUT_AMPL_WIDTH - 1),
		8623 => to_unsigned(24107, LUT_AMPL_WIDTH - 1),
		8624 => to_unsigned(24109, LUT_AMPL_WIDTH - 1),
		8625 => to_unsigned(24111, LUT_AMPL_WIDTH - 1),
		8626 => to_unsigned(24114, LUT_AMPL_WIDTH - 1),
		8627 => to_unsigned(24116, LUT_AMPL_WIDTH - 1),
		8628 => to_unsigned(24118, LUT_AMPL_WIDTH - 1),
		8629 => to_unsigned(24120, LUT_AMPL_WIDTH - 1),
		8630 => to_unsigned(24122, LUT_AMPL_WIDTH - 1),
		8631 => to_unsigned(24124, LUT_AMPL_WIDTH - 1),
		8632 => to_unsigned(24126, LUT_AMPL_WIDTH - 1),
		8633 => to_unsigned(24128, LUT_AMPL_WIDTH - 1),
		8634 => to_unsigned(24131, LUT_AMPL_WIDTH - 1),
		8635 => to_unsigned(24133, LUT_AMPL_WIDTH - 1),
		8636 => to_unsigned(24135, LUT_AMPL_WIDTH - 1),
		8637 => to_unsigned(24137, LUT_AMPL_WIDTH - 1),
		8638 => to_unsigned(24139, LUT_AMPL_WIDTH - 1),
		8639 => to_unsigned(24141, LUT_AMPL_WIDTH - 1),
		8640 => to_unsigned(24143, LUT_AMPL_WIDTH - 1),
		8641 => to_unsigned(24145, LUT_AMPL_WIDTH - 1),
		8642 => to_unsigned(24148, LUT_AMPL_WIDTH - 1),
		8643 => to_unsigned(24150, LUT_AMPL_WIDTH - 1),
		8644 => to_unsigned(24152, LUT_AMPL_WIDTH - 1),
		8645 => to_unsigned(24154, LUT_AMPL_WIDTH - 1),
		8646 => to_unsigned(24156, LUT_AMPL_WIDTH - 1),
		8647 => to_unsigned(24158, LUT_AMPL_WIDTH - 1),
		8648 => to_unsigned(24160, LUT_AMPL_WIDTH - 1),
		8649 => to_unsigned(24162, LUT_AMPL_WIDTH - 1),
		8650 => to_unsigned(24164, LUT_AMPL_WIDTH - 1),
		8651 => to_unsigned(24167, LUT_AMPL_WIDTH - 1),
		8652 => to_unsigned(24169, LUT_AMPL_WIDTH - 1),
		8653 => to_unsigned(24171, LUT_AMPL_WIDTH - 1),
		8654 => to_unsigned(24173, LUT_AMPL_WIDTH - 1),
		8655 => to_unsigned(24175, LUT_AMPL_WIDTH - 1),
		8656 => to_unsigned(24177, LUT_AMPL_WIDTH - 1),
		8657 => to_unsigned(24179, LUT_AMPL_WIDTH - 1),
		8658 => to_unsigned(24181, LUT_AMPL_WIDTH - 1),
		8659 => to_unsigned(24184, LUT_AMPL_WIDTH - 1),
		8660 => to_unsigned(24186, LUT_AMPL_WIDTH - 1),
		8661 => to_unsigned(24188, LUT_AMPL_WIDTH - 1),
		8662 => to_unsigned(24190, LUT_AMPL_WIDTH - 1),
		8663 => to_unsigned(24192, LUT_AMPL_WIDTH - 1),
		8664 => to_unsigned(24194, LUT_AMPL_WIDTH - 1),
		8665 => to_unsigned(24196, LUT_AMPL_WIDTH - 1),
		8666 => to_unsigned(24198, LUT_AMPL_WIDTH - 1),
		8667 => to_unsigned(24201, LUT_AMPL_WIDTH - 1),
		8668 => to_unsigned(24203, LUT_AMPL_WIDTH - 1),
		8669 => to_unsigned(24205, LUT_AMPL_WIDTH - 1),
		8670 => to_unsigned(24207, LUT_AMPL_WIDTH - 1),
		8671 => to_unsigned(24209, LUT_AMPL_WIDTH - 1),
		8672 => to_unsigned(24211, LUT_AMPL_WIDTH - 1),
		8673 => to_unsigned(24213, LUT_AMPL_WIDTH - 1),
		8674 => to_unsigned(24215, LUT_AMPL_WIDTH - 1),
		8675 => to_unsigned(24217, LUT_AMPL_WIDTH - 1),
		8676 => to_unsigned(24220, LUT_AMPL_WIDTH - 1),
		8677 => to_unsigned(24222, LUT_AMPL_WIDTH - 1),
		8678 => to_unsigned(24224, LUT_AMPL_WIDTH - 1),
		8679 => to_unsigned(24226, LUT_AMPL_WIDTH - 1),
		8680 => to_unsigned(24228, LUT_AMPL_WIDTH - 1),
		8681 => to_unsigned(24230, LUT_AMPL_WIDTH - 1),
		8682 => to_unsigned(24232, LUT_AMPL_WIDTH - 1),
		8683 => to_unsigned(24234, LUT_AMPL_WIDTH - 1),
		8684 => to_unsigned(24237, LUT_AMPL_WIDTH - 1),
		8685 => to_unsigned(24239, LUT_AMPL_WIDTH - 1),
		8686 => to_unsigned(24241, LUT_AMPL_WIDTH - 1),
		8687 => to_unsigned(24243, LUT_AMPL_WIDTH - 1),
		8688 => to_unsigned(24245, LUT_AMPL_WIDTH - 1),
		8689 => to_unsigned(24247, LUT_AMPL_WIDTH - 1),
		8690 => to_unsigned(24249, LUT_AMPL_WIDTH - 1),
		8691 => to_unsigned(24251, LUT_AMPL_WIDTH - 1),
		8692 => to_unsigned(24253, LUT_AMPL_WIDTH - 1),
		8693 => to_unsigned(24256, LUT_AMPL_WIDTH - 1),
		8694 => to_unsigned(24258, LUT_AMPL_WIDTH - 1),
		8695 => to_unsigned(24260, LUT_AMPL_WIDTH - 1),
		8696 => to_unsigned(24262, LUT_AMPL_WIDTH - 1),
		8697 => to_unsigned(24264, LUT_AMPL_WIDTH - 1),
		8698 => to_unsigned(24266, LUT_AMPL_WIDTH - 1),
		8699 => to_unsigned(24268, LUT_AMPL_WIDTH - 1),
		8700 => to_unsigned(24270, LUT_AMPL_WIDTH - 1),
		8701 => to_unsigned(24272, LUT_AMPL_WIDTH - 1),
		8702 => to_unsigned(24275, LUT_AMPL_WIDTH - 1),
		8703 => to_unsigned(24277, LUT_AMPL_WIDTH - 1),
		8704 => to_unsigned(24279, LUT_AMPL_WIDTH - 1),
		8705 => to_unsigned(24281, LUT_AMPL_WIDTH - 1),
		8706 => to_unsigned(24283, LUT_AMPL_WIDTH - 1),
		8707 => to_unsigned(24285, LUT_AMPL_WIDTH - 1),
		8708 => to_unsigned(24287, LUT_AMPL_WIDTH - 1),
		8709 => to_unsigned(24289, LUT_AMPL_WIDTH - 1),
		8710 => to_unsigned(24291, LUT_AMPL_WIDTH - 1),
		8711 => to_unsigned(24294, LUT_AMPL_WIDTH - 1),
		8712 => to_unsigned(24296, LUT_AMPL_WIDTH - 1),
		8713 => to_unsigned(24298, LUT_AMPL_WIDTH - 1),
		8714 => to_unsigned(24300, LUT_AMPL_WIDTH - 1),
		8715 => to_unsigned(24302, LUT_AMPL_WIDTH - 1),
		8716 => to_unsigned(24304, LUT_AMPL_WIDTH - 1),
		8717 => to_unsigned(24306, LUT_AMPL_WIDTH - 1),
		8718 => to_unsigned(24308, LUT_AMPL_WIDTH - 1),
		8719 => to_unsigned(24310, LUT_AMPL_WIDTH - 1),
		8720 => to_unsigned(24312, LUT_AMPL_WIDTH - 1),
		8721 => to_unsigned(24315, LUT_AMPL_WIDTH - 1),
		8722 => to_unsigned(24317, LUT_AMPL_WIDTH - 1),
		8723 => to_unsigned(24319, LUT_AMPL_WIDTH - 1),
		8724 => to_unsigned(24321, LUT_AMPL_WIDTH - 1),
		8725 => to_unsigned(24323, LUT_AMPL_WIDTH - 1),
		8726 => to_unsigned(24325, LUT_AMPL_WIDTH - 1),
		8727 => to_unsigned(24327, LUT_AMPL_WIDTH - 1),
		8728 => to_unsigned(24329, LUT_AMPL_WIDTH - 1),
		8729 => to_unsigned(24331, LUT_AMPL_WIDTH - 1),
		8730 => to_unsigned(24334, LUT_AMPL_WIDTH - 1),
		8731 => to_unsigned(24336, LUT_AMPL_WIDTH - 1),
		8732 => to_unsigned(24338, LUT_AMPL_WIDTH - 1),
		8733 => to_unsigned(24340, LUT_AMPL_WIDTH - 1),
		8734 => to_unsigned(24342, LUT_AMPL_WIDTH - 1),
		8735 => to_unsigned(24344, LUT_AMPL_WIDTH - 1),
		8736 => to_unsigned(24346, LUT_AMPL_WIDTH - 1),
		8737 => to_unsigned(24348, LUT_AMPL_WIDTH - 1),
		8738 => to_unsigned(24350, LUT_AMPL_WIDTH - 1),
		8739 => to_unsigned(24352, LUT_AMPL_WIDTH - 1),
		8740 => to_unsigned(24355, LUT_AMPL_WIDTH - 1),
		8741 => to_unsigned(24357, LUT_AMPL_WIDTH - 1),
		8742 => to_unsigned(24359, LUT_AMPL_WIDTH - 1),
		8743 => to_unsigned(24361, LUT_AMPL_WIDTH - 1),
		8744 => to_unsigned(24363, LUT_AMPL_WIDTH - 1),
		8745 => to_unsigned(24365, LUT_AMPL_WIDTH - 1),
		8746 => to_unsigned(24367, LUT_AMPL_WIDTH - 1),
		8747 => to_unsigned(24369, LUT_AMPL_WIDTH - 1),
		8748 => to_unsigned(24371, LUT_AMPL_WIDTH - 1),
		8749 => to_unsigned(24373, LUT_AMPL_WIDTH - 1),
		8750 => to_unsigned(24376, LUT_AMPL_WIDTH - 1),
		8751 => to_unsigned(24378, LUT_AMPL_WIDTH - 1),
		8752 => to_unsigned(24380, LUT_AMPL_WIDTH - 1),
		8753 => to_unsigned(24382, LUT_AMPL_WIDTH - 1),
		8754 => to_unsigned(24384, LUT_AMPL_WIDTH - 1),
		8755 => to_unsigned(24386, LUT_AMPL_WIDTH - 1),
		8756 => to_unsigned(24388, LUT_AMPL_WIDTH - 1),
		8757 => to_unsigned(24390, LUT_AMPL_WIDTH - 1),
		8758 => to_unsigned(24392, LUT_AMPL_WIDTH - 1),
		8759 => to_unsigned(24394, LUT_AMPL_WIDTH - 1),
		8760 => to_unsigned(24397, LUT_AMPL_WIDTH - 1),
		8761 => to_unsigned(24399, LUT_AMPL_WIDTH - 1),
		8762 => to_unsigned(24401, LUT_AMPL_WIDTH - 1),
		8763 => to_unsigned(24403, LUT_AMPL_WIDTH - 1),
		8764 => to_unsigned(24405, LUT_AMPL_WIDTH - 1),
		8765 => to_unsigned(24407, LUT_AMPL_WIDTH - 1),
		8766 => to_unsigned(24409, LUT_AMPL_WIDTH - 1),
		8767 => to_unsigned(24411, LUT_AMPL_WIDTH - 1),
		8768 => to_unsigned(24413, LUT_AMPL_WIDTH - 1),
		8769 => to_unsigned(24415, LUT_AMPL_WIDTH - 1),
		8770 => to_unsigned(24417, LUT_AMPL_WIDTH - 1),
		8771 => to_unsigned(24420, LUT_AMPL_WIDTH - 1),
		8772 => to_unsigned(24422, LUT_AMPL_WIDTH - 1),
		8773 => to_unsigned(24424, LUT_AMPL_WIDTH - 1),
		8774 => to_unsigned(24426, LUT_AMPL_WIDTH - 1),
		8775 => to_unsigned(24428, LUT_AMPL_WIDTH - 1),
		8776 => to_unsigned(24430, LUT_AMPL_WIDTH - 1),
		8777 => to_unsigned(24432, LUT_AMPL_WIDTH - 1),
		8778 => to_unsigned(24434, LUT_AMPL_WIDTH - 1),
		8779 => to_unsigned(24436, LUT_AMPL_WIDTH - 1),
		8780 => to_unsigned(24438, LUT_AMPL_WIDTH - 1),
		8781 => to_unsigned(24441, LUT_AMPL_WIDTH - 1),
		8782 => to_unsigned(24443, LUT_AMPL_WIDTH - 1),
		8783 => to_unsigned(24445, LUT_AMPL_WIDTH - 1),
		8784 => to_unsigned(24447, LUT_AMPL_WIDTH - 1),
		8785 => to_unsigned(24449, LUT_AMPL_WIDTH - 1),
		8786 => to_unsigned(24451, LUT_AMPL_WIDTH - 1),
		8787 => to_unsigned(24453, LUT_AMPL_WIDTH - 1),
		8788 => to_unsigned(24455, LUT_AMPL_WIDTH - 1),
		8789 => to_unsigned(24457, LUT_AMPL_WIDTH - 1),
		8790 => to_unsigned(24459, LUT_AMPL_WIDTH - 1),
		8791 => to_unsigned(24461, LUT_AMPL_WIDTH - 1),
		8792 => to_unsigned(24464, LUT_AMPL_WIDTH - 1),
		8793 => to_unsigned(24466, LUT_AMPL_WIDTH - 1),
		8794 => to_unsigned(24468, LUT_AMPL_WIDTH - 1),
		8795 => to_unsigned(24470, LUT_AMPL_WIDTH - 1),
		8796 => to_unsigned(24472, LUT_AMPL_WIDTH - 1),
		8797 => to_unsigned(24474, LUT_AMPL_WIDTH - 1),
		8798 => to_unsigned(24476, LUT_AMPL_WIDTH - 1),
		8799 => to_unsigned(24478, LUT_AMPL_WIDTH - 1),
		8800 => to_unsigned(24480, LUT_AMPL_WIDTH - 1),
		8801 => to_unsigned(24482, LUT_AMPL_WIDTH - 1),
		8802 => to_unsigned(24484, LUT_AMPL_WIDTH - 1),
		8803 => to_unsigned(24487, LUT_AMPL_WIDTH - 1),
		8804 => to_unsigned(24489, LUT_AMPL_WIDTH - 1),
		8805 => to_unsigned(24491, LUT_AMPL_WIDTH - 1),
		8806 => to_unsigned(24493, LUT_AMPL_WIDTH - 1),
		8807 => to_unsigned(24495, LUT_AMPL_WIDTH - 1),
		8808 => to_unsigned(24497, LUT_AMPL_WIDTH - 1),
		8809 => to_unsigned(24499, LUT_AMPL_WIDTH - 1),
		8810 => to_unsigned(24501, LUT_AMPL_WIDTH - 1),
		8811 => to_unsigned(24503, LUT_AMPL_WIDTH - 1),
		8812 => to_unsigned(24505, LUT_AMPL_WIDTH - 1),
		8813 => to_unsigned(24507, LUT_AMPL_WIDTH - 1),
		8814 => to_unsigned(24509, LUT_AMPL_WIDTH - 1),
		8815 => to_unsigned(24512, LUT_AMPL_WIDTH - 1),
		8816 => to_unsigned(24514, LUT_AMPL_WIDTH - 1),
		8817 => to_unsigned(24516, LUT_AMPL_WIDTH - 1),
		8818 => to_unsigned(24518, LUT_AMPL_WIDTH - 1),
		8819 => to_unsigned(24520, LUT_AMPL_WIDTH - 1),
		8820 => to_unsigned(24522, LUT_AMPL_WIDTH - 1),
		8821 => to_unsigned(24524, LUT_AMPL_WIDTH - 1),
		8822 => to_unsigned(24526, LUT_AMPL_WIDTH - 1),
		8823 => to_unsigned(24528, LUT_AMPL_WIDTH - 1),
		8824 => to_unsigned(24530, LUT_AMPL_WIDTH - 1),
		8825 => to_unsigned(24532, LUT_AMPL_WIDTH - 1),
		8826 => to_unsigned(24534, LUT_AMPL_WIDTH - 1),
		8827 => to_unsigned(24537, LUT_AMPL_WIDTH - 1),
		8828 => to_unsigned(24539, LUT_AMPL_WIDTH - 1),
		8829 => to_unsigned(24541, LUT_AMPL_WIDTH - 1),
		8830 => to_unsigned(24543, LUT_AMPL_WIDTH - 1),
		8831 => to_unsigned(24545, LUT_AMPL_WIDTH - 1),
		8832 => to_unsigned(24547, LUT_AMPL_WIDTH - 1),
		8833 => to_unsigned(24549, LUT_AMPL_WIDTH - 1),
		8834 => to_unsigned(24551, LUT_AMPL_WIDTH - 1),
		8835 => to_unsigned(24553, LUT_AMPL_WIDTH - 1),
		8836 => to_unsigned(24555, LUT_AMPL_WIDTH - 1),
		8837 => to_unsigned(24557, LUT_AMPL_WIDTH - 1),
		8838 => to_unsigned(24559, LUT_AMPL_WIDTH - 1),
		8839 => to_unsigned(24562, LUT_AMPL_WIDTH - 1),
		8840 => to_unsigned(24564, LUT_AMPL_WIDTH - 1),
		8841 => to_unsigned(24566, LUT_AMPL_WIDTH - 1),
		8842 => to_unsigned(24568, LUT_AMPL_WIDTH - 1),
		8843 => to_unsigned(24570, LUT_AMPL_WIDTH - 1),
		8844 => to_unsigned(24572, LUT_AMPL_WIDTH - 1),
		8845 => to_unsigned(24574, LUT_AMPL_WIDTH - 1),
		8846 => to_unsigned(24576, LUT_AMPL_WIDTH - 1),
		8847 => to_unsigned(24578, LUT_AMPL_WIDTH - 1),
		8848 => to_unsigned(24580, LUT_AMPL_WIDTH - 1),
		8849 => to_unsigned(24582, LUT_AMPL_WIDTH - 1),
		8850 => to_unsigned(24584, LUT_AMPL_WIDTH - 1),
		8851 => to_unsigned(24586, LUT_AMPL_WIDTH - 1),
		8852 => to_unsigned(24589, LUT_AMPL_WIDTH - 1),
		8853 => to_unsigned(24591, LUT_AMPL_WIDTH - 1),
		8854 => to_unsigned(24593, LUT_AMPL_WIDTH - 1),
		8855 => to_unsigned(24595, LUT_AMPL_WIDTH - 1),
		8856 => to_unsigned(24597, LUT_AMPL_WIDTH - 1),
		8857 => to_unsigned(24599, LUT_AMPL_WIDTH - 1),
		8858 => to_unsigned(24601, LUT_AMPL_WIDTH - 1),
		8859 => to_unsigned(24603, LUT_AMPL_WIDTH - 1),
		8860 => to_unsigned(24605, LUT_AMPL_WIDTH - 1),
		8861 => to_unsigned(24607, LUT_AMPL_WIDTH - 1),
		8862 => to_unsigned(24609, LUT_AMPL_WIDTH - 1),
		8863 => to_unsigned(24611, LUT_AMPL_WIDTH - 1),
		8864 => to_unsigned(24613, LUT_AMPL_WIDTH - 1),
		8865 => to_unsigned(24616, LUT_AMPL_WIDTH - 1),
		8866 => to_unsigned(24618, LUT_AMPL_WIDTH - 1),
		8867 => to_unsigned(24620, LUT_AMPL_WIDTH - 1),
		8868 => to_unsigned(24622, LUT_AMPL_WIDTH - 1),
		8869 => to_unsigned(24624, LUT_AMPL_WIDTH - 1),
		8870 => to_unsigned(24626, LUT_AMPL_WIDTH - 1),
		8871 => to_unsigned(24628, LUT_AMPL_WIDTH - 1),
		8872 => to_unsigned(24630, LUT_AMPL_WIDTH - 1),
		8873 => to_unsigned(24632, LUT_AMPL_WIDTH - 1),
		8874 => to_unsigned(24634, LUT_AMPL_WIDTH - 1),
		8875 => to_unsigned(24636, LUT_AMPL_WIDTH - 1),
		8876 => to_unsigned(24638, LUT_AMPL_WIDTH - 1),
		8877 => to_unsigned(24640, LUT_AMPL_WIDTH - 1),
		8878 => to_unsigned(24642, LUT_AMPL_WIDTH - 1),
		8879 => to_unsigned(24645, LUT_AMPL_WIDTH - 1),
		8880 => to_unsigned(24647, LUT_AMPL_WIDTH - 1),
		8881 => to_unsigned(24649, LUT_AMPL_WIDTH - 1),
		8882 => to_unsigned(24651, LUT_AMPL_WIDTH - 1),
		8883 => to_unsigned(24653, LUT_AMPL_WIDTH - 1),
		8884 => to_unsigned(24655, LUT_AMPL_WIDTH - 1),
		8885 => to_unsigned(24657, LUT_AMPL_WIDTH - 1),
		8886 => to_unsigned(24659, LUT_AMPL_WIDTH - 1),
		8887 => to_unsigned(24661, LUT_AMPL_WIDTH - 1),
		8888 => to_unsigned(24663, LUT_AMPL_WIDTH - 1),
		8889 => to_unsigned(24665, LUT_AMPL_WIDTH - 1),
		8890 => to_unsigned(24667, LUT_AMPL_WIDTH - 1),
		8891 => to_unsigned(24669, LUT_AMPL_WIDTH - 1),
		8892 => to_unsigned(24671, LUT_AMPL_WIDTH - 1),
		8893 => to_unsigned(24673, LUT_AMPL_WIDTH - 1),
		8894 => to_unsigned(24676, LUT_AMPL_WIDTH - 1),
		8895 => to_unsigned(24678, LUT_AMPL_WIDTH - 1),
		8896 => to_unsigned(24680, LUT_AMPL_WIDTH - 1),
		8897 => to_unsigned(24682, LUT_AMPL_WIDTH - 1),
		8898 => to_unsigned(24684, LUT_AMPL_WIDTH - 1),
		8899 => to_unsigned(24686, LUT_AMPL_WIDTH - 1),
		8900 => to_unsigned(24688, LUT_AMPL_WIDTH - 1),
		8901 => to_unsigned(24690, LUT_AMPL_WIDTH - 1),
		8902 => to_unsigned(24692, LUT_AMPL_WIDTH - 1),
		8903 => to_unsigned(24694, LUT_AMPL_WIDTH - 1),
		8904 => to_unsigned(24696, LUT_AMPL_WIDTH - 1),
		8905 => to_unsigned(24698, LUT_AMPL_WIDTH - 1),
		8906 => to_unsigned(24700, LUT_AMPL_WIDTH - 1),
		8907 => to_unsigned(24702, LUT_AMPL_WIDTH - 1),
		8908 => to_unsigned(24704, LUT_AMPL_WIDTH - 1),
		8909 => to_unsigned(24707, LUT_AMPL_WIDTH - 1),
		8910 => to_unsigned(24709, LUT_AMPL_WIDTH - 1),
		8911 => to_unsigned(24711, LUT_AMPL_WIDTH - 1),
		8912 => to_unsigned(24713, LUT_AMPL_WIDTH - 1),
		8913 => to_unsigned(24715, LUT_AMPL_WIDTH - 1),
		8914 => to_unsigned(24717, LUT_AMPL_WIDTH - 1),
		8915 => to_unsigned(24719, LUT_AMPL_WIDTH - 1),
		8916 => to_unsigned(24721, LUT_AMPL_WIDTH - 1),
		8917 => to_unsigned(24723, LUT_AMPL_WIDTH - 1),
		8918 => to_unsigned(24725, LUT_AMPL_WIDTH - 1),
		8919 => to_unsigned(24727, LUT_AMPL_WIDTH - 1),
		8920 => to_unsigned(24729, LUT_AMPL_WIDTH - 1),
		8921 => to_unsigned(24731, LUT_AMPL_WIDTH - 1),
		8922 => to_unsigned(24733, LUT_AMPL_WIDTH - 1),
		8923 => to_unsigned(24735, LUT_AMPL_WIDTH - 1),
		8924 => to_unsigned(24737, LUT_AMPL_WIDTH - 1),
		8925 => to_unsigned(24740, LUT_AMPL_WIDTH - 1),
		8926 => to_unsigned(24742, LUT_AMPL_WIDTH - 1),
		8927 => to_unsigned(24744, LUT_AMPL_WIDTH - 1),
		8928 => to_unsigned(24746, LUT_AMPL_WIDTH - 1),
		8929 => to_unsigned(24748, LUT_AMPL_WIDTH - 1),
		8930 => to_unsigned(24750, LUT_AMPL_WIDTH - 1),
		8931 => to_unsigned(24752, LUT_AMPL_WIDTH - 1),
		8932 => to_unsigned(24754, LUT_AMPL_WIDTH - 1),
		8933 => to_unsigned(24756, LUT_AMPL_WIDTH - 1),
		8934 => to_unsigned(24758, LUT_AMPL_WIDTH - 1),
		8935 => to_unsigned(24760, LUT_AMPL_WIDTH - 1),
		8936 => to_unsigned(24762, LUT_AMPL_WIDTH - 1),
		8937 => to_unsigned(24764, LUT_AMPL_WIDTH - 1),
		8938 => to_unsigned(24766, LUT_AMPL_WIDTH - 1),
		8939 => to_unsigned(24768, LUT_AMPL_WIDTH - 1),
		8940 => to_unsigned(24770, LUT_AMPL_WIDTH - 1),
		8941 => to_unsigned(24772, LUT_AMPL_WIDTH - 1),
		8942 => to_unsigned(24774, LUT_AMPL_WIDTH - 1),
		8943 => to_unsigned(24777, LUT_AMPL_WIDTH - 1),
		8944 => to_unsigned(24779, LUT_AMPL_WIDTH - 1),
		8945 => to_unsigned(24781, LUT_AMPL_WIDTH - 1),
		8946 => to_unsigned(24783, LUT_AMPL_WIDTH - 1),
		8947 => to_unsigned(24785, LUT_AMPL_WIDTH - 1),
		8948 => to_unsigned(24787, LUT_AMPL_WIDTH - 1),
		8949 => to_unsigned(24789, LUT_AMPL_WIDTH - 1),
		8950 => to_unsigned(24791, LUT_AMPL_WIDTH - 1),
		8951 => to_unsigned(24793, LUT_AMPL_WIDTH - 1),
		8952 => to_unsigned(24795, LUT_AMPL_WIDTH - 1),
		8953 => to_unsigned(24797, LUT_AMPL_WIDTH - 1),
		8954 => to_unsigned(24799, LUT_AMPL_WIDTH - 1),
		8955 => to_unsigned(24801, LUT_AMPL_WIDTH - 1),
		8956 => to_unsigned(24803, LUT_AMPL_WIDTH - 1),
		8957 => to_unsigned(24805, LUT_AMPL_WIDTH - 1),
		8958 => to_unsigned(24807, LUT_AMPL_WIDTH - 1),
		8959 => to_unsigned(24809, LUT_AMPL_WIDTH - 1),
		8960 => to_unsigned(24811, LUT_AMPL_WIDTH - 1),
		8961 => to_unsigned(24814, LUT_AMPL_WIDTH - 1),
		8962 => to_unsigned(24816, LUT_AMPL_WIDTH - 1),
		8963 => to_unsigned(24818, LUT_AMPL_WIDTH - 1),
		8964 => to_unsigned(24820, LUT_AMPL_WIDTH - 1),
		8965 => to_unsigned(24822, LUT_AMPL_WIDTH - 1),
		8966 => to_unsigned(24824, LUT_AMPL_WIDTH - 1),
		8967 => to_unsigned(24826, LUT_AMPL_WIDTH - 1),
		8968 => to_unsigned(24828, LUT_AMPL_WIDTH - 1),
		8969 => to_unsigned(24830, LUT_AMPL_WIDTH - 1),
		8970 => to_unsigned(24832, LUT_AMPL_WIDTH - 1),
		8971 => to_unsigned(24834, LUT_AMPL_WIDTH - 1),
		8972 => to_unsigned(24836, LUT_AMPL_WIDTH - 1),
		8973 => to_unsigned(24838, LUT_AMPL_WIDTH - 1),
		8974 => to_unsigned(24840, LUT_AMPL_WIDTH - 1),
		8975 => to_unsigned(24842, LUT_AMPL_WIDTH - 1),
		8976 => to_unsigned(24844, LUT_AMPL_WIDTH - 1),
		8977 => to_unsigned(24846, LUT_AMPL_WIDTH - 1),
		8978 => to_unsigned(24848, LUT_AMPL_WIDTH - 1),
		8979 => to_unsigned(24850, LUT_AMPL_WIDTH - 1),
		8980 => to_unsigned(24852, LUT_AMPL_WIDTH - 1),
		8981 => to_unsigned(24855, LUT_AMPL_WIDTH - 1),
		8982 => to_unsigned(24857, LUT_AMPL_WIDTH - 1),
		8983 => to_unsigned(24859, LUT_AMPL_WIDTH - 1),
		8984 => to_unsigned(24861, LUT_AMPL_WIDTH - 1),
		8985 => to_unsigned(24863, LUT_AMPL_WIDTH - 1),
		8986 => to_unsigned(24865, LUT_AMPL_WIDTH - 1),
		8987 => to_unsigned(24867, LUT_AMPL_WIDTH - 1),
		8988 => to_unsigned(24869, LUT_AMPL_WIDTH - 1),
		8989 => to_unsigned(24871, LUT_AMPL_WIDTH - 1),
		8990 => to_unsigned(24873, LUT_AMPL_WIDTH - 1),
		8991 => to_unsigned(24875, LUT_AMPL_WIDTH - 1),
		8992 => to_unsigned(24877, LUT_AMPL_WIDTH - 1),
		8993 => to_unsigned(24879, LUT_AMPL_WIDTH - 1),
		8994 => to_unsigned(24881, LUT_AMPL_WIDTH - 1),
		8995 => to_unsigned(24883, LUT_AMPL_WIDTH - 1),
		8996 => to_unsigned(24885, LUT_AMPL_WIDTH - 1),
		8997 => to_unsigned(24887, LUT_AMPL_WIDTH - 1),
		8998 => to_unsigned(24889, LUT_AMPL_WIDTH - 1),
		8999 => to_unsigned(24891, LUT_AMPL_WIDTH - 1),
		9000 => to_unsigned(24893, LUT_AMPL_WIDTH - 1),
		9001 => to_unsigned(24895, LUT_AMPL_WIDTH - 1),
		9002 => to_unsigned(24897, LUT_AMPL_WIDTH - 1),
		9003 => to_unsigned(24899, LUT_AMPL_WIDTH - 1),
		9004 => to_unsigned(24902, LUT_AMPL_WIDTH - 1),
		9005 => to_unsigned(24904, LUT_AMPL_WIDTH - 1),
		9006 => to_unsigned(24906, LUT_AMPL_WIDTH - 1),
		9007 => to_unsigned(24908, LUT_AMPL_WIDTH - 1),
		9008 => to_unsigned(24910, LUT_AMPL_WIDTH - 1),
		9009 => to_unsigned(24912, LUT_AMPL_WIDTH - 1),
		9010 => to_unsigned(24914, LUT_AMPL_WIDTH - 1),
		9011 => to_unsigned(24916, LUT_AMPL_WIDTH - 1),
		9012 => to_unsigned(24918, LUT_AMPL_WIDTH - 1),
		9013 => to_unsigned(24920, LUT_AMPL_WIDTH - 1),
		9014 => to_unsigned(24922, LUT_AMPL_WIDTH - 1),
		9015 => to_unsigned(24924, LUT_AMPL_WIDTH - 1),
		9016 => to_unsigned(24926, LUT_AMPL_WIDTH - 1),
		9017 => to_unsigned(24928, LUT_AMPL_WIDTH - 1),
		9018 => to_unsigned(24930, LUT_AMPL_WIDTH - 1),
		9019 => to_unsigned(24932, LUT_AMPL_WIDTH - 1),
		9020 => to_unsigned(24934, LUT_AMPL_WIDTH - 1),
		9021 => to_unsigned(24936, LUT_AMPL_WIDTH - 1),
		9022 => to_unsigned(24938, LUT_AMPL_WIDTH - 1),
		9023 => to_unsigned(24940, LUT_AMPL_WIDTH - 1),
		9024 => to_unsigned(24942, LUT_AMPL_WIDTH - 1),
		9025 => to_unsigned(24944, LUT_AMPL_WIDTH - 1),
		9026 => to_unsigned(24946, LUT_AMPL_WIDTH - 1),
		9027 => to_unsigned(24948, LUT_AMPL_WIDTH - 1),
		9028 => to_unsigned(24950, LUT_AMPL_WIDTH - 1),
		9029 => to_unsigned(24953, LUT_AMPL_WIDTH - 1),
		9030 => to_unsigned(24955, LUT_AMPL_WIDTH - 1),
		9031 => to_unsigned(24957, LUT_AMPL_WIDTH - 1),
		9032 => to_unsigned(24959, LUT_AMPL_WIDTH - 1),
		9033 => to_unsigned(24961, LUT_AMPL_WIDTH - 1),
		9034 => to_unsigned(24963, LUT_AMPL_WIDTH - 1),
		9035 => to_unsigned(24965, LUT_AMPL_WIDTH - 1),
		9036 => to_unsigned(24967, LUT_AMPL_WIDTH - 1),
		9037 => to_unsigned(24969, LUT_AMPL_WIDTH - 1),
		9038 => to_unsigned(24971, LUT_AMPL_WIDTH - 1),
		9039 => to_unsigned(24973, LUT_AMPL_WIDTH - 1),
		9040 => to_unsigned(24975, LUT_AMPL_WIDTH - 1),
		9041 => to_unsigned(24977, LUT_AMPL_WIDTH - 1),
		9042 => to_unsigned(24979, LUT_AMPL_WIDTH - 1),
		9043 => to_unsigned(24981, LUT_AMPL_WIDTH - 1),
		9044 => to_unsigned(24983, LUT_AMPL_WIDTH - 1),
		9045 => to_unsigned(24985, LUT_AMPL_WIDTH - 1),
		9046 => to_unsigned(24987, LUT_AMPL_WIDTH - 1),
		9047 => to_unsigned(24989, LUT_AMPL_WIDTH - 1),
		9048 => to_unsigned(24991, LUT_AMPL_WIDTH - 1),
		9049 => to_unsigned(24993, LUT_AMPL_WIDTH - 1),
		9050 => to_unsigned(24995, LUT_AMPL_WIDTH - 1),
		9051 => to_unsigned(24997, LUT_AMPL_WIDTH - 1),
		9052 => to_unsigned(24999, LUT_AMPL_WIDTH - 1),
		9053 => to_unsigned(25001, LUT_AMPL_WIDTH - 1),
		9054 => to_unsigned(25003, LUT_AMPL_WIDTH - 1),
		9055 => to_unsigned(25005, LUT_AMPL_WIDTH - 1),
		9056 => to_unsigned(25007, LUT_AMPL_WIDTH - 1),
		9057 => to_unsigned(25009, LUT_AMPL_WIDTH - 1),
		9058 => to_unsigned(25011, LUT_AMPL_WIDTH - 1),
		9059 => to_unsigned(25013, LUT_AMPL_WIDTH - 1),
		9060 => to_unsigned(25016, LUT_AMPL_WIDTH - 1),
		9061 => to_unsigned(25018, LUT_AMPL_WIDTH - 1),
		9062 => to_unsigned(25020, LUT_AMPL_WIDTH - 1),
		9063 => to_unsigned(25022, LUT_AMPL_WIDTH - 1),
		9064 => to_unsigned(25024, LUT_AMPL_WIDTH - 1),
		9065 => to_unsigned(25026, LUT_AMPL_WIDTH - 1),
		9066 => to_unsigned(25028, LUT_AMPL_WIDTH - 1),
		9067 => to_unsigned(25030, LUT_AMPL_WIDTH - 1),
		9068 => to_unsigned(25032, LUT_AMPL_WIDTH - 1),
		9069 => to_unsigned(25034, LUT_AMPL_WIDTH - 1),
		9070 => to_unsigned(25036, LUT_AMPL_WIDTH - 1),
		9071 => to_unsigned(25038, LUT_AMPL_WIDTH - 1),
		9072 => to_unsigned(25040, LUT_AMPL_WIDTH - 1),
		9073 => to_unsigned(25042, LUT_AMPL_WIDTH - 1),
		9074 => to_unsigned(25044, LUT_AMPL_WIDTH - 1),
		9075 => to_unsigned(25046, LUT_AMPL_WIDTH - 1),
		9076 => to_unsigned(25048, LUT_AMPL_WIDTH - 1),
		9077 => to_unsigned(25050, LUT_AMPL_WIDTH - 1),
		9078 => to_unsigned(25052, LUT_AMPL_WIDTH - 1),
		9079 => to_unsigned(25054, LUT_AMPL_WIDTH - 1),
		9080 => to_unsigned(25056, LUT_AMPL_WIDTH - 1),
		9081 => to_unsigned(25058, LUT_AMPL_WIDTH - 1),
		9082 => to_unsigned(25060, LUT_AMPL_WIDTH - 1),
		9083 => to_unsigned(25062, LUT_AMPL_WIDTH - 1),
		9084 => to_unsigned(25064, LUT_AMPL_WIDTH - 1),
		9085 => to_unsigned(25066, LUT_AMPL_WIDTH - 1),
		9086 => to_unsigned(25068, LUT_AMPL_WIDTH - 1),
		9087 => to_unsigned(25070, LUT_AMPL_WIDTH - 1),
		9088 => to_unsigned(25072, LUT_AMPL_WIDTH - 1),
		9089 => to_unsigned(25074, LUT_AMPL_WIDTH - 1),
		9090 => to_unsigned(25076, LUT_AMPL_WIDTH - 1),
		9091 => to_unsigned(25078, LUT_AMPL_WIDTH - 1),
		9092 => to_unsigned(25080, LUT_AMPL_WIDTH - 1),
		9093 => to_unsigned(25082, LUT_AMPL_WIDTH - 1),
		9094 => to_unsigned(25084, LUT_AMPL_WIDTH - 1),
		9095 => to_unsigned(25086, LUT_AMPL_WIDTH - 1),
		9096 => to_unsigned(25088, LUT_AMPL_WIDTH - 1),
		9097 => to_unsigned(25090, LUT_AMPL_WIDTH - 1),
		9098 => to_unsigned(25092, LUT_AMPL_WIDTH - 1),
		9099 => to_unsigned(25094, LUT_AMPL_WIDTH - 1),
		9100 => to_unsigned(25096, LUT_AMPL_WIDTH - 1),
		9101 => to_unsigned(25099, LUT_AMPL_WIDTH - 1),
		9102 => to_unsigned(25101, LUT_AMPL_WIDTH - 1),
		9103 => to_unsigned(25103, LUT_AMPL_WIDTH - 1),
		9104 => to_unsigned(25105, LUT_AMPL_WIDTH - 1),
		9105 => to_unsigned(25107, LUT_AMPL_WIDTH - 1),
		9106 => to_unsigned(25109, LUT_AMPL_WIDTH - 1),
		9107 => to_unsigned(25111, LUT_AMPL_WIDTH - 1),
		9108 => to_unsigned(25113, LUT_AMPL_WIDTH - 1),
		9109 => to_unsigned(25115, LUT_AMPL_WIDTH - 1),
		9110 => to_unsigned(25117, LUT_AMPL_WIDTH - 1),
		9111 => to_unsigned(25119, LUT_AMPL_WIDTH - 1),
		9112 => to_unsigned(25121, LUT_AMPL_WIDTH - 1),
		9113 => to_unsigned(25123, LUT_AMPL_WIDTH - 1),
		9114 => to_unsigned(25125, LUT_AMPL_WIDTH - 1),
		9115 => to_unsigned(25127, LUT_AMPL_WIDTH - 1),
		9116 => to_unsigned(25129, LUT_AMPL_WIDTH - 1),
		9117 => to_unsigned(25131, LUT_AMPL_WIDTH - 1),
		9118 => to_unsigned(25133, LUT_AMPL_WIDTH - 1),
		9119 => to_unsigned(25135, LUT_AMPL_WIDTH - 1),
		9120 => to_unsigned(25137, LUT_AMPL_WIDTH - 1),
		9121 => to_unsigned(25139, LUT_AMPL_WIDTH - 1),
		9122 => to_unsigned(25141, LUT_AMPL_WIDTH - 1),
		9123 => to_unsigned(25143, LUT_AMPL_WIDTH - 1),
		9124 => to_unsigned(25145, LUT_AMPL_WIDTH - 1),
		9125 => to_unsigned(25147, LUT_AMPL_WIDTH - 1),
		9126 => to_unsigned(25149, LUT_AMPL_WIDTH - 1),
		9127 => to_unsigned(25151, LUT_AMPL_WIDTH - 1),
		9128 => to_unsigned(25153, LUT_AMPL_WIDTH - 1),
		9129 => to_unsigned(25155, LUT_AMPL_WIDTH - 1),
		9130 => to_unsigned(25157, LUT_AMPL_WIDTH - 1),
		9131 => to_unsigned(25159, LUT_AMPL_WIDTH - 1),
		9132 => to_unsigned(25161, LUT_AMPL_WIDTH - 1),
		9133 => to_unsigned(25163, LUT_AMPL_WIDTH - 1),
		9134 => to_unsigned(25165, LUT_AMPL_WIDTH - 1),
		9135 => to_unsigned(25167, LUT_AMPL_WIDTH - 1),
		9136 => to_unsigned(25169, LUT_AMPL_WIDTH - 1),
		9137 => to_unsigned(25171, LUT_AMPL_WIDTH - 1),
		9138 => to_unsigned(25173, LUT_AMPL_WIDTH - 1),
		9139 => to_unsigned(25175, LUT_AMPL_WIDTH - 1),
		9140 => to_unsigned(25177, LUT_AMPL_WIDTH - 1),
		9141 => to_unsigned(25179, LUT_AMPL_WIDTH - 1),
		9142 => to_unsigned(25181, LUT_AMPL_WIDTH - 1),
		9143 => to_unsigned(25183, LUT_AMPL_WIDTH - 1),
		9144 => to_unsigned(25185, LUT_AMPL_WIDTH - 1),
		9145 => to_unsigned(25187, LUT_AMPL_WIDTH - 1),
		9146 => to_unsigned(25189, LUT_AMPL_WIDTH - 1),
		9147 => to_unsigned(25191, LUT_AMPL_WIDTH - 1),
		9148 => to_unsigned(25193, LUT_AMPL_WIDTH - 1),
		9149 => to_unsigned(25195, LUT_AMPL_WIDTH - 1),
		9150 => to_unsigned(25197, LUT_AMPL_WIDTH - 1),
		9151 => to_unsigned(25199, LUT_AMPL_WIDTH - 1),
		9152 => to_unsigned(25201, LUT_AMPL_WIDTH - 1),
		9153 => to_unsigned(25203, LUT_AMPL_WIDTH - 1),
		9154 => to_unsigned(25205, LUT_AMPL_WIDTH - 1),
		9155 => to_unsigned(25207, LUT_AMPL_WIDTH - 1),
		9156 => to_unsigned(25209, LUT_AMPL_WIDTH - 1),
		9157 => to_unsigned(25211, LUT_AMPL_WIDTH - 1),
		9158 => to_unsigned(25213, LUT_AMPL_WIDTH - 1),
		9159 => to_unsigned(25215, LUT_AMPL_WIDTH - 1),
		9160 => to_unsigned(25217, LUT_AMPL_WIDTH - 1),
		9161 => to_unsigned(25219, LUT_AMPL_WIDTH - 1),
		9162 => to_unsigned(25221, LUT_AMPL_WIDTH - 1),
		9163 => to_unsigned(25223, LUT_AMPL_WIDTH - 1),
		9164 => to_unsigned(25225, LUT_AMPL_WIDTH - 1),
		9165 => to_unsigned(25227, LUT_AMPL_WIDTH - 1),
		9166 => to_unsigned(25229, LUT_AMPL_WIDTH - 1),
		9167 => to_unsigned(25231, LUT_AMPL_WIDTH - 1),
		9168 => to_unsigned(25233, LUT_AMPL_WIDTH - 1),
		9169 => to_unsigned(25235, LUT_AMPL_WIDTH - 1),
		9170 => to_unsigned(25237, LUT_AMPL_WIDTH - 1),
		9171 => to_unsigned(25239, LUT_AMPL_WIDTH - 1),
		9172 => to_unsigned(25241, LUT_AMPL_WIDTH - 1),
		9173 => to_unsigned(25243, LUT_AMPL_WIDTH - 1),
		9174 => to_unsigned(25245, LUT_AMPL_WIDTH - 1),
		9175 => to_unsigned(25247, LUT_AMPL_WIDTH - 1),
		9176 => to_unsigned(25249, LUT_AMPL_WIDTH - 1),
		9177 => to_unsigned(25251, LUT_AMPL_WIDTH - 1),
		9178 => to_unsigned(25253, LUT_AMPL_WIDTH - 1),
		9179 => to_unsigned(25255, LUT_AMPL_WIDTH - 1),
		9180 => to_unsigned(25257, LUT_AMPL_WIDTH - 1),
		9181 => to_unsigned(25259, LUT_AMPL_WIDTH - 1),
		9182 => to_unsigned(25261, LUT_AMPL_WIDTH - 1),
		9183 => to_unsigned(25263, LUT_AMPL_WIDTH - 1),
		9184 => to_unsigned(25265, LUT_AMPL_WIDTH - 1),
		9185 => to_unsigned(25267, LUT_AMPL_WIDTH - 1),
		9186 => to_unsigned(25269, LUT_AMPL_WIDTH - 1),
		9187 => to_unsigned(25271, LUT_AMPL_WIDTH - 1),
		9188 => to_unsigned(25273, LUT_AMPL_WIDTH - 1),
		9189 => to_unsigned(25275, LUT_AMPL_WIDTH - 1),
		9190 => to_unsigned(25277, LUT_AMPL_WIDTH - 1),
		9191 => to_unsigned(25279, LUT_AMPL_WIDTH - 1),
		9192 => to_unsigned(25281, LUT_AMPL_WIDTH - 1),
		9193 => to_unsigned(25283, LUT_AMPL_WIDTH - 1),
		9194 => to_unsigned(25285, LUT_AMPL_WIDTH - 1),
		9195 => to_unsigned(25287, LUT_AMPL_WIDTH - 1),
		9196 => to_unsigned(25289, LUT_AMPL_WIDTH - 1),
		9197 => to_unsigned(25291, LUT_AMPL_WIDTH - 1),
		9198 => to_unsigned(25293, LUT_AMPL_WIDTH - 1),
		9199 => to_unsigned(25295, LUT_AMPL_WIDTH - 1),
		9200 => to_unsigned(25297, LUT_AMPL_WIDTH - 1),
		9201 => to_unsigned(25299, LUT_AMPL_WIDTH - 1),
		9202 => to_unsigned(25301, LUT_AMPL_WIDTH - 1),
		9203 => to_unsigned(25303, LUT_AMPL_WIDTH - 1),
		9204 => to_unsigned(25305, LUT_AMPL_WIDTH - 1),
		9205 => to_unsigned(25307, LUT_AMPL_WIDTH - 1),
		9206 => to_unsigned(25309, LUT_AMPL_WIDTH - 1),
		9207 => to_unsigned(25311, LUT_AMPL_WIDTH - 1),
		9208 => to_unsigned(25313, LUT_AMPL_WIDTH - 1),
		9209 => to_unsigned(25315, LUT_AMPL_WIDTH - 1),
		9210 => to_unsigned(25317, LUT_AMPL_WIDTH - 1),
		9211 => to_unsigned(25319, LUT_AMPL_WIDTH - 1),
		9212 => to_unsigned(25321, LUT_AMPL_WIDTH - 1),
		9213 => to_unsigned(25323, LUT_AMPL_WIDTH - 1),
		9214 => to_unsigned(25325, LUT_AMPL_WIDTH - 1),
		9215 => to_unsigned(25327, LUT_AMPL_WIDTH - 1),
		9216 => to_unsigned(25329, LUT_AMPL_WIDTH - 1),
		9217 => to_unsigned(25331, LUT_AMPL_WIDTH - 1),
		9218 => to_unsigned(25333, LUT_AMPL_WIDTH - 1),
		9219 => to_unsigned(25335, LUT_AMPL_WIDTH - 1),
		9220 => to_unsigned(25337, LUT_AMPL_WIDTH - 1),
		9221 => to_unsigned(25339, LUT_AMPL_WIDTH - 1),
		9222 => to_unsigned(25341, LUT_AMPL_WIDTH - 1),
		9223 => to_unsigned(25343, LUT_AMPL_WIDTH - 1),
		9224 => to_unsigned(25345, LUT_AMPL_WIDTH - 1),
		9225 => to_unsigned(25347, LUT_AMPL_WIDTH - 1),
		9226 => to_unsigned(25349, LUT_AMPL_WIDTH - 1),
		9227 => to_unsigned(25351, LUT_AMPL_WIDTH - 1),
		9228 => to_unsigned(25353, LUT_AMPL_WIDTH - 1),
		9229 => to_unsigned(25355, LUT_AMPL_WIDTH - 1),
		9230 => to_unsigned(25357, LUT_AMPL_WIDTH - 1),
		9231 => to_unsigned(25359, LUT_AMPL_WIDTH - 1),
		9232 => to_unsigned(25361, LUT_AMPL_WIDTH - 1),
		9233 => to_unsigned(25363, LUT_AMPL_WIDTH - 1),
		9234 => to_unsigned(25365, LUT_AMPL_WIDTH - 1),
		9235 => to_unsigned(25367, LUT_AMPL_WIDTH - 1),
		9236 => to_unsigned(25369, LUT_AMPL_WIDTH - 1),
		9237 => to_unsigned(25371, LUT_AMPL_WIDTH - 1),
		9238 => to_unsigned(25373, LUT_AMPL_WIDTH - 1),
		9239 => to_unsigned(25375, LUT_AMPL_WIDTH - 1),
		9240 => to_unsigned(25377, LUT_AMPL_WIDTH - 1),
		9241 => to_unsigned(25379, LUT_AMPL_WIDTH - 1),
		9242 => to_unsigned(25381, LUT_AMPL_WIDTH - 1),
		9243 => to_unsigned(25383, LUT_AMPL_WIDTH - 1),
		9244 => to_unsigned(25385, LUT_AMPL_WIDTH - 1),
		9245 => to_unsigned(25387, LUT_AMPL_WIDTH - 1),
		9246 => to_unsigned(25389, LUT_AMPL_WIDTH - 1),
		9247 => to_unsigned(25391, LUT_AMPL_WIDTH - 1),
		9248 => to_unsigned(25393, LUT_AMPL_WIDTH - 1),
		9249 => to_unsigned(25395, LUT_AMPL_WIDTH - 1),
		9250 => to_unsigned(25397, LUT_AMPL_WIDTH - 1),
		9251 => to_unsigned(25399, LUT_AMPL_WIDTH - 1),
		9252 => to_unsigned(25401, LUT_AMPL_WIDTH - 1),
		9253 => to_unsigned(25403, LUT_AMPL_WIDTH - 1),
		9254 => to_unsigned(25405, LUT_AMPL_WIDTH - 1),
		9255 => to_unsigned(25407, LUT_AMPL_WIDTH - 1),
		9256 => to_unsigned(25409, LUT_AMPL_WIDTH - 1),
		9257 => to_unsigned(25411, LUT_AMPL_WIDTH - 1),
		9258 => to_unsigned(25413, LUT_AMPL_WIDTH - 1),
		9259 => to_unsigned(25415, LUT_AMPL_WIDTH - 1),
		9260 => to_unsigned(25417, LUT_AMPL_WIDTH - 1),
		9261 => to_unsigned(25419, LUT_AMPL_WIDTH - 1),
		9262 => to_unsigned(25421, LUT_AMPL_WIDTH - 1),
		9263 => to_unsigned(25423, LUT_AMPL_WIDTH - 1),
		9264 => to_unsigned(25425, LUT_AMPL_WIDTH - 1),
		9265 => to_unsigned(25427, LUT_AMPL_WIDTH - 1),
		9266 => to_unsigned(25429, LUT_AMPL_WIDTH - 1),
		9267 => to_unsigned(25431, LUT_AMPL_WIDTH - 1),
		9268 => to_unsigned(25433, LUT_AMPL_WIDTH - 1),
		9269 => to_unsigned(25435, LUT_AMPL_WIDTH - 1),
		9270 => to_unsigned(25437, LUT_AMPL_WIDTH - 1),
		9271 => to_unsigned(25438, LUT_AMPL_WIDTH - 1),
		9272 => to_unsigned(25440, LUT_AMPL_WIDTH - 1),
		9273 => to_unsigned(25442, LUT_AMPL_WIDTH - 1),
		9274 => to_unsigned(25444, LUT_AMPL_WIDTH - 1),
		9275 => to_unsigned(25446, LUT_AMPL_WIDTH - 1),
		9276 => to_unsigned(25448, LUT_AMPL_WIDTH - 1),
		9277 => to_unsigned(25450, LUT_AMPL_WIDTH - 1),
		9278 => to_unsigned(25452, LUT_AMPL_WIDTH - 1),
		9279 => to_unsigned(25454, LUT_AMPL_WIDTH - 1),
		9280 => to_unsigned(25456, LUT_AMPL_WIDTH - 1),
		9281 => to_unsigned(25458, LUT_AMPL_WIDTH - 1),
		9282 => to_unsigned(25460, LUT_AMPL_WIDTH - 1),
		9283 => to_unsigned(25462, LUT_AMPL_WIDTH - 1),
		9284 => to_unsigned(25464, LUT_AMPL_WIDTH - 1),
		9285 => to_unsigned(25466, LUT_AMPL_WIDTH - 1),
		9286 => to_unsigned(25468, LUT_AMPL_WIDTH - 1),
		9287 => to_unsigned(25470, LUT_AMPL_WIDTH - 1),
		9288 => to_unsigned(25472, LUT_AMPL_WIDTH - 1),
		9289 => to_unsigned(25474, LUT_AMPL_WIDTH - 1),
		9290 => to_unsigned(25476, LUT_AMPL_WIDTH - 1),
		9291 => to_unsigned(25478, LUT_AMPL_WIDTH - 1),
		9292 => to_unsigned(25480, LUT_AMPL_WIDTH - 1),
		9293 => to_unsigned(25482, LUT_AMPL_WIDTH - 1),
		9294 => to_unsigned(25484, LUT_AMPL_WIDTH - 1),
		9295 => to_unsigned(25486, LUT_AMPL_WIDTH - 1),
		9296 => to_unsigned(25488, LUT_AMPL_WIDTH - 1),
		9297 => to_unsigned(25490, LUT_AMPL_WIDTH - 1),
		9298 => to_unsigned(25492, LUT_AMPL_WIDTH - 1),
		9299 => to_unsigned(25494, LUT_AMPL_WIDTH - 1),
		9300 => to_unsigned(25496, LUT_AMPL_WIDTH - 1),
		9301 => to_unsigned(25498, LUT_AMPL_WIDTH - 1),
		9302 => to_unsigned(25500, LUT_AMPL_WIDTH - 1),
		9303 => to_unsigned(25502, LUT_AMPL_WIDTH - 1),
		9304 => to_unsigned(25504, LUT_AMPL_WIDTH - 1),
		9305 => to_unsigned(25506, LUT_AMPL_WIDTH - 1),
		9306 => to_unsigned(25508, LUT_AMPL_WIDTH - 1),
		9307 => to_unsigned(25510, LUT_AMPL_WIDTH - 1),
		9308 => to_unsigned(25512, LUT_AMPL_WIDTH - 1),
		9309 => to_unsigned(25514, LUT_AMPL_WIDTH - 1),
		9310 => to_unsigned(25516, LUT_AMPL_WIDTH - 1),
		9311 => to_unsigned(25518, LUT_AMPL_WIDTH - 1),
		9312 => to_unsigned(25519, LUT_AMPL_WIDTH - 1),
		9313 => to_unsigned(25521, LUT_AMPL_WIDTH - 1),
		9314 => to_unsigned(25523, LUT_AMPL_WIDTH - 1),
		9315 => to_unsigned(25525, LUT_AMPL_WIDTH - 1),
		9316 => to_unsigned(25527, LUT_AMPL_WIDTH - 1),
		9317 => to_unsigned(25529, LUT_AMPL_WIDTH - 1),
		9318 => to_unsigned(25531, LUT_AMPL_WIDTH - 1),
		9319 => to_unsigned(25533, LUT_AMPL_WIDTH - 1),
		9320 => to_unsigned(25535, LUT_AMPL_WIDTH - 1),
		9321 => to_unsigned(25537, LUT_AMPL_WIDTH - 1),
		9322 => to_unsigned(25539, LUT_AMPL_WIDTH - 1),
		9323 => to_unsigned(25541, LUT_AMPL_WIDTH - 1),
		9324 => to_unsigned(25543, LUT_AMPL_WIDTH - 1),
		9325 => to_unsigned(25545, LUT_AMPL_WIDTH - 1),
		9326 => to_unsigned(25547, LUT_AMPL_WIDTH - 1),
		9327 => to_unsigned(25549, LUT_AMPL_WIDTH - 1),
		9328 => to_unsigned(25551, LUT_AMPL_WIDTH - 1),
		9329 => to_unsigned(25553, LUT_AMPL_WIDTH - 1),
		9330 => to_unsigned(25555, LUT_AMPL_WIDTH - 1),
		9331 => to_unsigned(25557, LUT_AMPL_WIDTH - 1),
		9332 => to_unsigned(25559, LUT_AMPL_WIDTH - 1),
		9333 => to_unsigned(25561, LUT_AMPL_WIDTH - 1),
		9334 => to_unsigned(25563, LUT_AMPL_WIDTH - 1),
		9335 => to_unsigned(25565, LUT_AMPL_WIDTH - 1),
		9336 => to_unsigned(25567, LUT_AMPL_WIDTH - 1),
		9337 => to_unsigned(25569, LUT_AMPL_WIDTH - 1),
		9338 => to_unsigned(25571, LUT_AMPL_WIDTH - 1),
		9339 => to_unsigned(25573, LUT_AMPL_WIDTH - 1),
		9340 => to_unsigned(25575, LUT_AMPL_WIDTH - 1),
		9341 => to_unsigned(25577, LUT_AMPL_WIDTH - 1),
		9342 => to_unsigned(25578, LUT_AMPL_WIDTH - 1),
		9343 => to_unsigned(25580, LUT_AMPL_WIDTH - 1),
		9344 => to_unsigned(25582, LUT_AMPL_WIDTH - 1),
		9345 => to_unsigned(25584, LUT_AMPL_WIDTH - 1),
		9346 => to_unsigned(25586, LUT_AMPL_WIDTH - 1),
		9347 => to_unsigned(25588, LUT_AMPL_WIDTH - 1),
		9348 => to_unsigned(25590, LUT_AMPL_WIDTH - 1),
		9349 => to_unsigned(25592, LUT_AMPL_WIDTH - 1),
		9350 => to_unsigned(25594, LUT_AMPL_WIDTH - 1),
		9351 => to_unsigned(25596, LUT_AMPL_WIDTH - 1),
		9352 => to_unsigned(25598, LUT_AMPL_WIDTH - 1),
		9353 => to_unsigned(25600, LUT_AMPL_WIDTH - 1),
		9354 => to_unsigned(25602, LUT_AMPL_WIDTH - 1),
		9355 => to_unsigned(25604, LUT_AMPL_WIDTH - 1),
		9356 => to_unsigned(25606, LUT_AMPL_WIDTH - 1),
		9357 => to_unsigned(25608, LUT_AMPL_WIDTH - 1),
		9358 => to_unsigned(25610, LUT_AMPL_WIDTH - 1),
		9359 => to_unsigned(25612, LUT_AMPL_WIDTH - 1),
		9360 => to_unsigned(25614, LUT_AMPL_WIDTH - 1),
		9361 => to_unsigned(25616, LUT_AMPL_WIDTH - 1),
		9362 => to_unsigned(25618, LUT_AMPL_WIDTH - 1),
		9363 => to_unsigned(25620, LUT_AMPL_WIDTH - 1),
		9364 => to_unsigned(25622, LUT_AMPL_WIDTH - 1),
		9365 => to_unsigned(25624, LUT_AMPL_WIDTH - 1),
		9366 => to_unsigned(25626, LUT_AMPL_WIDTH - 1),
		9367 => to_unsigned(25628, LUT_AMPL_WIDTH - 1),
		9368 => to_unsigned(25629, LUT_AMPL_WIDTH - 1),
		9369 => to_unsigned(25631, LUT_AMPL_WIDTH - 1),
		9370 => to_unsigned(25633, LUT_AMPL_WIDTH - 1),
		9371 => to_unsigned(25635, LUT_AMPL_WIDTH - 1),
		9372 => to_unsigned(25637, LUT_AMPL_WIDTH - 1),
		9373 => to_unsigned(25639, LUT_AMPL_WIDTH - 1),
		9374 => to_unsigned(25641, LUT_AMPL_WIDTH - 1),
		9375 => to_unsigned(25643, LUT_AMPL_WIDTH - 1),
		9376 => to_unsigned(25645, LUT_AMPL_WIDTH - 1),
		9377 => to_unsigned(25647, LUT_AMPL_WIDTH - 1),
		9378 => to_unsigned(25649, LUT_AMPL_WIDTH - 1),
		9379 => to_unsigned(25651, LUT_AMPL_WIDTH - 1),
		9380 => to_unsigned(25653, LUT_AMPL_WIDTH - 1),
		9381 => to_unsigned(25655, LUT_AMPL_WIDTH - 1),
		9382 => to_unsigned(25657, LUT_AMPL_WIDTH - 1),
		9383 => to_unsigned(25659, LUT_AMPL_WIDTH - 1),
		9384 => to_unsigned(25661, LUT_AMPL_WIDTH - 1),
		9385 => to_unsigned(25663, LUT_AMPL_WIDTH - 1),
		9386 => to_unsigned(25665, LUT_AMPL_WIDTH - 1),
		9387 => to_unsigned(25667, LUT_AMPL_WIDTH - 1),
		9388 => to_unsigned(25669, LUT_AMPL_WIDTH - 1),
		9389 => to_unsigned(25671, LUT_AMPL_WIDTH - 1),
		9390 => to_unsigned(25672, LUT_AMPL_WIDTH - 1),
		9391 => to_unsigned(25674, LUT_AMPL_WIDTH - 1),
		9392 => to_unsigned(25676, LUT_AMPL_WIDTH - 1),
		9393 => to_unsigned(25678, LUT_AMPL_WIDTH - 1),
		9394 => to_unsigned(25680, LUT_AMPL_WIDTH - 1),
		9395 => to_unsigned(25682, LUT_AMPL_WIDTH - 1),
		9396 => to_unsigned(25684, LUT_AMPL_WIDTH - 1),
		9397 => to_unsigned(25686, LUT_AMPL_WIDTH - 1),
		9398 => to_unsigned(25688, LUT_AMPL_WIDTH - 1),
		9399 => to_unsigned(25690, LUT_AMPL_WIDTH - 1),
		9400 => to_unsigned(25692, LUT_AMPL_WIDTH - 1),
		9401 => to_unsigned(25694, LUT_AMPL_WIDTH - 1),
		9402 => to_unsigned(25696, LUT_AMPL_WIDTH - 1),
		9403 => to_unsigned(25698, LUT_AMPL_WIDTH - 1),
		9404 => to_unsigned(25700, LUT_AMPL_WIDTH - 1),
		9405 => to_unsigned(25702, LUT_AMPL_WIDTH - 1),
		9406 => to_unsigned(25704, LUT_AMPL_WIDTH - 1),
		9407 => to_unsigned(25706, LUT_AMPL_WIDTH - 1),
		9408 => to_unsigned(25708, LUT_AMPL_WIDTH - 1),
		9409 => to_unsigned(25710, LUT_AMPL_WIDTH - 1),
		9410 => to_unsigned(25711, LUT_AMPL_WIDTH - 1),
		9411 => to_unsigned(25713, LUT_AMPL_WIDTH - 1),
		9412 => to_unsigned(25715, LUT_AMPL_WIDTH - 1),
		9413 => to_unsigned(25717, LUT_AMPL_WIDTH - 1),
		9414 => to_unsigned(25719, LUT_AMPL_WIDTH - 1),
		9415 => to_unsigned(25721, LUT_AMPL_WIDTH - 1),
		9416 => to_unsigned(25723, LUT_AMPL_WIDTH - 1),
		9417 => to_unsigned(25725, LUT_AMPL_WIDTH - 1),
		9418 => to_unsigned(25727, LUT_AMPL_WIDTH - 1),
		9419 => to_unsigned(25729, LUT_AMPL_WIDTH - 1),
		9420 => to_unsigned(25731, LUT_AMPL_WIDTH - 1),
		9421 => to_unsigned(25733, LUT_AMPL_WIDTH - 1),
		9422 => to_unsigned(25735, LUT_AMPL_WIDTH - 1),
		9423 => to_unsigned(25737, LUT_AMPL_WIDTH - 1),
		9424 => to_unsigned(25739, LUT_AMPL_WIDTH - 1),
		9425 => to_unsigned(25741, LUT_AMPL_WIDTH - 1),
		9426 => to_unsigned(25743, LUT_AMPL_WIDTH - 1),
		9427 => to_unsigned(25745, LUT_AMPL_WIDTH - 1),
		9428 => to_unsigned(25746, LUT_AMPL_WIDTH - 1),
		9429 => to_unsigned(25748, LUT_AMPL_WIDTH - 1),
		9430 => to_unsigned(25750, LUT_AMPL_WIDTH - 1),
		9431 => to_unsigned(25752, LUT_AMPL_WIDTH - 1),
		9432 => to_unsigned(25754, LUT_AMPL_WIDTH - 1),
		9433 => to_unsigned(25756, LUT_AMPL_WIDTH - 1),
		9434 => to_unsigned(25758, LUT_AMPL_WIDTH - 1),
		9435 => to_unsigned(25760, LUT_AMPL_WIDTH - 1),
		9436 => to_unsigned(25762, LUT_AMPL_WIDTH - 1),
		9437 => to_unsigned(25764, LUT_AMPL_WIDTH - 1),
		9438 => to_unsigned(25766, LUT_AMPL_WIDTH - 1),
		9439 => to_unsigned(25768, LUT_AMPL_WIDTH - 1),
		9440 => to_unsigned(25770, LUT_AMPL_WIDTH - 1),
		9441 => to_unsigned(25772, LUT_AMPL_WIDTH - 1),
		9442 => to_unsigned(25774, LUT_AMPL_WIDTH - 1),
		9443 => to_unsigned(25776, LUT_AMPL_WIDTH - 1),
		9444 => to_unsigned(25778, LUT_AMPL_WIDTH - 1),
		9445 => to_unsigned(25779, LUT_AMPL_WIDTH - 1),
		9446 => to_unsigned(25781, LUT_AMPL_WIDTH - 1),
		9447 => to_unsigned(25783, LUT_AMPL_WIDTH - 1),
		9448 => to_unsigned(25785, LUT_AMPL_WIDTH - 1),
		9449 => to_unsigned(25787, LUT_AMPL_WIDTH - 1),
		9450 => to_unsigned(25789, LUT_AMPL_WIDTH - 1),
		9451 => to_unsigned(25791, LUT_AMPL_WIDTH - 1),
		9452 => to_unsigned(25793, LUT_AMPL_WIDTH - 1),
		9453 => to_unsigned(25795, LUT_AMPL_WIDTH - 1),
		9454 => to_unsigned(25797, LUT_AMPL_WIDTH - 1),
		9455 => to_unsigned(25799, LUT_AMPL_WIDTH - 1),
		9456 => to_unsigned(25801, LUT_AMPL_WIDTH - 1),
		9457 => to_unsigned(25803, LUT_AMPL_WIDTH - 1),
		9458 => to_unsigned(25805, LUT_AMPL_WIDTH - 1),
		9459 => to_unsigned(25807, LUT_AMPL_WIDTH - 1),
		9460 => to_unsigned(25809, LUT_AMPL_WIDTH - 1),
		9461 => to_unsigned(25810, LUT_AMPL_WIDTH - 1),
		9462 => to_unsigned(25812, LUT_AMPL_WIDTH - 1),
		9463 => to_unsigned(25814, LUT_AMPL_WIDTH - 1),
		9464 => to_unsigned(25816, LUT_AMPL_WIDTH - 1),
		9465 => to_unsigned(25818, LUT_AMPL_WIDTH - 1),
		9466 => to_unsigned(25820, LUT_AMPL_WIDTH - 1),
		9467 => to_unsigned(25822, LUT_AMPL_WIDTH - 1),
		9468 => to_unsigned(25824, LUT_AMPL_WIDTH - 1),
		9469 => to_unsigned(25826, LUT_AMPL_WIDTH - 1),
		9470 => to_unsigned(25828, LUT_AMPL_WIDTH - 1),
		9471 => to_unsigned(25830, LUT_AMPL_WIDTH - 1),
		9472 => to_unsigned(25832, LUT_AMPL_WIDTH - 1),
		9473 => to_unsigned(25834, LUT_AMPL_WIDTH - 1),
		9474 => to_unsigned(25836, LUT_AMPL_WIDTH - 1),
		9475 => to_unsigned(25838, LUT_AMPL_WIDTH - 1),
		9476 => to_unsigned(25839, LUT_AMPL_WIDTH - 1),
		9477 => to_unsigned(25841, LUT_AMPL_WIDTH - 1),
		9478 => to_unsigned(25843, LUT_AMPL_WIDTH - 1),
		9479 => to_unsigned(25845, LUT_AMPL_WIDTH - 1),
		9480 => to_unsigned(25847, LUT_AMPL_WIDTH - 1),
		9481 => to_unsigned(25849, LUT_AMPL_WIDTH - 1),
		9482 => to_unsigned(25851, LUT_AMPL_WIDTH - 1),
		9483 => to_unsigned(25853, LUT_AMPL_WIDTH - 1),
		9484 => to_unsigned(25855, LUT_AMPL_WIDTH - 1),
		9485 => to_unsigned(25857, LUT_AMPL_WIDTH - 1),
		9486 => to_unsigned(25859, LUT_AMPL_WIDTH - 1),
		9487 => to_unsigned(25861, LUT_AMPL_WIDTH - 1),
		9488 => to_unsigned(25863, LUT_AMPL_WIDTH - 1),
		9489 => to_unsigned(25865, LUT_AMPL_WIDTH - 1),
		9490 => to_unsigned(25866, LUT_AMPL_WIDTH - 1),
		9491 => to_unsigned(25868, LUT_AMPL_WIDTH - 1),
		9492 => to_unsigned(25870, LUT_AMPL_WIDTH - 1),
		9493 => to_unsigned(25872, LUT_AMPL_WIDTH - 1),
		9494 => to_unsigned(25874, LUT_AMPL_WIDTH - 1),
		9495 => to_unsigned(25876, LUT_AMPL_WIDTH - 1),
		9496 => to_unsigned(25878, LUT_AMPL_WIDTH - 1),
		9497 => to_unsigned(25880, LUT_AMPL_WIDTH - 1),
		9498 => to_unsigned(25882, LUT_AMPL_WIDTH - 1),
		9499 => to_unsigned(25884, LUT_AMPL_WIDTH - 1),
		9500 => to_unsigned(25886, LUT_AMPL_WIDTH - 1),
		9501 => to_unsigned(25888, LUT_AMPL_WIDTH - 1),
		9502 => to_unsigned(25890, LUT_AMPL_WIDTH - 1),
		9503 => to_unsigned(25892, LUT_AMPL_WIDTH - 1),
		9504 => to_unsigned(25893, LUT_AMPL_WIDTH - 1),
		9505 => to_unsigned(25895, LUT_AMPL_WIDTH - 1),
		9506 => to_unsigned(25897, LUT_AMPL_WIDTH - 1),
		9507 => to_unsigned(25899, LUT_AMPL_WIDTH - 1),
		9508 => to_unsigned(25901, LUT_AMPL_WIDTH - 1),
		9509 => to_unsigned(25903, LUT_AMPL_WIDTH - 1),
		9510 => to_unsigned(25905, LUT_AMPL_WIDTH - 1),
		9511 => to_unsigned(25907, LUT_AMPL_WIDTH - 1),
		9512 => to_unsigned(25909, LUT_AMPL_WIDTH - 1),
		9513 => to_unsigned(25911, LUT_AMPL_WIDTH - 1),
		9514 => to_unsigned(25913, LUT_AMPL_WIDTH - 1),
		9515 => to_unsigned(25915, LUT_AMPL_WIDTH - 1),
		9516 => to_unsigned(25917, LUT_AMPL_WIDTH - 1),
		9517 => to_unsigned(25918, LUT_AMPL_WIDTH - 1),
		9518 => to_unsigned(25920, LUT_AMPL_WIDTH - 1),
		9519 => to_unsigned(25922, LUT_AMPL_WIDTH - 1),
		9520 => to_unsigned(25924, LUT_AMPL_WIDTH - 1),
		9521 => to_unsigned(25926, LUT_AMPL_WIDTH - 1),
		9522 => to_unsigned(25928, LUT_AMPL_WIDTH - 1),
		9523 => to_unsigned(25930, LUT_AMPL_WIDTH - 1),
		9524 => to_unsigned(25932, LUT_AMPL_WIDTH - 1),
		9525 => to_unsigned(25934, LUT_AMPL_WIDTH - 1),
		9526 => to_unsigned(25936, LUT_AMPL_WIDTH - 1),
		9527 => to_unsigned(25938, LUT_AMPL_WIDTH - 1),
		9528 => to_unsigned(25940, LUT_AMPL_WIDTH - 1),
		9529 => to_unsigned(25942, LUT_AMPL_WIDTH - 1),
		9530 => to_unsigned(25943, LUT_AMPL_WIDTH - 1),
		9531 => to_unsigned(25945, LUT_AMPL_WIDTH - 1),
		9532 => to_unsigned(25947, LUT_AMPL_WIDTH - 1),
		9533 => to_unsigned(25949, LUT_AMPL_WIDTH - 1),
		9534 => to_unsigned(25951, LUT_AMPL_WIDTH - 1),
		9535 => to_unsigned(25953, LUT_AMPL_WIDTH - 1),
		9536 => to_unsigned(25955, LUT_AMPL_WIDTH - 1),
		9537 => to_unsigned(25957, LUT_AMPL_WIDTH - 1),
		9538 => to_unsigned(25959, LUT_AMPL_WIDTH - 1),
		9539 => to_unsigned(25961, LUT_AMPL_WIDTH - 1),
		9540 => to_unsigned(25963, LUT_AMPL_WIDTH - 1),
		9541 => to_unsigned(25965, LUT_AMPL_WIDTH - 1),
		9542 => to_unsigned(25966, LUT_AMPL_WIDTH - 1),
		9543 => to_unsigned(25968, LUT_AMPL_WIDTH - 1),
		9544 => to_unsigned(25970, LUT_AMPL_WIDTH - 1),
		9545 => to_unsigned(25972, LUT_AMPL_WIDTH - 1),
		9546 => to_unsigned(25974, LUT_AMPL_WIDTH - 1),
		9547 => to_unsigned(25976, LUT_AMPL_WIDTH - 1),
		9548 => to_unsigned(25978, LUT_AMPL_WIDTH - 1),
		9549 => to_unsigned(25980, LUT_AMPL_WIDTH - 1),
		9550 => to_unsigned(25982, LUT_AMPL_WIDTH - 1),
		9551 => to_unsigned(25984, LUT_AMPL_WIDTH - 1),
		9552 => to_unsigned(25986, LUT_AMPL_WIDTH - 1),
		9553 => to_unsigned(25988, LUT_AMPL_WIDTH - 1),
		9554 => to_unsigned(25989, LUT_AMPL_WIDTH - 1),
		9555 => to_unsigned(25991, LUT_AMPL_WIDTH - 1),
		9556 => to_unsigned(25993, LUT_AMPL_WIDTH - 1),
		9557 => to_unsigned(25995, LUT_AMPL_WIDTH - 1),
		9558 => to_unsigned(25997, LUT_AMPL_WIDTH - 1),
		9559 => to_unsigned(25999, LUT_AMPL_WIDTH - 1),
		9560 => to_unsigned(26001, LUT_AMPL_WIDTH - 1),
		9561 => to_unsigned(26003, LUT_AMPL_WIDTH - 1),
		9562 => to_unsigned(26005, LUT_AMPL_WIDTH - 1),
		9563 => to_unsigned(26007, LUT_AMPL_WIDTH - 1),
		9564 => to_unsigned(26009, LUT_AMPL_WIDTH - 1),
		9565 => to_unsigned(26010, LUT_AMPL_WIDTH - 1),
		9566 => to_unsigned(26012, LUT_AMPL_WIDTH - 1),
		9567 => to_unsigned(26014, LUT_AMPL_WIDTH - 1),
		9568 => to_unsigned(26016, LUT_AMPL_WIDTH - 1),
		9569 => to_unsigned(26018, LUT_AMPL_WIDTH - 1),
		9570 => to_unsigned(26020, LUT_AMPL_WIDTH - 1),
		9571 => to_unsigned(26022, LUT_AMPL_WIDTH - 1),
		9572 => to_unsigned(26024, LUT_AMPL_WIDTH - 1),
		9573 => to_unsigned(26026, LUT_AMPL_WIDTH - 1),
		9574 => to_unsigned(26028, LUT_AMPL_WIDTH - 1),
		9575 => to_unsigned(26030, LUT_AMPL_WIDTH - 1),
		9576 => to_unsigned(26031, LUT_AMPL_WIDTH - 1),
		9577 => to_unsigned(26033, LUT_AMPL_WIDTH - 1),
		9578 => to_unsigned(26035, LUT_AMPL_WIDTH - 1),
		9579 => to_unsigned(26037, LUT_AMPL_WIDTH - 1),
		9580 => to_unsigned(26039, LUT_AMPL_WIDTH - 1),
		9581 => to_unsigned(26041, LUT_AMPL_WIDTH - 1),
		9582 => to_unsigned(26043, LUT_AMPL_WIDTH - 1),
		9583 => to_unsigned(26045, LUT_AMPL_WIDTH - 1),
		9584 => to_unsigned(26047, LUT_AMPL_WIDTH - 1),
		9585 => to_unsigned(26049, LUT_AMPL_WIDTH - 1),
		9586 => to_unsigned(26051, LUT_AMPL_WIDTH - 1),
		9587 => to_unsigned(26052, LUT_AMPL_WIDTH - 1),
		9588 => to_unsigned(26054, LUT_AMPL_WIDTH - 1),
		9589 => to_unsigned(26056, LUT_AMPL_WIDTH - 1),
		9590 => to_unsigned(26058, LUT_AMPL_WIDTH - 1),
		9591 => to_unsigned(26060, LUT_AMPL_WIDTH - 1),
		9592 => to_unsigned(26062, LUT_AMPL_WIDTH - 1),
		9593 => to_unsigned(26064, LUT_AMPL_WIDTH - 1),
		9594 => to_unsigned(26066, LUT_AMPL_WIDTH - 1),
		9595 => to_unsigned(26068, LUT_AMPL_WIDTH - 1),
		9596 => to_unsigned(26070, LUT_AMPL_WIDTH - 1),
		9597 => to_unsigned(26071, LUT_AMPL_WIDTH - 1),
		9598 => to_unsigned(26073, LUT_AMPL_WIDTH - 1),
		9599 => to_unsigned(26075, LUT_AMPL_WIDTH - 1),
		9600 => to_unsigned(26077, LUT_AMPL_WIDTH - 1),
		9601 => to_unsigned(26079, LUT_AMPL_WIDTH - 1),
		9602 => to_unsigned(26081, LUT_AMPL_WIDTH - 1),
		9603 => to_unsigned(26083, LUT_AMPL_WIDTH - 1),
		9604 => to_unsigned(26085, LUT_AMPL_WIDTH - 1),
		9605 => to_unsigned(26087, LUT_AMPL_WIDTH - 1),
		9606 => to_unsigned(26089, LUT_AMPL_WIDTH - 1),
		9607 => to_unsigned(26090, LUT_AMPL_WIDTH - 1),
		9608 => to_unsigned(26092, LUT_AMPL_WIDTH - 1),
		9609 => to_unsigned(26094, LUT_AMPL_WIDTH - 1),
		9610 => to_unsigned(26096, LUT_AMPL_WIDTH - 1),
		9611 => to_unsigned(26098, LUT_AMPL_WIDTH - 1),
		9612 => to_unsigned(26100, LUT_AMPL_WIDTH - 1),
		9613 => to_unsigned(26102, LUT_AMPL_WIDTH - 1),
		9614 => to_unsigned(26104, LUT_AMPL_WIDTH - 1),
		9615 => to_unsigned(26106, LUT_AMPL_WIDTH - 1),
		9616 => to_unsigned(26108, LUT_AMPL_WIDTH - 1),
		9617 => to_unsigned(26109, LUT_AMPL_WIDTH - 1),
		9618 => to_unsigned(26111, LUT_AMPL_WIDTH - 1),
		9619 => to_unsigned(26113, LUT_AMPL_WIDTH - 1),
		9620 => to_unsigned(26115, LUT_AMPL_WIDTH - 1),
		9621 => to_unsigned(26117, LUT_AMPL_WIDTH - 1),
		9622 => to_unsigned(26119, LUT_AMPL_WIDTH - 1),
		9623 => to_unsigned(26121, LUT_AMPL_WIDTH - 1),
		9624 => to_unsigned(26123, LUT_AMPL_WIDTH - 1),
		9625 => to_unsigned(26125, LUT_AMPL_WIDTH - 1),
		9626 => to_unsigned(26127, LUT_AMPL_WIDTH - 1),
		9627 => to_unsigned(26128, LUT_AMPL_WIDTH - 1),
		9628 => to_unsigned(26130, LUT_AMPL_WIDTH - 1),
		9629 => to_unsigned(26132, LUT_AMPL_WIDTH - 1),
		9630 => to_unsigned(26134, LUT_AMPL_WIDTH - 1),
		9631 => to_unsigned(26136, LUT_AMPL_WIDTH - 1),
		9632 => to_unsigned(26138, LUT_AMPL_WIDTH - 1),
		9633 => to_unsigned(26140, LUT_AMPL_WIDTH - 1),
		9634 => to_unsigned(26142, LUT_AMPL_WIDTH - 1),
		9635 => to_unsigned(26144, LUT_AMPL_WIDTH - 1),
		9636 => to_unsigned(26146, LUT_AMPL_WIDTH - 1),
		9637 => to_unsigned(26147, LUT_AMPL_WIDTH - 1),
		9638 => to_unsigned(26149, LUT_AMPL_WIDTH - 1),
		9639 => to_unsigned(26151, LUT_AMPL_WIDTH - 1),
		9640 => to_unsigned(26153, LUT_AMPL_WIDTH - 1),
		9641 => to_unsigned(26155, LUT_AMPL_WIDTH - 1),
		9642 => to_unsigned(26157, LUT_AMPL_WIDTH - 1),
		9643 => to_unsigned(26159, LUT_AMPL_WIDTH - 1),
		9644 => to_unsigned(26161, LUT_AMPL_WIDTH - 1),
		9645 => to_unsigned(26163, LUT_AMPL_WIDTH - 1),
		9646 => to_unsigned(26164, LUT_AMPL_WIDTH - 1),
		9647 => to_unsigned(26166, LUT_AMPL_WIDTH - 1),
		9648 => to_unsigned(26168, LUT_AMPL_WIDTH - 1),
		9649 => to_unsigned(26170, LUT_AMPL_WIDTH - 1),
		9650 => to_unsigned(26172, LUT_AMPL_WIDTH - 1),
		9651 => to_unsigned(26174, LUT_AMPL_WIDTH - 1),
		9652 => to_unsigned(26176, LUT_AMPL_WIDTH - 1),
		9653 => to_unsigned(26178, LUT_AMPL_WIDTH - 1),
		9654 => to_unsigned(26180, LUT_AMPL_WIDTH - 1),
		9655 => to_unsigned(26181, LUT_AMPL_WIDTH - 1),
		9656 => to_unsigned(26183, LUT_AMPL_WIDTH - 1),
		9657 => to_unsigned(26185, LUT_AMPL_WIDTH - 1),
		9658 => to_unsigned(26187, LUT_AMPL_WIDTH - 1),
		9659 => to_unsigned(26189, LUT_AMPL_WIDTH - 1),
		9660 => to_unsigned(26191, LUT_AMPL_WIDTH - 1),
		9661 => to_unsigned(26193, LUT_AMPL_WIDTH - 1),
		9662 => to_unsigned(26195, LUT_AMPL_WIDTH - 1),
		9663 => to_unsigned(26197, LUT_AMPL_WIDTH - 1),
		9664 => to_unsigned(26198, LUT_AMPL_WIDTH - 1),
		9665 => to_unsigned(26200, LUT_AMPL_WIDTH - 1),
		9666 => to_unsigned(26202, LUT_AMPL_WIDTH - 1),
		9667 => to_unsigned(26204, LUT_AMPL_WIDTH - 1),
		9668 => to_unsigned(26206, LUT_AMPL_WIDTH - 1),
		9669 => to_unsigned(26208, LUT_AMPL_WIDTH - 1),
		9670 => to_unsigned(26210, LUT_AMPL_WIDTH - 1),
		9671 => to_unsigned(26212, LUT_AMPL_WIDTH - 1),
		9672 => to_unsigned(26214, LUT_AMPL_WIDTH - 1),
		9673 => to_unsigned(26215, LUT_AMPL_WIDTH - 1),
		9674 => to_unsigned(26217, LUT_AMPL_WIDTH - 1),
		9675 => to_unsigned(26219, LUT_AMPL_WIDTH - 1),
		9676 => to_unsigned(26221, LUT_AMPL_WIDTH - 1),
		9677 => to_unsigned(26223, LUT_AMPL_WIDTH - 1),
		9678 => to_unsigned(26225, LUT_AMPL_WIDTH - 1),
		9679 => to_unsigned(26227, LUT_AMPL_WIDTH - 1),
		9680 => to_unsigned(26229, LUT_AMPL_WIDTH - 1),
		9681 => to_unsigned(26230, LUT_AMPL_WIDTH - 1),
		9682 => to_unsigned(26232, LUT_AMPL_WIDTH - 1),
		9683 => to_unsigned(26234, LUT_AMPL_WIDTH - 1),
		9684 => to_unsigned(26236, LUT_AMPL_WIDTH - 1),
		9685 => to_unsigned(26238, LUT_AMPL_WIDTH - 1),
		9686 => to_unsigned(26240, LUT_AMPL_WIDTH - 1),
		9687 => to_unsigned(26242, LUT_AMPL_WIDTH - 1),
		9688 => to_unsigned(26244, LUT_AMPL_WIDTH - 1),
		9689 => to_unsigned(26246, LUT_AMPL_WIDTH - 1),
		9690 => to_unsigned(26247, LUT_AMPL_WIDTH - 1),
		9691 => to_unsigned(26249, LUT_AMPL_WIDTH - 1),
		9692 => to_unsigned(26251, LUT_AMPL_WIDTH - 1),
		9693 => to_unsigned(26253, LUT_AMPL_WIDTH - 1),
		9694 => to_unsigned(26255, LUT_AMPL_WIDTH - 1),
		9695 => to_unsigned(26257, LUT_AMPL_WIDTH - 1),
		9696 => to_unsigned(26259, LUT_AMPL_WIDTH - 1),
		9697 => to_unsigned(26261, LUT_AMPL_WIDTH - 1),
		9698 => to_unsigned(26262, LUT_AMPL_WIDTH - 1),
		9699 => to_unsigned(26264, LUT_AMPL_WIDTH - 1),
		9700 => to_unsigned(26266, LUT_AMPL_WIDTH - 1),
		9701 => to_unsigned(26268, LUT_AMPL_WIDTH - 1),
		9702 => to_unsigned(26270, LUT_AMPL_WIDTH - 1),
		9703 => to_unsigned(26272, LUT_AMPL_WIDTH - 1),
		9704 => to_unsigned(26274, LUT_AMPL_WIDTH - 1),
		9705 => to_unsigned(26276, LUT_AMPL_WIDTH - 1),
		9706 => to_unsigned(26277, LUT_AMPL_WIDTH - 1),
		9707 => to_unsigned(26279, LUT_AMPL_WIDTH - 1),
		9708 => to_unsigned(26281, LUT_AMPL_WIDTH - 1),
		9709 => to_unsigned(26283, LUT_AMPL_WIDTH - 1),
		9710 => to_unsigned(26285, LUT_AMPL_WIDTH - 1),
		9711 => to_unsigned(26287, LUT_AMPL_WIDTH - 1),
		9712 => to_unsigned(26289, LUT_AMPL_WIDTH - 1),
		9713 => to_unsigned(26291, LUT_AMPL_WIDTH - 1),
		9714 => to_unsigned(26292, LUT_AMPL_WIDTH - 1),
		9715 => to_unsigned(26294, LUT_AMPL_WIDTH - 1),
		9716 => to_unsigned(26296, LUT_AMPL_WIDTH - 1),
		9717 => to_unsigned(26298, LUT_AMPL_WIDTH - 1),
		9718 => to_unsigned(26300, LUT_AMPL_WIDTH - 1),
		9719 => to_unsigned(26302, LUT_AMPL_WIDTH - 1),
		9720 => to_unsigned(26304, LUT_AMPL_WIDTH - 1),
		9721 => to_unsigned(26306, LUT_AMPL_WIDTH - 1),
		9722 => to_unsigned(26307, LUT_AMPL_WIDTH - 1),
		9723 => to_unsigned(26309, LUT_AMPL_WIDTH - 1),
		9724 => to_unsigned(26311, LUT_AMPL_WIDTH - 1),
		9725 => to_unsigned(26313, LUT_AMPL_WIDTH - 1),
		9726 => to_unsigned(26315, LUT_AMPL_WIDTH - 1),
		9727 => to_unsigned(26317, LUT_AMPL_WIDTH - 1),
		9728 => to_unsigned(26319, LUT_AMPL_WIDTH - 1),
		9729 => to_unsigned(26321, LUT_AMPL_WIDTH - 1),
		9730 => to_unsigned(26322, LUT_AMPL_WIDTH - 1),
		9731 => to_unsigned(26324, LUT_AMPL_WIDTH - 1),
		9732 => to_unsigned(26326, LUT_AMPL_WIDTH - 1),
		9733 => to_unsigned(26328, LUT_AMPL_WIDTH - 1),
		9734 => to_unsigned(26330, LUT_AMPL_WIDTH - 1),
		9735 => to_unsigned(26332, LUT_AMPL_WIDTH - 1),
		9736 => to_unsigned(26334, LUT_AMPL_WIDTH - 1),
		9737 => to_unsigned(26336, LUT_AMPL_WIDTH - 1),
		9738 => to_unsigned(26337, LUT_AMPL_WIDTH - 1),
		9739 => to_unsigned(26339, LUT_AMPL_WIDTH - 1),
		9740 => to_unsigned(26341, LUT_AMPL_WIDTH - 1),
		9741 => to_unsigned(26343, LUT_AMPL_WIDTH - 1),
		9742 => to_unsigned(26345, LUT_AMPL_WIDTH - 1),
		9743 => to_unsigned(26347, LUT_AMPL_WIDTH - 1),
		9744 => to_unsigned(26349, LUT_AMPL_WIDTH - 1),
		9745 => to_unsigned(26350, LUT_AMPL_WIDTH - 1),
		9746 => to_unsigned(26352, LUT_AMPL_WIDTH - 1),
		9747 => to_unsigned(26354, LUT_AMPL_WIDTH - 1),
		9748 => to_unsigned(26356, LUT_AMPL_WIDTH - 1),
		9749 => to_unsigned(26358, LUT_AMPL_WIDTH - 1),
		9750 => to_unsigned(26360, LUT_AMPL_WIDTH - 1),
		9751 => to_unsigned(26362, LUT_AMPL_WIDTH - 1),
		9752 => to_unsigned(26364, LUT_AMPL_WIDTH - 1),
		9753 => to_unsigned(26365, LUT_AMPL_WIDTH - 1),
		9754 => to_unsigned(26367, LUT_AMPL_WIDTH - 1),
		9755 => to_unsigned(26369, LUT_AMPL_WIDTH - 1),
		9756 => to_unsigned(26371, LUT_AMPL_WIDTH - 1),
		9757 => to_unsigned(26373, LUT_AMPL_WIDTH - 1),
		9758 => to_unsigned(26375, LUT_AMPL_WIDTH - 1),
		9759 => to_unsigned(26377, LUT_AMPL_WIDTH - 1),
		9760 => to_unsigned(26378, LUT_AMPL_WIDTH - 1),
		9761 => to_unsigned(26380, LUT_AMPL_WIDTH - 1),
		9762 => to_unsigned(26382, LUT_AMPL_WIDTH - 1),
		9763 => to_unsigned(26384, LUT_AMPL_WIDTH - 1),
		9764 => to_unsigned(26386, LUT_AMPL_WIDTH - 1),
		9765 => to_unsigned(26388, LUT_AMPL_WIDTH - 1),
		9766 => to_unsigned(26390, LUT_AMPL_WIDTH - 1),
		9767 => to_unsigned(26392, LUT_AMPL_WIDTH - 1),
		9768 => to_unsigned(26393, LUT_AMPL_WIDTH - 1),
		9769 => to_unsigned(26395, LUT_AMPL_WIDTH - 1),
		9770 => to_unsigned(26397, LUT_AMPL_WIDTH - 1),
		9771 => to_unsigned(26399, LUT_AMPL_WIDTH - 1),
		9772 => to_unsigned(26401, LUT_AMPL_WIDTH - 1),
		9773 => to_unsigned(26403, LUT_AMPL_WIDTH - 1),
		9774 => to_unsigned(26405, LUT_AMPL_WIDTH - 1),
		9775 => to_unsigned(26406, LUT_AMPL_WIDTH - 1),
		9776 => to_unsigned(26408, LUT_AMPL_WIDTH - 1),
		9777 => to_unsigned(26410, LUT_AMPL_WIDTH - 1),
		9778 => to_unsigned(26412, LUT_AMPL_WIDTH - 1),
		9779 => to_unsigned(26414, LUT_AMPL_WIDTH - 1),
		9780 => to_unsigned(26416, LUT_AMPL_WIDTH - 1),
		9781 => to_unsigned(26418, LUT_AMPL_WIDTH - 1),
		9782 => to_unsigned(26419, LUT_AMPL_WIDTH - 1),
		9783 => to_unsigned(26421, LUT_AMPL_WIDTH - 1),
		9784 => to_unsigned(26423, LUT_AMPL_WIDTH - 1),
		9785 => to_unsigned(26425, LUT_AMPL_WIDTH - 1),
		9786 => to_unsigned(26427, LUT_AMPL_WIDTH - 1),
		9787 => to_unsigned(26429, LUT_AMPL_WIDTH - 1),
		9788 => to_unsigned(26431, LUT_AMPL_WIDTH - 1),
		9789 => to_unsigned(26432, LUT_AMPL_WIDTH - 1),
		9790 => to_unsigned(26434, LUT_AMPL_WIDTH - 1),
		9791 => to_unsigned(26436, LUT_AMPL_WIDTH - 1),
		9792 => to_unsigned(26438, LUT_AMPL_WIDTH - 1),
		9793 => to_unsigned(26440, LUT_AMPL_WIDTH - 1),
		9794 => to_unsigned(26442, LUT_AMPL_WIDTH - 1),
		9795 => to_unsigned(26444, LUT_AMPL_WIDTH - 1),
		9796 => to_unsigned(26445, LUT_AMPL_WIDTH - 1),
		9797 => to_unsigned(26447, LUT_AMPL_WIDTH - 1),
		9798 => to_unsigned(26449, LUT_AMPL_WIDTH - 1),
		9799 => to_unsigned(26451, LUT_AMPL_WIDTH - 1),
		9800 => to_unsigned(26453, LUT_AMPL_WIDTH - 1),
		9801 => to_unsigned(26455, LUT_AMPL_WIDTH - 1),
		9802 => to_unsigned(26457, LUT_AMPL_WIDTH - 1),
		9803 => to_unsigned(26458, LUT_AMPL_WIDTH - 1),
		9804 => to_unsigned(26460, LUT_AMPL_WIDTH - 1),
		9805 => to_unsigned(26462, LUT_AMPL_WIDTH - 1),
		9806 => to_unsigned(26464, LUT_AMPL_WIDTH - 1),
		9807 => to_unsigned(26466, LUT_AMPL_WIDTH - 1),
		9808 => to_unsigned(26468, LUT_AMPL_WIDTH - 1),
		9809 => to_unsigned(26469, LUT_AMPL_WIDTH - 1),
		9810 => to_unsigned(26471, LUT_AMPL_WIDTH - 1),
		9811 => to_unsigned(26473, LUT_AMPL_WIDTH - 1),
		9812 => to_unsigned(26475, LUT_AMPL_WIDTH - 1),
		9813 => to_unsigned(26477, LUT_AMPL_WIDTH - 1),
		9814 => to_unsigned(26479, LUT_AMPL_WIDTH - 1),
		9815 => to_unsigned(26481, LUT_AMPL_WIDTH - 1),
		9816 => to_unsigned(26482, LUT_AMPL_WIDTH - 1),
		9817 => to_unsigned(26484, LUT_AMPL_WIDTH - 1),
		9818 => to_unsigned(26486, LUT_AMPL_WIDTH - 1),
		9819 => to_unsigned(26488, LUT_AMPL_WIDTH - 1),
		9820 => to_unsigned(26490, LUT_AMPL_WIDTH - 1),
		9821 => to_unsigned(26492, LUT_AMPL_WIDTH - 1),
		9822 => to_unsigned(26494, LUT_AMPL_WIDTH - 1),
		9823 => to_unsigned(26495, LUT_AMPL_WIDTH - 1),
		9824 => to_unsigned(26497, LUT_AMPL_WIDTH - 1),
		9825 => to_unsigned(26499, LUT_AMPL_WIDTH - 1),
		9826 => to_unsigned(26501, LUT_AMPL_WIDTH - 1),
		9827 => to_unsigned(26503, LUT_AMPL_WIDTH - 1),
		9828 => to_unsigned(26505, LUT_AMPL_WIDTH - 1),
		9829 => to_unsigned(26506, LUT_AMPL_WIDTH - 1),
		9830 => to_unsigned(26508, LUT_AMPL_WIDTH - 1),
		9831 => to_unsigned(26510, LUT_AMPL_WIDTH - 1),
		9832 => to_unsigned(26512, LUT_AMPL_WIDTH - 1),
		9833 => to_unsigned(26514, LUT_AMPL_WIDTH - 1),
		9834 => to_unsigned(26516, LUT_AMPL_WIDTH - 1),
		9835 => to_unsigned(26518, LUT_AMPL_WIDTH - 1),
		9836 => to_unsigned(26519, LUT_AMPL_WIDTH - 1),
		9837 => to_unsigned(26521, LUT_AMPL_WIDTH - 1),
		9838 => to_unsigned(26523, LUT_AMPL_WIDTH - 1),
		9839 => to_unsigned(26525, LUT_AMPL_WIDTH - 1),
		9840 => to_unsigned(26527, LUT_AMPL_WIDTH - 1),
		9841 => to_unsigned(26529, LUT_AMPL_WIDTH - 1),
		9842 => to_unsigned(26530, LUT_AMPL_WIDTH - 1),
		9843 => to_unsigned(26532, LUT_AMPL_WIDTH - 1),
		9844 => to_unsigned(26534, LUT_AMPL_WIDTH - 1),
		9845 => to_unsigned(26536, LUT_AMPL_WIDTH - 1),
		9846 => to_unsigned(26538, LUT_AMPL_WIDTH - 1),
		9847 => to_unsigned(26540, LUT_AMPL_WIDTH - 1),
		9848 => to_unsigned(26542, LUT_AMPL_WIDTH - 1),
		9849 => to_unsigned(26543, LUT_AMPL_WIDTH - 1),
		9850 => to_unsigned(26545, LUT_AMPL_WIDTH - 1),
		9851 => to_unsigned(26547, LUT_AMPL_WIDTH - 1),
		9852 => to_unsigned(26549, LUT_AMPL_WIDTH - 1),
		9853 => to_unsigned(26551, LUT_AMPL_WIDTH - 1),
		9854 => to_unsigned(26553, LUT_AMPL_WIDTH - 1),
		9855 => to_unsigned(26554, LUT_AMPL_WIDTH - 1),
		9856 => to_unsigned(26556, LUT_AMPL_WIDTH - 1),
		9857 => to_unsigned(26558, LUT_AMPL_WIDTH - 1),
		9858 => to_unsigned(26560, LUT_AMPL_WIDTH - 1),
		9859 => to_unsigned(26562, LUT_AMPL_WIDTH - 1),
		9860 => to_unsigned(26564, LUT_AMPL_WIDTH - 1),
		9861 => to_unsigned(26565, LUT_AMPL_WIDTH - 1),
		9862 => to_unsigned(26567, LUT_AMPL_WIDTH - 1),
		9863 => to_unsigned(26569, LUT_AMPL_WIDTH - 1),
		9864 => to_unsigned(26571, LUT_AMPL_WIDTH - 1),
		9865 => to_unsigned(26573, LUT_AMPL_WIDTH - 1),
		9866 => to_unsigned(26575, LUT_AMPL_WIDTH - 1),
		9867 => to_unsigned(26576, LUT_AMPL_WIDTH - 1),
		9868 => to_unsigned(26578, LUT_AMPL_WIDTH - 1),
		9869 => to_unsigned(26580, LUT_AMPL_WIDTH - 1),
		9870 => to_unsigned(26582, LUT_AMPL_WIDTH - 1),
		9871 => to_unsigned(26584, LUT_AMPL_WIDTH - 1),
		9872 => to_unsigned(26586, LUT_AMPL_WIDTH - 1),
		9873 => to_unsigned(26588, LUT_AMPL_WIDTH - 1),
		9874 => to_unsigned(26589, LUT_AMPL_WIDTH - 1),
		9875 => to_unsigned(26591, LUT_AMPL_WIDTH - 1),
		9876 => to_unsigned(26593, LUT_AMPL_WIDTH - 1),
		9877 => to_unsigned(26595, LUT_AMPL_WIDTH - 1),
		9878 => to_unsigned(26597, LUT_AMPL_WIDTH - 1),
		9879 => to_unsigned(26599, LUT_AMPL_WIDTH - 1),
		9880 => to_unsigned(26600, LUT_AMPL_WIDTH - 1),
		9881 => to_unsigned(26602, LUT_AMPL_WIDTH - 1),
		9882 => to_unsigned(26604, LUT_AMPL_WIDTH - 1),
		9883 => to_unsigned(26606, LUT_AMPL_WIDTH - 1),
		9884 => to_unsigned(26608, LUT_AMPL_WIDTH - 1),
		9885 => to_unsigned(26610, LUT_AMPL_WIDTH - 1),
		9886 => to_unsigned(26611, LUT_AMPL_WIDTH - 1),
		9887 => to_unsigned(26613, LUT_AMPL_WIDTH - 1),
		9888 => to_unsigned(26615, LUT_AMPL_WIDTH - 1),
		9889 => to_unsigned(26617, LUT_AMPL_WIDTH - 1),
		9890 => to_unsigned(26619, LUT_AMPL_WIDTH - 1),
		9891 => to_unsigned(26621, LUT_AMPL_WIDTH - 1),
		9892 => to_unsigned(26622, LUT_AMPL_WIDTH - 1),
		9893 => to_unsigned(26624, LUT_AMPL_WIDTH - 1),
		9894 => to_unsigned(26626, LUT_AMPL_WIDTH - 1),
		9895 => to_unsigned(26628, LUT_AMPL_WIDTH - 1),
		9896 => to_unsigned(26630, LUT_AMPL_WIDTH - 1),
		9897 => to_unsigned(26631, LUT_AMPL_WIDTH - 1),
		9898 => to_unsigned(26633, LUT_AMPL_WIDTH - 1),
		9899 => to_unsigned(26635, LUT_AMPL_WIDTH - 1),
		9900 => to_unsigned(26637, LUT_AMPL_WIDTH - 1),
		9901 => to_unsigned(26639, LUT_AMPL_WIDTH - 1),
		9902 => to_unsigned(26641, LUT_AMPL_WIDTH - 1),
		9903 => to_unsigned(26642, LUT_AMPL_WIDTH - 1),
		9904 => to_unsigned(26644, LUT_AMPL_WIDTH - 1),
		9905 => to_unsigned(26646, LUT_AMPL_WIDTH - 1),
		9906 => to_unsigned(26648, LUT_AMPL_WIDTH - 1),
		9907 => to_unsigned(26650, LUT_AMPL_WIDTH - 1),
		9908 => to_unsigned(26652, LUT_AMPL_WIDTH - 1),
		9909 => to_unsigned(26653, LUT_AMPL_WIDTH - 1),
		9910 => to_unsigned(26655, LUT_AMPL_WIDTH - 1),
		9911 => to_unsigned(26657, LUT_AMPL_WIDTH - 1),
		9912 => to_unsigned(26659, LUT_AMPL_WIDTH - 1),
		9913 => to_unsigned(26661, LUT_AMPL_WIDTH - 1),
		9914 => to_unsigned(26663, LUT_AMPL_WIDTH - 1),
		9915 => to_unsigned(26664, LUT_AMPL_WIDTH - 1),
		9916 => to_unsigned(26666, LUT_AMPL_WIDTH - 1),
		9917 => to_unsigned(26668, LUT_AMPL_WIDTH - 1),
		9918 => to_unsigned(26670, LUT_AMPL_WIDTH - 1),
		9919 => to_unsigned(26672, LUT_AMPL_WIDTH - 1),
		9920 => to_unsigned(26674, LUT_AMPL_WIDTH - 1),
		9921 => to_unsigned(26675, LUT_AMPL_WIDTH - 1),
		9922 => to_unsigned(26677, LUT_AMPL_WIDTH - 1),
		9923 => to_unsigned(26679, LUT_AMPL_WIDTH - 1),
		9924 => to_unsigned(26681, LUT_AMPL_WIDTH - 1),
		9925 => to_unsigned(26683, LUT_AMPL_WIDTH - 1),
		9926 => to_unsigned(26684, LUT_AMPL_WIDTH - 1),
		9927 => to_unsigned(26686, LUT_AMPL_WIDTH - 1),
		9928 => to_unsigned(26688, LUT_AMPL_WIDTH - 1),
		9929 => to_unsigned(26690, LUT_AMPL_WIDTH - 1),
		9930 => to_unsigned(26692, LUT_AMPL_WIDTH - 1),
		9931 => to_unsigned(26694, LUT_AMPL_WIDTH - 1),
		9932 => to_unsigned(26695, LUT_AMPL_WIDTH - 1),
		9933 => to_unsigned(26697, LUT_AMPL_WIDTH - 1),
		9934 => to_unsigned(26699, LUT_AMPL_WIDTH - 1),
		9935 => to_unsigned(26701, LUT_AMPL_WIDTH - 1),
		9936 => to_unsigned(26703, LUT_AMPL_WIDTH - 1),
		9937 => to_unsigned(26705, LUT_AMPL_WIDTH - 1),
		9938 => to_unsigned(26706, LUT_AMPL_WIDTH - 1),
		9939 => to_unsigned(26708, LUT_AMPL_WIDTH - 1),
		9940 => to_unsigned(26710, LUT_AMPL_WIDTH - 1),
		9941 => to_unsigned(26712, LUT_AMPL_WIDTH - 1),
		9942 => to_unsigned(26714, LUT_AMPL_WIDTH - 1),
		9943 => to_unsigned(26715, LUT_AMPL_WIDTH - 1),
		9944 => to_unsigned(26717, LUT_AMPL_WIDTH - 1),
		9945 => to_unsigned(26719, LUT_AMPL_WIDTH - 1),
		9946 => to_unsigned(26721, LUT_AMPL_WIDTH - 1),
		9947 => to_unsigned(26723, LUT_AMPL_WIDTH - 1),
		9948 => to_unsigned(26725, LUT_AMPL_WIDTH - 1),
		9949 => to_unsigned(26726, LUT_AMPL_WIDTH - 1),
		9950 => to_unsigned(26728, LUT_AMPL_WIDTH - 1),
		9951 => to_unsigned(26730, LUT_AMPL_WIDTH - 1),
		9952 => to_unsigned(26732, LUT_AMPL_WIDTH - 1),
		9953 => to_unsigned(26734, LUT_AMPL_WIDTH - 1),
		9954 => to_unsigned(26735, LUT_AMPL_WIDTH - 1),
		9955 => to_unsigned(26737, LUT_AMPL_WIDTH - 1),
		9956 => to_unsigned(26739, LUT_AMPL_WIDTH - 1),
		9957 => to_unsigned(26741, LUT_AMPL_WIDTH - 1),
		9958 => to_unsigned(26743, LUT_AMPL_WIDTH - 1),
		9959 => to_unsigned(26745, LUT_AMPL_WIDTH - 1),
		9960 => to_unsigned(26746, LUT_AMPL_WIDTH - 1),
		9961 => to_unsigned(26748, LUT_AMPL_WIDTH - 1),
		9962 => to_unsigned(26750, LUT_AMPL_WIDTH - 1),
		9963 => to_unsigned(26752, LUT_AMPL_WIDTH - 1),
		9964 => to_unsigned(26754, LUT_AMPL_WIDTH - 1),
		9965 => to_unsigned(26755, LUT_AMPL_WIDTH - 1),
		9966 => to_unsigned(26757, LUT_AMPL_WIDTH - 1),
		9967 => to_unsigned(26759, LUT_AMPL_WIDTH - 1),
		9968 => to_unsigned(26761, LUT_AMPL_WIDTH - 1),
		9969 => to_unsigned(26763, LUT_AMPL_WIDTH - 1),
		9970 => to_unsigned(26764, LUT_AMPL_WIDTH - 1),
		9971 => to_unsigned(26766, LUT_AMPL_WIDTH - 1),
		9972 => to_unsigned(26768, LUT_AMPL_WIDTH - 1),
		9973 => to_unsigned(26770, LUT_AMPL_WIDTH - 1),
		9974 => to_unsigned(26772, LUT_AMPL_WIDTH - 1),
		9975 => to_unsigned(26774, LUT_AMPL_WIDTH - 1),
		9976 => to_unsigned(26775, LUT_AMPL_WIDTH - 1),
		9977 => to_unsigned(26777, LUT_AMPL_WIDTH - 1),
		9978 => to_unsigned(26779, LUT_AMPL_WIDTH - 1),
		9979 => to_unsigned(26781, LUT_AMPL_WIDTH - 1),
		9980 => to_unsigned(26783, LUT_AMPL_WIDTH - 1),
		9981 => to_unsigned(26784, LUT_AMPL_WIDTH - 1),
		9982 => to_unsigned(26786, LUT_AMPL_WIDTH - 1),
		9983 => to_unsigned(26788, LUT_AMPL_WIDTH - 1),
		9984 => to_unsigned(26790, LUT_AMPL_WIDTH - 1),
		9985 => to_unsigned(26792, LUT_AMPL_WIDTH - 1),
		9986 => to_unsigned(26793, LUT_AMPL_WIDTH - 1),
		9987 => to_unsigned(26795, LUT_AMPL_WIDTH - 1),
		9988 => to_unsigned(26797, LUT_AMPL_WIDTH - 1),
		9989 => to_unsigned(26799, LUT_AMPL_WIDTH - 1),
		9990 => to_unsigned(26801, LUT_AMPL_WIDTH - 1),
		9991 => to_unsigned(26802, LUT_AMPL_WIDTH - 1),
		9992 => to_unsigned(26804, LUT_AMPL_WIDTH - 1),
		9993 => to_unsigned(26806, LUT_AMPL_WIDTH - 1),
		9994 => to_unsigned(26808, LUT_AMPL_WIDTH - 1),
		9995 => to_unsigned(26810, LUT_AMPL_WIDTH - 1),
		9996 => to_unsigned(26811, LUT_AMPL_WIDTH - 1),
		9997 => to_unsigned(26813, LUT_AMPL_WIDTH - 1),
		9998 => to_unsigned(26815, LUT_AMPL_WIDTH - 1),
		9999 => to_unsigned(26817, LUT_AMPL_WIDTH - 1),
		10000 => to_unsigned(26819, LUT_AMPL_WIDTH - 1),
		10001 => to_unsigned(26821, LUT_AMPL_WIDTH - 1),
		10002 => to_unsigned(26822, LUT_AMPL_WIDTH - 1),
		10003 => to_unsigned(26824, LUT_AMPL_WIDTH - 1),
		10004 => to_unsigned(26826, LUT_AMPL_WIDTH - 1),
		10005 => to_unsigned(26828, LUT_AMPL_WIDTH - 1),
		10006 => to_unsigned(26830, LUT_AMPL_WIDTH - 1),
		10007 => to_unsigned(26831, LUT_AMPL_WIDTH - 1),
		10008 => to_unsigned(26833, LUT_AMPL_WIDTH - 1),
		10009 => to_unsigned(26835, LUT_AMPL_WIDTH - 1),
		10010 => to_unsigned(26837, LUT_AMPL_WIDTH - 1),
		10011 => to_unsigned(26839, LUT_AMPL_WIDTH - 1),
		10012 => to_unsigned(26840, LUT_AMPL_WIDTH - 1),
		10013 => to_unsigned(26842, LUT_AMPL_WIDTH - 1),
		10014 => to_unsigned(26844, LUT_AMPL_WIDTH - 1),
		10015 => to_unsigned(26846, LUT_AMPL_WIDTH - 1),
		10016 => to_unsigned(26848, LUT_AMPL_WIDTH - 1),
		10017 => to_unsigned(26849, LUT_AMPL_WIDTH - 1),
		10018 => to_unsigned(26851, LUT_AMPL_WIDTH - 1),
		10019 => to_unsigned(26853, LUT_AMPL_WIDTH - 1),
		10020 => to_unsigned(26855, LUT_AMPL_WIDTH - 1),
		10021 => to_unsigned(26857, LUT_AMPL_WIDTH - 1),
		10022 => to_unsigned(26858, LUT_AMPL_WIDTH - 1),
		10023 => to_unsigned(26860, LUT_AMPL_WIDTH - 1),
		10024 => to_unsigned(26862, LUT_AMPL_WIDTH - 1),
		10025 => to_unsigned(26864, LUT_AMPL_WIDTH - 1),
		10026 => to_unsigned(26866, LUT_AMPL_WIDTH - 1),
		10027 => to_unsigned(26867, LUT_AMPL_WIDTH - 1),
		10028 => to_unsigned(26869, LUT_AMPL_WIDTH - 1),
		10029 => to_unsigned(26871, LUT_AMPL_WIDTH - 1),
		10030 => to_unsigned(26873, LUT_AMPL_WIDTH - 1),
		10031 => to_unsigned(26875, LUT_AMPL_WIDTH - 1),
		10032 => to_unsigned(26876, LUT_AMPL_WIDTH - 1),
		10033 => to_unsigned(26878, LUT_AMPL_WIDTH - 1),
		10034 => to_unsigned(26880, LUT_AMPL_WIDTH - 1),
		10035 => to_unsigned(26882, LUT_AMPL_WIDTH - 1),
		10036 => to_unsigned(26884, LUT_AMPL_WIDTH - 1),
		10037 => to_unsigned(26885, LUT_AMPL_WIDTH - 1),
		10038 => to_unsigned(26887, LUT_AMPL_WIDTH - 1),
		10039 => to_unsigned(26889, LUT_AMPL_WIDTH - 1),
		10040 => to_unsigned(26891, LUT_AMPL_WIDTH - 1),
		10041 => to_unsigned(26893, LUT_AMPL_WIDTH - 1),
		10042 => to_unsigned(26894, LUT_AMPL_WIDTH - 1),
		10043 => to_unsigned(26896, LUT_AMPL_WIDTH - 1),
		10044 => to_unsigned(26898, LUT_AMPL_WIDTH - 1),
		10045 => to_unsigned(26900, LUT_AMPL_WIDTH - 1),
		10046 => to_unsigned(26901, LUT_AMPL_WIDTH - 1),
		10047 => to_unsigned(26903, LUT_AMPL_WIDTH - 1),
		10048 => to_unsigned(26905, LUT_AMPL_WIDTH - 1),
		10049 => to_unsigned(26907, LUT_AMPL_WIDTH - 1),
		10050 => to_unsigned(26909, LUT_AMPL_WIDTH - 1),
		10051 => to_unsigned(26910, LUT_AMPL_WIDTH - 1),
		10052 => to_unsigned(26912, LUT_AMPL_WIDTH - 1),
		10053 => to_unsigned(26914, LUT_AMPL_WIDTH - 1),
		10054 => to_unsigned(26916, LUT_AMPL_WIDTH - 1),
		10055 => to_unsigned(26918, LUT_AMPL_WIDTH - 1),
		10056 => to_unsigned(26919, LUT_AMPL_WIDTH - 1),
		10057 => to_unsigned(26921, LUT_AMPL_WIDTH - 1),
		10058 => to_unsigned(26923, LUT_AMPL_WIDTH - 1),
		10059 => to_unsigned(26925, LUT_AMPL_WIDTH - 1),
		10060 => to_unsigned(26927, LUT_AMPL_WIDTH - 1),
		10061 => to_unsigned(26928, LUT_AMPL_WIDTH - 1),
		10062 => to_unsigned(26930, LUT_AMPL_WIDTH - 1),
		10063 => to_unsigned(26932, LUT_AMPL_WIDTH - 1),
		10064 => to_unsigned(26934, LUT_AMPL_WIDTH - 1),
		10065 => to_unsigned(26936, LUT_AMPL_WIDTH - 1),
		10066 => to_unsigned(26937, LUT_AMPL_WIDTH - 1),
		10067 => to_unsigned(26939, LUT_AMPL_WIDTH - 1),
		10068 => to_unsigned(26941, LUT_AMPL_WIDTH - 1),
		10069 => to_unsigned(26943, LUT_AMPL_WIDTH - 1),
		10070 => to_unsigned(26944, LUT_AMPL_WIDTH - 1),
		10071 => to_unsigned(26946, LUT_AMPL_WIDTH - 1),
		10072 => to_unsigned(26948, LUT_AMPL_WIDTH - 1),
		10073 => to_unsigned(26950, LUT_AMPL_WIDTH - 1),
		10074 => to_unsigned(26952, LUT_AMPL_WIDTH - 1),
		10075 => to_unsigned(26953, LUT_AMPL_WIDTH - 1),
		10076 => to_unsigned(26955, LUT_AMPL_WIDTH - 1),
		10077 => to_unsigned(26957, LUT_AMPL_WIDTH - 1),
		10078 => to_unsigned(26959, LUT_AMPL_WIDTH - 1),
		10079 => to_unsigned(26961, LUT_AMPL_WIDTH - 1),
		10080 => to_unsigned(26962, LUT_AMPL_WIDTH - 1),
		10081 => to_unsigned(26964, LUT_AMPL_WIDTH - 1),
		10082 => to_unsigned(26966, LUT_AMPL_WIDTH - 1),
		10083 => to_unsigned(26968, LUT_AMPL_WIDTH - 1),
		10084 => to_unsigned(26969, LUT_AMPL_WIDTH - 1),
		10085 => to_unsigned(26971, LUT_AMPL_WIDTH - 1),
		10086 => to_unsigned(26973, LUT_AMPL_WIDTH - 1),
		10087 => to_unsigned(26975, LUT_AMPL_WIDTH - 1),
		10088 => to_unsigned(26977, LUT_AMPL_WIDTH - 1),
		10089 => to_unsigned(26978, LUT_AMPL_WIDTH - 1),
		10090 => to_unsigned(26980, LUT_AMPL_WIDTH - 1),
		10091 => to_unsigned(26982, LUT_AMPL_WIDTH - 1),
		10092 => to_unsigned(26984, LUT_AMPL_WIDTH - 1),
		10093 => to_unsigned(26986, LUT_AMPL_WIDTH - 1),
		10094 => to_unsigned(26987, LUT_AMPL_WIDTH - 1),
		10095 => to_unsigned(26989, LUT_AMPL_WIDTH - 1),
		10096 => to_unsigned(26991, LUT_AMPL_WIDTH - 1),
		10097 => to_unsigned(26993, LUT_AMPL_WIDTH - 1),
		10098 => to_unsigned(26994, LUT_AMPL_WIDTH - 1),
		10099 => to_unsigned(26996, LUT_AMPL_WIDTH - 1),
		10100 => to_unsigned(26998, LUT_AMPL_WIDTH - 1),
		10101 => to_unsigned(27000, LUT_AMPL_WIDTH - 1),
		10102 => to_unsigned(27002, LUT_AMPL_WIDTH - 1),
		10103 => to_unsigned(27003, LUT_AMPL_WIDTH - 1),
		10104 => to_unsigned(27005, LUT_AMPL_WIDTH - 1),
		10105 => to_unsigned(27007, LUT_AMPL_WIDTH - 1),
		10106 => to_unsigned(27009, LUT_AMPL_WIDTH - 1),
		10107 => to_unsigned(27010, LUT_AMPL_WIDTH - 1),
		10108 => to_unsigned(27012, LUT_AMPL_WIDTH - 1),
		10109 => to_unsigned(27014, LUT_AMPL_WIDTH - 1),
		10110 => to_unsigned(27016, LUT_AMPL_WIDTH - 1),
		10111 => to_unsigned(27018, LUT_AMPL_WIDTH - 1),
		10112 => to_unsigned(27019, LUT_AMPL_WIDTH - 1),
		10113 => to_unsigned(27021, LUT_AMPL_WIDTH - 1),
		10114 => to_unsigned(27023, LUT_AMPL_WIDTH - 1),
		10115 => to_unsigned(27025, LUT_AMPL_WIDTH - 1),
		10116 => to_unsigned(27026, LUT_AMPL_WIDTH - 1),
		10117 => to_unsigned(27028, LUT_AMPL_WIDTH - 1),
		10118 => to_unsigned(27030, LUT_AMPL_WIDTH - 1),
		10119 => to_unsigned(27032, LUT_AMPL_WIDTH - 1),
		10120 => to_unsigned(27034, LUT_AMPL_WIDTH - 1),
		10121 => to_unsigned(27035, LUT_AMPL_WIDTH - 1),
		10122 => to_unsigned(27037, LUT_AMPL_WIDTH - 1),
		10123 => to_unsigned(27039, LUT_AMPL_WIDTH - 1),
		10124 => to_unsigned(27041, LUT_AMPL_WIDTH - 1),
		10125 => to_unsigned(27042, LUT_AMPL_WIDTH - 1),
		10126 => to_unsigned(27044, LUT_AMPL_WIDTH - 1),
		10127 => to_unsigned(27046, LUT_AMPL_WIDTH - 1),
		10128 => to_unsigned(27048, LUT_AMPL_WIDTH - 1),
		10129 => to_unsigned(27049, LUT_AMPL_WIDTH - 1),
		10130 => to_unsigned(27051, LUT_AMPL_WIDTH - 1),
		10131 => to_unsigned(27053, LUT_AMPL_WIDTH - 1),
		10132 => to_unsigned(27055, LUT_AMPL_WIDTH - 1),
		10133 => to_unsigned(27057, LUT_AMPL_WIDTH - 1),
		10134 => to_unsigned(27058, LUT_AMPL_WIDTH - 1),
		10135 => to_unsigned(27060, LUT_AMPL_WIDTH - 1),
		10136 => to_unsigned(27062, LUT_AMPL_WIDTH - 1),
		10137 => to_unsigned(27064, LUT_AMPL_WIDTH - 1),
		10138 => to_unsigned(27065, LUT_AMPL_WIDTH - 1),
		10139 => to_unsigned(27067, LUT_AMPL_WIDTH - 1),
		10140 => to_unsigned(27069, LUT_AMPL_WIDTH - 1),
		10141 => to_unsigned(27071, LUT_AMPL_WIDTH - 1),
		10142 => to_unsigned(27073, LUT_AMPL_WIDTH - 1),
		10143 => to_unsigned(27074, LUT_AMPL_WIDTH - 1),
		10144 => to_unsigned(27076, LUT_AMPL_WIDTH - 1),
		10145 => to_unsigned(27078, LUT_AMPL_WIDTH - 1),
		10146 => to_unsigned(27080, LUT_AMPL_WIDTH - 1),
		10147 => to_unsigned(27081, LUT_AMPL_WIDTH - 1),
		10148 => to_unsigned(27083, LUT_AMPL_WIDTH - 1),
		10149 => to_unsigned(27085, LUT_AMPL_WIDTH - 1),
		10150 => to_unsigned(27087, LUT_AMPL_WIDTH - 1),
		10151 => to_unsigned(27088, LUT_AMPL_WIDTH - 1),
		10152 => to_unsigned(27090, LUT_AMPL_WIDTH - 1),
		10153 => to_unsigned(27092, LUT_AMPL_WIDTH - 1),
		10154 => to_unsigned(27094, LUT_AMPL_WIDTH - 1),
		10155 => to_unsigned(27096, LUT_AMPL_WIDTH - 1),
		10156 => to_unsigned(27097, LUT_AMPL_WIDTH - 1),
		10157 => to_unsigned(27099, LUT_AMPL_WIDTH - 1),
		10158 => to_unsigned(27101, LUT_AMPL_WIDTH - 1),
		10159 => to_unsigned(27103, LUT_AMPL_WIDTH - 1),
		10160 => to_unsigned(27104, LUT_AMPL_WIDTH - 1),
		10161 => to_unsigned(27106, LUT_AMPL_WIDTH - 1),
		10162 => to_unsigned(27108, LUT_AMPL_WIDTH - 1),
		10163 => to_unsigned(27110, LUT_AMPL_WIDTH - 1),
		10164 => to_unsigned(27111, LUT_AMPL_WIDTH - 1),
		10165 => to_unsigned(27113, LUT_AMPL_WIDTH - 1),
		10166 => to_unsigned(27115, LUT_AMPL_WIDTH - 1),
		10167 => to_unsigned(27117, LUT_AMPL_WIDTH - 1),
		10168 => to_unsigned(27118, LUT_AMPL_WIDTH - 1),
		10169 => to_unsigned(27120, LUT_AMPL_WIDTH - 1),
		10170 => to_unsigned(27122, LUT_AMPL_WIDTH - 1),
		10171 => to_unsigned(27124, LUT_AMPL_WIDTH - 1),
		10172 => to_unsigned(27126, LUT_AMPL_WIDTH - 1),
		10173 => to_unsigned(27127, LUT_AMPL_WIDTH - 1),
		10174 => to_unsigned(27129, LUT_AMPL_WIDTH - 1),
		10175 => to_unsigned(27131, LUT_AMPL_WIDTH - 1),
		10176 => to_unsigned(27133, LUT_AMPL_WIDTH - 1),
		10177 => to_unsigned(27134, LUT_AMPL_WIDTH - 1),
		10178 => to_unsigned(27136, LUT_AMPL_WIDTH - 1),
		10179 => to_unsigned(27138, LUT_AMPL_WIDTH - 1),
		10180 => to_unsigned(27140, LUT_AMPL_WIDTH - 1),
		10181 => to_unsigned(27141, LUT_AMPL_WIDTH - 1),
		10182 => to_unsigned(27143, LUT_AMPL_WIDTH - 1),
		10183 => to_unsigned(27145, LUT_AMPL_WIDTH - 1),
		10184 => to_unsigned(27147, LUT_AMPL_WIDTH - 1),
		10185 => to_unsigned(27148, LUT_AMPL_WIDTH - 1),
		10186 => to_unsigned(27150, LUT_AMPL_WIDTH - 1),
		10187 => to_unsigned(27152, LUT_AMPL_WIDTH - 1),
		10188 => to_unsigned(27154, LUT_AMPL_WIDTH - 1),
		10189 => to_unsigned(27155, LUT_AMPL_WIDTH - 1),
		10190 => to_unsigned(27157, LUT_AMPL_WIDTH - 1),
		10191 => to_unsigned(27159, LUT_AMPL_WIDTH - 1),
		10192 => to_unsigned(27161, LUT_AMPL_WIDTH - 1),
		10193 => to_unsigned(27162, LUT_AMPL_WIDTH - 1),
		10194 => to_unsigned(27164, LUT_AMPL_WIDTH - 1),
		10195 => to_unsigned(27166, LUT_AMPL_WIDTH - 1),
		10196 => to_unsigned(27168, LUT_AMPL_WIDTH - 1),
		10197 => to_unsigned(27169, LUT_AMPL_WIDTH - 1),
		10198 => to_unsigned(27171, LUT_AMPL_WIDTH - 1),
		10199 => to_unsigned(27173, LUT_AMPL_WIDTH - 1),
		10200 => to_unsigned(27175, LUT_AMPL_WIDTH - 1),
		10201 => to_unsigned(27177, LUT_AMPL_WIDTH - 1),
		10202 => to_unsigned(27178, LUT_AMPL_WIDTH - 1),
		10203 => to_unsigned(27180, LUT_AMPL_WIDTH - 1),
		10204 => to_unsigned(27182, LUT_AMPL_WIDTH - 1),
		10205 => to_unsigned(27184, LUT_AMPL_WIDTH - 1),
		10206 => to_unsigned(27185, LUT_AMPL_WIDTH - 1),
		10207 => to_unsigned(27187, LUT_AMPL_WIDTH - 1),
		10208 => to_unsigned(27189, LUT_AMPL_WIDTH - 1),
		10209 => to_unsigned(27191, LUT_AMPL_WIDTH - 1),
		10210 => to_unsigned(27192, LUT_AMPL_WIDTH - 1),
		10211 => to_unsigned(27194, LUT_AMPL_WIDTH - 1),
		10212 => to_unsigned(27196, LUT_AMPL_WIDTH - 1),
		10213 => to_unsigned(27198, LUT_AMPL_WIDTH - 1),
		10214 => to_unsigned(27199, LUT_AMPL_WIDTH - 1),
		10215 => to_unsigned(27201, LUT_AMPL_WIDTH - 1),
		10216 => to_unsigned(27203, LUT_AMPL_WIDTH - 1),
		10217 => to_unsigned(27205, LUT_AMPL_WIDTH - 1),
		10218 => to_unsigned(27206, LUT_AMPL_WIDTH - 1),
		10219 => to_unsigned(27208, LUT_AMPL_WIDTH - 1),
		10220 => to_unsigned(27210, LUT_AMPL_WIDTH - 1),
		10221 => to_unsigned(27212, LUT_AMPL_WIDTH - 1),
		10222 => to_unsigned(27213, LUT_AMPL_WIDTH - 1),
		10223 => to_unsigned(27215, LUT_AMPL_WIDTH - 1),
		10224 => to_unsigned(27217, LUT_AMPL_WIDTH - 1),
		10225 => to_unsigned(27219, LUT_AMPL_WIDTH - 1),
		10226 => to_unsigned(27220, LUT_AMPL_WIDTH - 1),
		10227 => to_unsigned(27222, LUT_AMPL_WIDTH - 1),
		10228 => to_unsigned(27224, LUT_AMPL_WIDTH - 1),
		10229 => to_unsigned(27226, LUT_AMPL_WIDTH - 1),
		10230 => to_unsigned(27227, LUT_AMPL_WIDTH - 1),
		10231 => to_unsigned(27229, LUT_AMPL_WIDTH - 1),
		10232 => to_unsigned(27231, LUT_AMPL_WIDTH - 1),
		10233 => to_unsigned(27233, LUT_AMPL_WIDTH - 1),
		10234 => to_unsigned(27234, LUT_AMPL_WIDTH - 1),
		10235 => to_unsigned(27236, LUT_AMPL_WIDTH - 1),
		10236 => to_unsigned(27238, LUT_AMPL_WIDTH - 1),
		10237 => to_unsigned(27240, LUT_AMPL_WIDTH - 1),
		10238 => to_unsigned(27241, LUT_AMPL_WIDTH - 1),
		10239 => to_unsigned(27243, LUT_AMPL_WIDTH - 1),
		10240 => to_unsigned(27245, LUT_AMPL_WIDTH - 1),
		10241 => to_unsigned(27247, LUT_AMPL_WIDTH - 1),
		10242 => to_unsigned(27248, LUT_AMPL_WIDTH - 1),
		10243 => to_unsigned(27250, LUT_AMPL_WIDTH - 1),
		10244 => to_unsigned(27252, LUT_AMPL_WIDTH - 1),
		10245 => to_unsigned(27253, LUT_AMPL_WIDTH - 1),
		10246 => to_unsigned(27255, LUT_AMPL_WIDTH - 1),
		10247 => to_unsigned(27257, LUT_AMPL_WIDTH - 1),
		10248 => to_unsigned(27259, LUT_AMPL_WIDTH - 1),
		10249 => to_unsigned(27260, LUT_AMPL_WIDTH - 1),
		10250 => to_unsigned(27262, LUT_AMPL_WIDTH - 1),
		10251 => to_unsigned(27264, LUT_AMPL_WIDTH - 1),
		10252 => to_unsigned(27266, LUT_AMPL_WIDTH - 1),
		10253 => to_unsigned(27267, LUT_AMPL_WIDTH - 1),
		10254 => to_unsigned(27269, LUT_AMPL_WIDTH - 1),
		10255 => to_unsigned(27271, LUT_AMPL_WIDTH - 1),
		10256 => to_unsigned(27273, LUT_AMPL_WIDTH - 1),
		10257 => to_unsigned(27274, LUT_AMPL_WIDTH - 1),
		10258 => to_unsigned(27276, LUT_AMPL_WIDTH - 1),
		10259 => to_unsigned(27278, LUT_AMPL_WIDTH - 1),
		10260 => to_unsigned(27280, LUT_AMPL_WIDTH - 1),
		10261 => to_unsigned(27281, LUT_AMPL_WIDTH - 1),
		10262 => to_unsigned(27283, LUT_AMPL_WIDTH - 1),
		10263 => to_unsigned(27285, LUT_AMPL_WIDTH - 1),
		10264 => to_unsigned(27287, LUT_AMPL_WIDTH - 1),
		10265 => to_unsigned(27288, LUT_AMPL_WIDTH - 1),
		10266 => to_unsigned(27290, LUT_AMPL_WIDTH - 1),
		10267 => to_unsigned(27292, LUT_AMPL_WIDTH - 1),
		10268 => to_unsigned(27294, LUT_AMPL_WIDTH - 1),
		10269 => to_unsigned(27295, LUT_AMPL_WIDTH - 1),
		10270 => to_unsigned(27297, LUT_AMPL_WIDTH - 1),
		10271 => to_unsigned(27299, LUT_AMPL_WIDTH - 1),
		10272 => to_unsigned(27300, LUT_AMPL_WIDTH - 1),
		10273 => to_unsigned(27302, LUT_AMPL_WIDTH - 1),
		10274 => to_unsigned(27304, LUT_AMPL_WIDTH - 1),
		10275 => to_unsigned(27306, LUT_AMPL_WIDTH - 1),
		10276 => to_unsigned(27307, LUT_AMPL_WIDTH - 1),
		10277 => to_unsigned(27309, LUT_AMPL_WIDTH - 1),
		10278 => to_unsigned(27311, LUT_AMPL_WIDTH - 1),
		10279 => to_unsigned(27313, LUT_AMPL_WIDTH - 1),
		10280 => to_unsigned(27314, LUT_AMPL_WIDTH - 1),
		10281 => to_unsigned(27316, LUT_AMPL_WIDTH - 1),
		10282 => to_unsigned(27318, LUT_AMPL_WIDTH - 1),
		10283 => to_unsigned(27320, LUT_AMPL_WIDTH - 1),
		10284 => to_unsigned(27321, LUT_AMPL_WIDTH - 1),
		10285 => to_unsigned(27323, LUT_AMPL_WIDTH - 1),
		10286 => to_unsigned(27325, LUT_AMPL_WIDTH - 1),
		10287 => to_unsigned(27327, LUT_AMPL_WIDTH - 1),
		10288 => to_unsigned(27328, LUT_AMPL_WIDTH - 1),
		10289 => to_unsigned(27330, LUT_AMPL_WIDTH - 1),
		10290 => to_unsigned(27332, LUT_AMPL_WIDTH - 1),
		10291 => to_unsigned(27333, LUT_AMPL_WIDTH - 1),
		10292 => to_unsigned(27335, LUT_AMPL_WIDTH - 1),
		10293 => to_unsigned(27337, LUT_AMPL_WIDTH - 1),
		10294 => to_unsigned(27339, LUT_AMPL_WIDTH - 1),
		10295 => to_unsigned(27340, LUT_AMPL_WIDTH - 1),
		10296 => to_unsigned(27342, LUT_AMPL_WIDTH - 1),
		10297 => to_unsigned(27344, LUT_AMPL_WIDTH - 1),
		10298 => to_unsigned(27346, LUT_AMPL_WIDTH - 1),
		10299 => to_unsigned(27347, LUT_AMPL_WIDTH - 1),
		10300 => to_unsigned(27349, LUT_AMPL_WIDTH - 1),
		10301 => to_unsigned(27351, LUT_AMPL_WIDTH - 1),
		10302 => to_unsigned(27352, LUT_AMPL_WIDTH - 1),
		10303 => to_unsigned(27354, LUT_AMPL_WIDTH - 1),
		10304 => to_unsigned(27356, LUT_AMPL_WIDTH - 1),
		10305 => to_unsigned(27358, LUT_AMPL_WIDTH - 1),
		10306 => to_unsigned(27359, LUT_AMPL_WIDTH - 1),
		10307 => to_unsigned(27361, LUT_AMPL_WIDTH - 1),
		10308 => to_unsigned(27363, LUT_AMPL_WIDTH - 1),
		10309 => to_unsigned(27365, LUT_AMPL_WIDTH - 1),
		10310 => to_unsigned(27366, LUT_AMPL_WIDTH - 1),
		10311 => to_unsigned(27368, LUT_AMPL_WIDTH - 1),
		10312 => to_unsigned(27370, LUT_AMPL_WIDTH - 1),
		10313 => to_unsigned(27372, LUT_AMPL_WIDTH - 1),
		10314 => to_unsigned(27373, LUT_AMPL_WIDTH - 1),
		10315 => to_unsigned(27375, LUT_AMPL_WIDTH - 1),
		10316 => to_unsigned(27377, LUT_AMPL_WIDTH - 1),
		10317 => to_unsigned(27378, LUT_AMPL_WIDTH - 1),
		10318 => to_unsigned(27380, LUT_AMPL_WIDTH - 1),
		10319 => to_unsigned(27382, LUT_AMPL_WIDTH - 1),
		10320 => to_unsigned(27384, LUT_AMPL_WIDTH - 1),
		10321 => to_unsigned(27385, LUT_AMPL_WIDTH - 1),
		10322 => to_unsigned(27387, LUT_AMPL_WIDTH - 1),
		10323 => to_unsigned(27389, LUT_AMPL_WIDTH - 1),
		10324 => to_unsigned(27390, LUT_AMPL_WIDTH - 1),
		10325 => to_unsigned(27392, LUT_AMPL_WIDTH - 1),
		10326 => to_unsigned(27394, LUT_AMPL_WIDTH - 1),
		10327 => to_unsigned(27396, LUT_AMPL_WIDTH - 1),
		10328 => to_unsigned(27397, LUT_AMPL_WIDTH - 1),
		10329 => to_unsigned(27399, LUT_AMPL_WIDTH - 1),
		10330 => to_unsigned(27401, LUT_AMPL_WIDTH - 1),
		10331 => to_unsigned(27403, LUT_AMPL_WIDTH - 1),
		10332 => to_unsigned(27404, LUT_AMPL_WIDTH - 1),
		10333 => to_unsigned(27406, LUT_AMPL_WIDTH - 1),
		10334 => to_unsigned(27408, LUT_AMPL_WIDTH - 1),
		10335 => to_unsigned(27409, LUT_AMPL_WIDTH - 1),
		10336 => to_unsigned(27411, LUT_AMPL_WIDTH - 1),
		10337 => to_unsigned(27413, LUT_AMPL_WIDTH - 1),
		10338 => to_unsigned(27415, LUT_AMPL_WIDTH - 1),
		10339 => to_unsigned(27416, LUT_AMPL_WIDTH - 1),
		10340 => to_unsigned(27418, LUT_AMPL_WIDTH - 1),
		10341 => to_unsigned(27420, LUT_AMPL_WIDTH - 1),
		10342 => to_unsigned(27421, LUT_AMPL_WIDTH - 1),
		10343 => to_unsigned(27423, LUT_AMPL_WIDTH - 1),
		10344 => to_unsigned(27425, LUT_AMPL_WIDTH - 1),
		10345 => to_unsigned(27427, LUT_AMPL_WIDTH - 1),
		10346 => to_unsigned(27428, LUT_AMPL_WIDTH - 1),
		10347 => to_unsigned(27430, LUT_AMPL_WIDTH - 1),
		10348 => to_unsigned(27432, LUT_AMPL_WIDTH - 1),
		10349 => to_unsigned(27434, LUT_AMPL_WIDTH - 1),
		10350 => to_unsigned(27435, LUT_AMPL_WIDTH - 1),
		10351 => to_unsigned(27437, LUT_AMPL_WIDTH - 1),
		10352 => to_unsigned(27439, LUT_AMPL_WIDTH - 1),
		10353 => to_unsigned(27440, LUT_AMPL_WIDTH - 1),
		10354 => to_unsigned(27442, LUT_AMPL_WIDTH - 1),
		10355 => to_unsigned(27444, LUT_AMPL_WIDTH - 1),
		10356 => to_unsigned(27446, LUT_AMPL_WIDTH - 1),
		10357 => to_unsigned(27447, LUT_AMPL_WIDTH - 1),
		10358 => to_unsigned(27449, LUT_AMPL_WIDTH - 1),
		10359 => to_unsigned(27451, LUT_AMPL_WIDTH - 1),
		10360 => to_unsigned(27452, LUT_AMPL_WIDTH - 1),
		10361 => to_unsigned(27454, LUT_AMPL_WIDTH - 1),
		10362 => to_unsigned(27456, LUT_AMPL_WIDTH - 1),
		10363 => to_unsigned(27458, LUT_AMPL_WIDTH - 1),
		10364 => to_unsigned(27459, LUT_AMPL_WIDTH - 1),
		10365 => to_unsigned(27461, LUT_AMPL_WIDTH - 1),
		10366 => to_unsigned(27463, LUT_AMPL_WIDTH - 1),
		10367 => to_unsigned(27464, LUT_AMPL_WIDTH - 1),
		10368 => to_unsigned(27466, LUT_AMPL_WIDTH - 1),
		10369 => to_unsigned(27468, LUT_AMPL_WIDTH - 1),
		10370 => to_unsigned(27470, LUT_AMPL_WIDTH - 1),
		10371 => to_unsigned(27471, LUT_AMPL_WIDTH - 1),
		10372 => to_unsigned(27473, LUT_AMPL_WIDTH - 1),
		10373 => to_unsigned(27475, LUT_AMPL_WIDTH - 1),
		10374 => to_unsigned(27476, LUT_AMPL_WIDTH - 1),
		10375 => to_unsigned(27478, LUT_AMPL_WIDTH - 1),
		10376 => to_unsigned(27480, LUT_AMPL_WIDTH - 1),
		10377 => to_unsigned(27482, LUT_AMPL_WIDTH - 1),
		10378 => to_unsigned(27483, LUT_AMPL_WIDTH - 1),
		10379 => to_unsigned(27485, LUT_AMPL_WIDTH - 1),
		10380 => to_unsigned(27487, LUT_AMPL_WIDTH - 1),
		10381 => to_unsigned(27488, LUT_AMPL_WIDTH - 1),
		10382 => to_unsigned(27490, LUT_AMPL_WIDTH - 1),
		10383 => to_unsigned(27492, LUT_AMPL_WIDTH - 1),
		10384 => to_unsigned(27493, LUT_AMPL_WIDTH - 1),
		10385 => to_unsigned(27495, LUT_AMPL_WIDTH - 1),
		10386 => to_unsigned(27497, LUT_AMPL_WIDTH - 1),
		10387 => to_unsigned(27499, LUT_AMPL_WIDTH - 1),
		10388 => to_unsigned(27500, LUT_AMPL_WIDTH - 1),
		10389 => to_unsigned(27502, LUT_AMPL_WIDTH - 1),
		10390 => to_unsigned(27504, LUT_AMPL_WIDTH - 1),
		10391 => to_unsigned(27505, LUT_AMPL_WIDTH - 1),
		10392 => to_unsigned(27507, LUT_AMPL_WIDTH - 1),
		10393 => to_unsigned(27509, LUT_AMPL_WIDTH - 1),
		10394 => to_unsigned(27511, LUT_AMPL_WIDTH - 1),
		10395 => to_unsigned(27512, LUT_AMPL_WIDTH - 1),
		10396 => to_unsigned(27514, LUT_AMPL_WIDTH - 1),
		10397 => to_unsigned(27516, LUT_AMPL_WIDTH - 1),
		10398 => to_unsigned(27517, LUT_AMPL_WIDTH - 1),
		10399 => to_unsigned(27519, LUT_AMPL_WIDTH - 1),
		10400 => to_unsigned(27521, LUT_AMPL_WIDTH - 1),
		10401 => to_unsigned(27523, LUT_AMPL_WIDTH - 1),
		10402 => to_unsigned(27524, LUT_AMPL_WIDTH - 1),
		10403 => to_unsigned(27526, LUT_AMPL_WIDTH - 1),
		10404 => to_unsigned(27528, LUT_AMPL_WIDTH - 1),
		10405 => to_unsigned(27529, LUT_AMPL_WIDTH - 1),
		10406 => to_unsigned(27531, LUT_AMPL_WIDTH - 1),
		10407 => to_unsigned(27533, LUT_AMPL_WIDTH - 1),
		10408 => to_unsigned(27534, LUT_AMPL_WIDTH - 1),
		10409 => to_unsigned(27536, LUT_AMPL_WIDTH - 1),
		10410 => to_unsigned(27538, LUT_AMPL_WIDTH - 1),
		10411 => to_unsigned(27540, LUT_AMPL_WIDTH - 1),
		10412 => to_unsigned(27541, LUT_AMPL_WIDTH - 1),
		10413 => to_unsigned(27543, LUT_AMPL_WIDTH - 1),
		10414 => to_unsigned(27545, LUT_AMPL_WIDTH - 1),
		10415 => to_unsigned(27546, LUT_AMPL_WIDTH - 1),
		10416 => to_unsigned(27548, LUT_AMPL_WIDTH - 1),
		10417 => to_unsigned(27550, LUT_AMPL_WIDTH - 1),
		10418 => to_unsigned(27551, LUT_AMPL_WIDTH - 1),
		10419 => to_unsigned(27553, LUT_AMPL_WIDTH - 1),
		10420 => to_unsigned(27555, LUT_AMPL_WIDTH - 1),
		10421 => to_unsigned(27557, LUT_AMPL_WIDTH - 1),
		10422 => to_unsigned(27558, LUT_AMPL_WIDTH - 1),
		10423 => to_unsigned(27560, LUT_AMPL_WIDTH - 1),
		10424 => to_unsigned(27562, LUT_AMPL_WIDTH - 1),
		10425 => to_unsigned(27563, LUT_AMPL_WIDTH - 1),
		10426 => to_unsigned(27565, LUT_AMPL_WIDTH - 1),
		10427 => to_unsigned(27567, LUT_AMPL_WIDTH - 1),
		10428 => to_unsigned(27568, LUT_AMPL_WIDTH - 1),
		10429 => to_unsigned(27570, LUT_AMPL_WIDTH - 1),
		10430 => to_unsigned(27572, LUT_AMPL_WIDTH - 1),
		10431 => to_unsigned(27574, LUT_AMPL_WIDTH - 1),
		10432 => to_unsigned(27575, LUT_AMPL_WIDTH - 1),
		10433 => to_unsigned(27577, LUT_AMPL_WIDTH - 1),
		10434 => to_unsigned(27579, LUT_AMPL_WIDTH - 1),
		10435 => to_unsigned(27580, LUT_AMPL_WIDTH - 1),
		10436 => to_unsigned(27582, LUT_AMPL_WIDTH - 1),
		10437 => to_unsigned(27584, LUT_AMPL_WIDTH - 1),
		10438 => to_unsigned(27585, LUT_AMPL_WIDTH - 1),
		10439 => to_unsigned(27587, LUT_AMPL_WIDTH - 1),
		10440 => to_unsigned(27589, LUT_AMPL_WIDTH - 1),
		10441 => to_unsigned(27590, LUT_AMPL_WIDTH - 1),
		10442 => to_unsigned(27592, LUT_AMPL_WIDTH - 1),
		10443 => to_unsigned(27594, LUT_AMPL_WIDTH - 1),
		10444 => to_unsigned(27596, LUT_AMPL_WIDTH - 1),
		10445 => to_unsigned(27597, LUT_AMPL_WIDTH - 1),
		10446 => to_unsigned(27599, LUT_AMPL_WIDTH - 1),
		10447 => to_unsigned(27601, LUT_AMPL_WIDTH - 1),
		10448 => to_unsigned(27602, LUT_AMPL_WIDTH - 1),
		10449 => to_unsigned(27604, LUT_AMPL_WIDTH - 1),
		10450 => to_unsigned(27606, LUT_AMPL_WIDTH - 1),
		10451 => to_unsigned(27607, LUT_AMPL_WIDTH - 1),
		10452 => to_unsigned(27609, LUT_AMPL_WIDTH - 1),
		10453 => to_unsigned(27611, LUT_AMPL_WIDTH - 1),
		10454 => to_unsigned(27613, LUT_AMPL_WIDTH - 1),
		10455 => to_unsigned(27614, LUT_AMPL_WIDTH - 1),
		10456 => to_unsigned(27616, LUT_AMPL_WIDTH - 1),
		10457 => to_unsigned(27618, LUT_AMPL_WIDTH - 1),
		10458 => to_unsigned(27619, LUT_AMPL_WIDTH - 1),
		10459 => to_unsigned(27621, LUT_AMPL_WIDTH - 1),
		10460 => to_unsigned(27623, LUT_AMPL_WIDTH - 1),
		10461 => to_unsigned(27624, LUT_AMPL_WIDTH - 1),
		10462 => to_unsigned(27626, LUT_AMPL_WIDTH - 1),
		10463 => to_unsigned(27628, LUT_AMPL_WIDTH - 1),
		10464 => to_unsigned(27629, LUT_AMPL_WIDTH - 1),
		10465 => to_unsigned(27631, LUT_AMPL_WIDTH - 1),
		10466 => to_unsigned(27633, LUT_AMPL_WIDTH - 1),
		10467 => to_unsigned(27634, LUT_AMPL_WIDTH - 1),
		10468 => to_unsigned(27636, LUT_AMPL_WIDTH - 1),
		10469 => to_unsigned(27638, LUT_AMPL_WIDTH - 1),
		10470 => to_unsigned(27640, LUT_AMPL_WIDTH - 1),
		10471 => to_unsigned(27641, LUT_AMPL_WIDTH - 1),
		10472 => to_unsigned(27643, LUT_AMPL_WIDTH - 1),
		10473 => to_unsigned(27645, LUT_AMPL_WIDTH - 1),
		10474 => to_unsigned(27646, LUT_AMPL_WIDTH - 1),
		10475 => to_unsigned(27648, LUT_AMPL_WIDTH - 1),
		10476 => to_unsigned(27650, LUT_AMPL_WIDTH - 1),
		10477 => to_unsigned(27651, LUT_AMPL_WIDTH - 1),
		10478 => to_unsigned(27653, LUT_AMPL_WIDTH - 1),
		10479 => to_unsigned(27655, LUT_AMPL_WIDTH - 1),
		10480 => to_unsigned(27656, LUT_AMPL_WIDTH - 1),
		10481 => to_unsigned(27658, LUT_AMPL_WIDTH - 1),
		10482 => to_unsigned(27660, LUT_AMPL_WIDTH - 1),
		10483 => to_unsigned(27661, LUT_AMPL_WIDTH - 1),
		10484 => to_unsigned(27663, LUT_AMPL_WIDTH - 1),
		10485 => to_unsigned(27665, LUT_AMPL_WIDTH - 1),
		10486 => to_unsigned(27666, LUT_AMPL_WIDTH - 1),
		10487 => to_unsigned(27668, LUT_AMPL_WIDTH - 1),
		10488 => to_unsigned(27670, LUT_AMPL_WIDTH - 1),
		10489 => to_unsigned(27672, LUT_AMPL_WIDTH - 1),
		10490 => to_unsigned(27673, LUT_AMPL_WIDTH - 1),
		10491 => to_unsigned(27675, LUT_AMPL_WIDTH - 1),
		10492 => to_unsigned(27677, LUT_AMPL_WIDTH - 1),
		10493 => to_unsigned(27678, LUT_AMPL_WIDTH - 1),
		10494 => to_unsigned(27680, LUT_AMPL_WIDTH - 1),
		10495 => to_unsigned(27682, LUT_AMPL_WIDTH - 1),
		10496 => to_unsigned(27683, LUT_AMPL_WIDTH - 1),
		10497 => to_unsigned(27685, LUT_AMPL_WIDTH - 1),
		10498 => to_unsigned(27687, LUT_AMPL_WIDTH - 1),
		10499 => to_unsigned(27688, LUT_AMPL_WIDTH - 1),
		10500 => to_unsigned(27690, LUT_AMPL_WIDTH - 1),
		10501 => to_unsigned(27692, LUT_AMPL_WIDTH - 1),
		10502 => to_unsigned(27693, LUT_AMPL_WIDTH - 1),
		10503 => to_unsigned(27695, LUT_AMPL_WIDTH - 1),
		10504 => to_unsigned(27697, LUT_AMPL_WIDTH - 1),
		10505 => to_unsigned(27698, LUT_AMPL_WIDTH - 1),
		10506 => to_unsigned(27700, LUT_AMPL_WIDTH - 1),
		10507 => to_unsigned(27702, LUT_AMPL_WIDTH - 1),
		10508 => to_unsigned(27703, LUT_AMPL_WIDTH - 1),
		10509 => to_unsigned(27705, LUT_AMPL_WIDTH - 1),
		10510 => to_unsigned(27707, LUT_AMPL_WIDTH - 1),
		10511 => to_unsigned(27708, LUT_AMPL_WIDTH - 1),
		10512 => to_unsigned(27710, LUT_AMPL_WIDTH - 1),
		10513 => to_unsigned(27712, LUT_AMPL_WIDTH - 1),
		10514 => to_unsigned(27714, LUT_AMPL_WIDTH - 1),
		10515 => to_unsigned(27715, LUT_AMPL_WIDTH - 1),
		10516 => to_unsigned(27717, LUT_AMPL_WIDTH - 1),
		10517 => to_unsigned(27719, LUT_AMPL_WIDTH - 1),
		10518 => to_unsigned(27720, LUT_AMPL_WIDTH - 1),
		10519 => to_unsigned(27722, LUT_AMPL_WIDTH - 1),
		10520 => to_unsigned(27724, LUT_AMPL_WIDTH - 1),
		10521 => to_unsigned(27725, LUT_AMPL_WIDTH - 1),
		10522 => to_unsigned(27727, LUT_AMPL_WIDTH - 1),
		10523 => to_unsigned(27729, LUT_AMPL_WIDTH - 1),
		10524 => to_unsigned(27730, LUT_AMPL_WIDTH - 1),
		10525 => to_unsigned(27732, LUT_AMPL_WIDTH - 1),
		10526 => to_unsigned(27734, LUT_AMPL_WIDTH - 1),
		10527 => to_unsigned(27735, LUT_AMPL_WIDTH - 1),
		10528 => to_unsigned(27737, LUT_AMPL_WIDTH - 1),
		10529 => to_unsigned(27739, LUT_AMPL_WIDTH - 1),
		10530 => to_unsigned(27740, LUT_AMPL_WIDTH - 1),
		10531 => to_unsigned(27742, LUT_AMPL_WIDTH - 1),
		10532 => to_unsigned(27744, LUT_AMPL_WIDTH - 1),
		10533 => to_unsigned(27745, LUT_AMPL_WIDTH - 1),
		10534 => to_unsigned(27747, LUT_AMPL_WIDTH - 1),
		10535 => to_unsigned(27749, LUT_AMPL_WIDTH - 1),
		10536 => to_unsigned(27750, LUT_AMPL_WIDTH - 1),
		10537 => to_unsigned(27752, LUT_AMPL_WIDTH - 1),
		10538 => to_unsigned(27754, LUT_AMPL_WIDTH - 1),
		10539 => to_unsigned(27755, LUT_AMPL_WIDTH - 1),
		10540 => to_unsigned(27757, LUT_AMPL_WIDTH - 1),
		10541 => to_unsigned(27759, LUT_AMPL_WIDTH - 1),
		10542 => to_unsigned(27760, LUT_AMPL_WIDTH - 1),
		10543 => to_unsigned(27762, LUT_AMPL_WIDTH - 1),
		10544 => to_unsigned(27764, LUT_AMPL_WIDTH - 1),
		10545 => to_unsigned(27765, LUT_AMPL_WIDTH - 1),
		10546 => to_unsigned(27767, LUT_AMPL_WIDTH - 1),
		10547 => to_unsigned(27769, LUT_AMPL_WIDTH - 1),
		10548 => to_unsigned(27770, LUT_AMPL_WIDTH - 1),
		10549 => to_unsigned(27772, LUT_AMPL_WIDTH - 1),
		10550 => to_unsigned(27774, LUT_AMPL_WIDTH - 1),
		10551 => to_unsigned(27775, LUT_AMPL_WIDTH - 1),
		10552 => to_unsigned(27777, LUT_AMPL_WIDTH - 1),
		10553 => to_unsigned(27779, LUT_AMPL_WIDTH - 1),
		10554 => to_unsigned(27780, LUT_AMPL_WIDTH - 1),
		10555 => to_unsigned(27782, LUT_AMPL_WIDTH - 1),
		10556 => to_unsigned(27784, LUT_AMPL_WIDTH - 1),
		10557 => to_unsigned(27785, LUT_AMPL_WIDTH - 1),
		10558 => to_unsigned(27787, LUT_AMPL_WIDTH - 1),
		10559 => to_unsigned(27789, LUT_AMPL_WIDTH - 1),
		10560 => to_unsigned(27790, LUT_AMPL_WIDTH - 1),
		10561 => to_unsigned(27792, LUT_AMPL_WIDTH - 1),
		10562 => to_unsigned(27794, LUT_AMPL_WIDTH - 1),
		10563 => to_unsigned(27795, LUT_AMPL_WIDTH - 1),
		10564 => to_unsigned(27797, LUT_AMPL_WIDTH - 1),
		10565 => to_unsigned(27799, LUT_AMPL_WIDTH - 1),
		10566 => to_unsigned(27800, LUT_AMPL_WIDTH - 1),
		10567 => to_unsigned(27802, LUT_AMPL_WIDTH - 1),
		10568 => to_unsigned(27804, LUT_AMPL_WIDTH - 1),
		10569 => to_unsigned(27805, LUT_AMPL_WIDTH - 1),
		10570 => to_unsigned(27807, LUT_AMPL_WIDTH - 1),
		10571 => to_unsigned(27809, LUT_AMPL_WIDTH - 1),
		10572 => to_unsigned(27810, LUT_AMPL_WIDTH - 1),
		10573 => to_unsigned(27812, LUT_AMPL_WIDTH - 1),
		10574 => to_unsigned(27814, LUT_AMPL_WIDTH - 1),
		10575 => to_unsigned(27815, LUT_AMPL_WIDTH - 1),
		10576 => to_unsigned(27817, LUT_AMPL_WIDTH - 1),
		10577 => to_unsigned(27819, LUT_AMPL_WIDTH - 1),
		10578 => to_unsigned(27820, LUT_AMPL_WIDTH - 1),
		10579 => to_unsigned(27822, LUT_AMPL_WIDTH - 1),
		10580 => to_unsigned(27824, LUT_AMPL_WIDTH - 1),
		10581 => to_unsigned(27825, LUT_AMPL_WIDTH - 1),
		10582 => to_unsigned(27827, LUT_AMPL_WIDTH - 1),
		10583 => to_unsigned(27829, LUT_AMPL_WIDTH - 1),
		10584 => to_unsigned(27830, LUT_AMPL_WIDTH - 1),
		10585 => to_unsigned(27832, LUT_AMPL_WIDTH - 1),
		10586 => to_unsigned(27834, LUT_AMPL_WIDTH - 1),
		10587 => to_unsigned(27835, LUT_AMPL_WIDTH - 1),
		10588 => to_unsigned(27837, LUT_AMPL_WIDTH - 1),
		10589 => to_unsigned(27839, LUT_AMPL_WIDTH - 1),
		10590 => to_unsigned(27840, LUT_AMPL_WIDTH - 1),
		10591 => to_unsigned(27842, LUT_AMPL_WIDTH - 1),
		10592 => to_unsigned(27843, LUT_AMPL_WIDTH - 1),
		10593 => to_unsigned(27845, LUT_AMPL_WIDTH - 1),
		10594 => to_unsigned(27847, LUT_AMPL_WIDTH - 1),
		10595 => to_unsigned(27848, LUT_AMPL_WIDTH - 1),
		10596 => to_unsigned(27850, LUT_AMPL_WIDTH - 1),
		10597 => to_unsigned(27852, LUT_AMPL_WIDTH - 1),
		10598 => to_unsigned(27853, LUT_AMPL_WIDTH - 1),
		10599 => to_unsigned(27855, LUT_AMPL_WIDTH - 1),
		10600 => to_unsigned(27857, LUT_AMPL_WIDTH - 1),
		10601 => to_unsigned(27858, LUT_AMPL_WIDTH - 1),
		10602 => to_unsigned(27860, LUT_AMPL_WIDTH - 1),
		10603 => to_unsigned(27862, LUT_AMPL_WIDTH - 1),
		10604 => to_unsigned(27863, LUT_AMPL_WIDTH - 1),
		10605 => to_unsigned(27865, LUT_AMPL_WIDTH - 1),
		10606 => to_unsigned(27867, LUT_AMPL_WIDTH - 1),
		10607 => to_unsigned(27868, LUT_AMPL_WIDTH - 1),
		10608 => to_unsigned(27870, LUT_AMPL_WIDTH - 1),
		10609 => to_unsigned(27872, LUT_AMPL_WIDTH - 1),
		10610 => to_unsigned(27873, LUT_AMPL_WIDTH - 1),
		10611 => to_unsigned(27875, LUT_AMPL_WIDTH - 1),
		10612 => to_unsigned(27877, LUT_AMPL_WIDTH - 1),
		10613 => to_unsigned(27878, LUT_AMPL_WIDTH - 1),
		10614 => to_unsigned(27880, LUT_AMPL_WIDTH - 1),
		10615 => to_unsigned(27882, LUT_AMPL_WIDTH - 1),
		10616 => to_unsigned(27883, LUT_AMPL_WIDTH - 1),
		10617 => to_unsigned(27885, LUT_AMPL_WIDTH - 1),
		10618 => to_unsigned(27886, LUT_AMPL_WIDTH - 1),
		10619 => to_unsigned(27888, LUT_AMPL_WIDTH - 1),
		10620 => to_unsigned(27890, LUT_AMPL_WIDTH - 1),
		10621 => to_unsigned(27891, LUT_AMPL_WIDTH - 1),
		10622 => to_unsigned(27893, LUT_AMPL_WIDTH - 1),
		10623 => to_unsigned(27895, LUT_AMPL_WIDTH - 1),
		10624 => to_unsigned(27896, LUT_AMPL_WIDTH - 1),
		10625 => to_unsigned(27898, LUT_AMPL_WIDTH - 1),
		10626 => to_unsigned(27900, LUT_AMPL_WIDTH - 1),
		10627 => to_unsigned(27901, LUT_AMPL_WIDTH - 1),
		10628 => to_unsigned(27903, LUT_AMPL_WIDTH - 1),
		10629 => to_unsigned(27905, LUT_AMPL_WIDTH - 1),
		10630 => to_unsigned(27906, LUT_AMPL_WIDTH - 1),
		10631 => to_unsigned(27908, LUT_AMPL_WIDTH - 1),
		10632 => to_unsigned(27910, LUT_AMPL_WIDTH - 1),
		10633 => to_unsigned(27911, LUT_AMPL_WIDTH - 1),
		10634 => to_unsigned(27913, LUT_AMPL_WIDTH - 1),
		10635 => to_unsigned(27914, LUT_AMPL_WIDTH - 1),
		10636 => to_unsigned(27916, LUT_AMPL_WIDTH - 1),
		10637 => to_unsigned(27918, LUT_AMPL_WIDTH - 1),
		10638 => to_unsigned(27919, LUT_AMPL_WIDTH - 1),
		10639 => to_unsigned(27921, LUT_AMPL_WIDTH - 1),
		10640 => to_unsigned(27923, LUT_AMPL_WIDTH - 1),
		10641 => to_unsigned(27924, LUT_AMPL_WIDTH - 1),
		10642 => to_unsigned(27926, LUT_AMPL_WIDTH - 1),
		10643 => to_unsigned(27928, LUT_AMPL_WIDTH - 1),
		10644 => to_unsigned(27929, LUT_AMPL_WIDTH - 1),
		10645 => to_unsigned(27931, LUT_AMPL_WIDTH - 1),
		10646 => to_unsigned(27933, LUT_AMPL_WIDTH - 1),
		10647 => to_unsigned(27934, LUT_AMPL_WIDTH - 1),
		10648 => to_unsigned(27936, LUT_AMPL_WIDTH - 1),
		10649 => to_unsigned(27937, LUT_AMPL_WIDTH - 1),
		10650 => to_unsigned(27939, LUT_AMPL_WIDTH - 1),
		10651 => to_unsigned(27941, LUT_AMPL_WIDTH - 1),
		10652 => to_unsigned(27942, LUT_AMPL_WIDTH - 1),
		10653 => to_unsigned(27944, LUT_AMPL_WIDTH - 1),
		10654 => to_unsigned(27946, LUT_AMPL_WIDTH - 1),
		10655 => to_unsigned(27947, LUT_AMPL_WIDTH - 1),
		10656 => to_unsigned(27949, LUT_AMPL_WIDTH - 1),
		10657 => to_unsigned(27951, LUT_AMPL_WIDTH - 1),
		10658 => to_unsigned(27952, LUT_AMPL_WIDTH - 1),
		10659 => to_unsigned(27954, LUT_AMPL_WIDTH - 1),
		10660 => to_unsigned(27956, LUT_AMPL_WIDTH - 1),
		10661 => to_unsigned(27957, LUT_AMPL_WIDTH - 1),
		10662 => to_unsigned(27959, LUT_AMPL_WIDTH - 1),
		10663 => to_unsigned(27960, LUT_AMPL_WIDTH - 1),
		10664 => to_unsigned(27962, LUT_AMPL_WIDTH - 1),
		10665 => to_unsigned(27964, LUT_AMPL_WIDTH - 1),
		10666 => to_unsigned(27965, LUT_AMPL_WIDTH - 1),
		10667 => to_unsigned(27967, LUT_AMPL_WIDTH - 1),
		10668 => to_unsigned(27969, LUT_AMPL_WIDTH - 1),
		10669 => to_unsigned(27970, LUT_AMPL_WIDTH - 1),
		10670 => to_unsigned(27972, LUT_AMPL_WIDTH - 1),
		10671 => to_unsigned(27974, LUT_AMPL_WIDTH - 1),
		10672 => to_unsigned(27975, LUT_AMPL_WIDTH - 1),
		10673 => to_unsigned(27977, LUT_AMPL_WIDTH - 1),
		10674 => to_unsigned(27978, LUT_AMPL_WIDTH - 1),
		10675 => to_unsigned(27980, LUT_AMPL_WIDTH - 1),
		10676 => to_unsigned(27982, LUT_AMPL_WIDTH - 1),
		10677 => to_unsigned(27983, LUT_AMPL_WIDTH - 1),
		10678 => to_unsigned(27985, LUT_AMPL_WIDTH - 1),
		10679 => to_unsigned(27987, LUT_AMPL_WIDTH - 1),
		10680 => to_unsigned(27988, LUT_AMPL_WIDTH - 1),
		10681 => to_unsigned(27990, LUT_AMPL_WIDTH - 1),
		10682 => to_unsigned(27992, LUT_AMPL_WIDTH - 1),
		10683 => to_unsigned(27993, LUT_AMPL_WIDTH - 1),
		10684 => to_unsigned(27995, LUT_AMPL_WIDTH - 1),
		10685 => to_unsigned(27996, LUT_AMPL_WIDTH - 1),
		10686 => to_unsigned(27998, LUT_AMPL_WIDTH - 1),
		10687 => to_unsigned(28000, LUT_AMPL_WIDTH - 1),
		10688 => to_unsigned(28001, LUT_AMPL_WIDTH - 1),
		10689 => to_unsigned(28003, LUT_AMPL_WIDTH - 1),
		10690 => to_unsigned(28005, LUT_AMPL_WIDTH - 1),
		10691 => to_unsigned(28006, LUT_AMPL_WIDTH - 1),
		10692 => to_unsigned(28008, LUT_AMPL_WIDTH - 1),
		10693 => to_unsigned(28009, LUT_AMPL_WIDTH - 1),
		10694 => to_unsigned(28011, LUT_AMPL_WIDTH - 1),
		10695 => to_unsigned(28013, LUT_AMPL_WIDTH - 1),
		10696 => to_unsigned(28014, LUT_AMPL_WIDTH - 1),
		10697 => to_unsigned(28016, LUT_AMPL_WIDTH - 1),
		10698 => to_unsigned(28018, LUT_AMPL_WIDTH - 1),
		10699 => to_unsigned(28019, LUT_AMPL_WIDTH - 1),
		10700 => to_unsigned(28021, LUT_AMPL_WIDTH - 1),
		10701 => to_unsigned(28022, LUT_AMPL_WIDTH - 1),
		10702 => to_unsigned(28024, LUT_AMPL_WIDTH - 1),
		10703 => to_unsigned(28026, LUT_AMPL_WIDTH - 1),
		10704 => to_unsigned(28027, LUT_AMPL_WIDTH - 1),
		10705 => to_unsigned(28029, LUT_AMPL_WIDTH - 1),
		10706 => to_unsigned(28031, LUT_AMPL_WIDTH - 1),
		10707 => to_unsigned(28032, LUT_AMPL_WIDTH - 1),
		10708 => to_unsigned(28034, LUT_AMPL_WIDTH - 1),
		10709 => to_unsigned(28036, LUT_AMPL_WIDTH - 1),
		10710 => to_unsigned(28037, LUT_AMPL_WIDTH - 1),
		10711 => to_unsigned(28039, LUT_AMPL_WIDTH - 1),
		10712 => to_unsigned(28040, LUT_AMPL_WIDTH - 1),
		10713 => to_unsigned(28042, LUT_AMPL_WIDTH - 1),
		10714 => to_unsigned(28044, LUT_AMPL_WIDTH - 1),
		10715 => to_unsigned(28045, LUT_AMPL_WIDTH - 1),
		10716 => to_unsigned(28047, LUT_AMPL_WIDTH - 1),
		10717 => to_unsigned(28049, LUT_AMPL_WIDTH - 1),
		10718 => to_unsigned(28050, LUT_AMPL_WIDTH - 1),
		10719 => to_unsigned(28052, LUT_AMPL_WIDTH - 1),
		10720 => to_unsigned(28053, LUT_AMPL_WIDTH - 1),
		10721 => to_unsigned(28055, LUT_AMPL_WIDTH - 1),
		10722 => to_unsigned(28057, LUT_AMPL_WIDTH - 1),
		10723 => to_unsigned(28058, LUT_AMPL_WIDTH - 1),
		10724 => to_unsigned(28060, LUT_AMPL_WIDTH - 1),
		10725 => to_unsigned(28061, LUT_AMPL_WIDTH - 1),
		10726 => to_unsigned(28063, LUT_AMPL_WIDTH - 1),
		10727 => to_unsigned(28065, LUT_AMPL_WIDTH - 1),
		10728 => to_unsigned(28066, LUT_AMPL_WIDTH - 1),
		10729 => to_unsigned(28068, LUT_AMPL_WIDTH - 1),
		10730 => to_unsigned(28070, LUT_AMPL_WIDTH - 1),
		10731 => to_unsigned(28071, LUT_AMPL_WIDTH - 1),
		10732 => to_unsigned(28073, LUT_AMPL_WIDTH - 1),
		10733 => to_unsigned(28074, LUT_AMPL_WIDTH - 1),
		10734 => to_unsigned(28076, LUT_AMPL_WIDTH - 1),
		10735 => to_unsigned(28078, LUT_AMPL_WIDTH - 1),
		10736 => to_unsigned(28079, LUT_AMPL_WIDTH - 1),
		10737 => to_unsigned(28081, LUT_AMPL_WIDTH - 1),
		10738 => to_unsigned(28083, LUT_AMPL_WIDTH - 1),
		10739 => to_unsigned(28084, LUT_AMPL_WIDTH - 1),
		10740 => to_unsigned(28086, LUT_AMPL_WIDTH - 1),
		10741 => to_unsigned(28087, LUT_AMPL_WIDTH - 1),
		10742 => to_unsigned(28089, LUT_AMPL_WIDTH - 1),
		10743 => to_unsigned(28091, LUT_AMPL_WIDTH - 1),
		10744 => to_unsigned(28092, LUT_AMPL_WIDTH - 1),
		10745 => to_unsigned(28094, LUT_AMPL_WIDTH - 1),
		10746 => to_unsigned(28095, LUT_AMPL_WIDTH - 1),
		10747 => to_unsigned(28097, LUT_AMPL_WIDTH - 1),
		10748 => to_unsigned(28099, LUT_AMPL_WIDTH - 1),
		10749 => to_unsigned(28100, LUT_AMPL_WIDTH - 1),
		10750 => to_unsigned(28102, LUT_AMPL_WIDTH - 1),
		10751 => to_unsigned(28104, LUT_AMPL_WIDTH - 1),
		10752 => to_unsigned(28105, LUT_AMPL_WIDTH - 1),
		10753 => to_unsigned(28107, LUT_AMPL_WIDTH - 1),
		10754 => to_unsigned(28108, LUT_AMPL_WIDTH - 1),
		10755 => to_unsigned(28110, LUT_AMPL_WIDTH - 1),
		10756 => to_unsigned(28112, LUT_AMPL_WIDTH - 1),
		10757 => to_unsigned(28113, LUT_AMPL_WIDTH - 1),
		10758 => to_unsigned(28115, LUT_AMPL_WIDTH - 1),
		10759 => to_unsigned(28116, LUT_AMPL_WIDTH - 1),
		10760 => to_unsigned(28118, LUT_AMPL_WIDTH - 1),
		10761 => to_unsigned(28120, LUT_AMPL_WIDTH - 1),
		10762 => to_unsigned(28121, LUT_AMPL_WIDTH - 1),
		10763 => to_unsigned(28123, LUT_AMPL_WIDTH - 1),
		10764 => to_unsigned(28125, LUT_AMPL_WIDTH - 1),
		10765 => to_unsigned(28126, LUT_AMPL_WIDTH - 1),
		10766 => to_unsigned(28128, LUT_AMPL_WIDTH - 1),
		10767 => to_unsigned(28129, LUT_AMPL_WIDTH - 1),
		10768 => to_unsigned(28131, LUT_AMPL_WIDTH - 1),
		10769 => to_unsigned(28133, LUT_AMPL_WIDTH - 1),
		10770 => to_unsigned(28134, LUT_AMPL_WIDTH - 1),
		10771 => to_unsigned(28136, LUT_AMPL_WIDTH - 1),
		10772 => to_unsigned(28137, LUT_AMPL_WIDTH - 1),
		10773 => to_unsigned(28139, LUT_AMPL_WIDTH - 1),
		10774 => to_unsigned(28141, LUT_AMPL_WIDTH - 1),
		10775 => to_unsigned(28142, LUT_AMPL_WIDTH - 1),
		10776 => to_unsigned(28144, LUT_AMPL_WIDTH - 1),
		10777 => to_unsigned(28145, LUT_AMPL_WIDTH - 1),
		10778 => to_unsigned(28147, LUT_AMPL_WIDTH - 1),
		10779 => to_unsigned(28149, LUT_AMPL_WIDTH - 1),
		10780 => to_unsigned(28150, LUT_AMPL_WIDTH - 1),
		10781 => to_unsigned(28152, LUT_AMPL_WIDTH - 1),
		10782 => to_unsigned(28154, LUT_AMPL_WIDTH - 1),
		10783 => to_unsigned(28155, LUT_AMPL_WIDTH - 1),
		10784 => to_unsigned(28157, LUT_AMPL_WIDTH - 1),
		10785 => to_unsigned(28158, LUT_AMPL_WIDTH - 1),
		10786 => to_unsigned(28160, LUT_AMPL_WIDTH - 1),
		10787 => to_unsigned(28162, LUT_AMPL_WIDTH - 1),
		10788 => to_unsigned(28163, LUT_AMPL_WIDTH - 1),
		10789 => to_unsigned(28165, LUT_AMPL_WIDTH - 1),
		10790 => to_unsigned(28166, LUT_AMPL_WIDTH - 1),
		10791 => to_unsigned(28168, LUT_AMPL_WIDTH - 1),
		10792 => to_unsigned(28170, LUT_AMPL_WIDTH - 1),
		10793 => to_unsigned(28171, LUT_AMPL_WIDTH - 1),
		10794 => to_unsigned(28173, LUT_AMPL_WIDTH - 1),
		10795 => to_unsigned(28174, LUT_AMPL_WIDTH - 1),
		10796 => to_unsigned(28176, LUT_AMPL_WIDTH - 1),
		10797 => to_unsigned(28178, LUT_AMPL_WIDTH - 1),
		10798 => to_unsigned(28179, LUT_AMPL_WIDTH - 1),
		10799 => to_unsigned(28181, LUT_AMPL_WIDTH - 1),
		10800 => to_unsigned(28182, LUT_AMPL_WIDTH - 1),
		10801 => to_unsigned(28184, LUT_AMPL_WIDTH - 1),
		10802 => to_unsigned(28186, LUT_AMPL_WIDTH - 1),
		10803 => to_unsigned(28187, LUT_AMPL_WIDTH - 1),
		10804 => to_unsigned(28189, LUT_AMPL_WIDTH - 1),
		10805 => to_unsigned(28190, LUT_AMPL_WIDTH - 1),
		10806 => to_unsigned(28192, LUT_AMPL_WIDTH - 1),
		10807 => to_unsigned(28194, LUT_AMPL_WIDTH - 1),
		10808 => to_unsigned(28195, LUT_AMPL_WIDTH - 1),
		10809 => to_unsigned(28197, LUT_AMPL_WIDTH - 1),
		10810 => to_unsigned(28198, LUT_AMPL_WIDTH - 1),
		10811 => to_unsigned(28200, LUT_AMPL_WIDTH - 1),
		10812 => to_unsigned(28202, LUT_AMPL_WIDTH - 1),
		10813 => to_unsigned(28203, LUT_AMPL_WIDTH - 1),
		10814 => to_unsigned(28205, LUT_AMPL_WIDTH - 1),
		10815 => to_unsigned(28206, LUT_AMPL_WIDTH - 1),
		10816 => to_unsigned(28208, LUT_AMPL_WIDTH - 1),
		10817 => to_unsigned(28210, LUT_AMPL_WIDTH - 1),
		10818 => to_unsigned(28211, LUT_AMPL_WIDTH - 1),
		10819 => to_unsigned(28213, LUT_AMPL_WIDTH - 1),
		10820 => to_unsigned(28214, LUT_AMPL_WIDTH - 1),
		10821 => to_unsigned(28216, LUT_AMPL_WIDTH - 1),
		10822 => to_unsigned(28218, LUT_AMPL_WIDTH - 1),
		10823 => to_unsigned(28219, LUT_AMPL_WIDTH - 1),
		10824 => to_unsigned(28221, LUT_AMPL_WIDTH - 1),
		10825 => to_unsigned(28222, LUT_AMPL_WIDTH - 1),
		10826 => to_unsigned(28224, LUT_AMPL_WIDTH - 1),
		10827 => to_unsigned(28226, LUT_AMPL_WIDTH - 1),
		10828 => to_unsigned(28227, LUT_AMPL_WIDTH - 1),
		10829 => to_unsigned(28229, LUT_AMPL_WIDTH - 1),
		10830 => to_unsigned(28230, LUT_AMPL_WIDTH - 1),
		10831 => to_unsigned(28232, LUT_AMPL_WIDTH - 1),
		10832 => to_unsigned(28234, LUT_AMPL_WIDTH - 1),
		10833 => to_unsigned(28235, LUT_AMPL_WIDTH - 1),
		10834 => to_unsigned(28237, LUT_AMPL_WIDTH - 1),
		10835 => to_unsigned(28238, LUT_AMPL_WIDTH - 1),
		10836 => to_unsigned(28240, LUT_AMPL_WIDTH - 1),
		10837 => to_unsigned(28242, LUT_AMPL_WIDTH - 1),
		10838 => to_unsigned(28243, LUT_AMPL_WIDTH - 1),
		10839 => to_unsigned(28245, LUT_AMPL_WIDTH - 1),
		10840 => to_unsigned(28246, LUT_AMPL_WIDTH - 1),
		10841 => to_unsigned(28248, LUT_AMPL_WIDTH - 1),
		10842 => to_unsigned(28249, LUT_AMPL_WIDTH - 1),
		10843 => to_unsigned(28251, LUT_AMPL_WIDTH - 1),
		10844 => to_unsigned(28253, LUT_AMPL_WIDTH - 1),
		10845 => to_unsigned(28254, LUT_AMPL_WIDTH - 1),
		10846 => to_unsigned(28256, LUT_AMPL_WIDTH - 1),
		10847 => to_unsigned(28257, LUT_AMPL_WIDTH - 1),
		10848 => to_unsigned(28259, LUT_AMPL_WIDTH - 1),
		10849 => to_unsigned(28261, LUT_AMPL_WIDTH - 1),
		10850 => to_unsigned(28262, LUT_AMPL_WIDTH - 1),
		10851 => to_unsigned(28264, LUT_AMPL_WIDTH - 1),
		10852 => to_unsigned(28265, LUT_AMPL_WIDTH - 1),
		10853 => to_unsigned(28267, LUT_AMPL_WIDTH - 1),
		10854 => to_unsigned(28269, LUT_AMPL_WIDTH - 1),
		10855 => to_unsigned(28270, LUT_AMPL_WIDTH - 1),
		10856 => to_unsigned(28272, LUT_AMPL_WIDTH - 1),
		10857 => to_unsigned(28273, LUT_AMPL_WIDTH - 1),
		10858 => to_unsigned(28275, LUT_AMPL_WIDTH - 1),
		10859 => to_unsigned(28277, LUT_AMPL_WIDTH - 1),
		10860 => to_unsigned(28278, LUT_AMPL_WIDTH - 1),
		10861 => to_unsigned(28280, LUT_AMPL_WIDTH - 1),
		10862 => to_unsigned(28281, LUT_AMPL_WIDTH - 1),
		10863 => to_unsigned(28283, LUT_AMPL_WIDTH - 1),
		10864 => to_unsigned(28284, LUT_AMPL_WIDTH - 1),
		10865 => to_unsigned(28286, LUT_AMPL_WIDTH - 1),
		10866 => to_unsigned(28288, LUT_AMPL_WIDTH - 1),
		10867 => to_unsigned(28289, LUT_AMPL_WIDTH - 1),
		10868 => to_unsigned(28291, LUT_AMPL_WIDTH - 1),
		10869 => to_unsigned(28292, LUT_AMPL_WIDTH - 1),
		10870 => to_unsigned(28294, LUT_AMPL_WIDTH - 1),
		10871 => to_unsigned(28296, LUT_AMPL_WIDTH - 1),
		10872 => to_unsigned(28297, LUT_AMPL_WIDTH - 1),
		10873 => to_unsigned(28299, LUT_AMPL_WIDTH - 1),
		10874 => to_unsigned(28300, LUT_AMPL_WIDTH - 1),
		10875 => to_unsigned(28302, LUT_AMPL_WIDTH - 1),
		10876 => to_unsigned(28303, LUT_AMPL_WIDTH - 1),
		10877 => to_unsigned(28305, LUT_AMPL_WIDTH - 1),
		10878 => to_unsigned(28307, LUT_AMPL_WIDTH - 1),
		10879 => to_unsigned(28308, LUT_AMPL_WIDTH - 1),
		10880 => to_unsigned(28310, LUT_AMPL_WIDTH - 1),
		10881 => to_unsigned(28311, LUT_AMPL_WIDTH - 1),
		10882 => to_unsigned(28313, LUT_AMPL_WIDTH - 1),
		10883 => to_unsigned(28315, LUT_AMPL_WIDTH - 1),
		10884 => to_unsigned(28316, LUT_AMPL_WIDTH - 1),
		10885 => to_unsigned(28318, LUT_AMPL_WIDTH - 1),
		10886 => to_unsigned(28319, LUT_AMPL_WIDTH - 1),
		10887 => to_unsigned(28321, LUT_AMPL_WIDTH - 1),
		10888 => to_unsigned(28322, LUT_AMPL_WIDTH - 1),
		10889 => to_unsigned(28324, LUT_AMPL_WIDTH - 1),
		10890 => to_unsigned(28326, LUT_AMPL_WIDTH - 1),
		10891 => to_unsigned(28327, LUT_AMPL_WIDTH - 1),
		10892 => to_unsigned(28329, LUT_AMPL_WIDTH - 1),
		10893 => to_unsigned(28330, LUT_AMPL_WIDTH - 1),
		10894 => to_unsigned(28332, LUT_AMPL_WIDTH - 1),
		10895 => to_unsigned(28333, LUT_AMPL_WIDTH - 1),
		10896 => to_unsigned(28335, LUT_AMPL_WIDTH - 1),
		10897 => to_unsigned(28337, LUT_AMPL_WIDTH - 1),
		10898 => to_unsigned(28338, LUT_AMPL_WIDTH - 1),
		10899 => to_unsigned(28340, LUT_AMPL_WIDTH - 1),
		10900 => to_unsigned(28341, LUT_AMPL_WIDTH - 1),
		10901 => to_unsigned(28343, LUT_AMPL_WIDTH - 1),
		10902 => to_unsigned(28345, LUT_AMPL_WIDTH - 1),
		10903 => to_unsigned(28346, LUT_AMPL_WIDTH - 1),
		10904 => to_unsigned(28348, LUT_AMPL_WIDTH - 1),
		10905 => to_unsigned(28349, LUT_AMPL_WIDTH - 1),
		10906 => to_unsigned(28351, LUT_AMPL_WIDTH - 1),
		10907 => to_unsigned(28352, LUT_AMPL_WIDTH - 1),
		10908 => to_unsigned(28354, LUT_AMPL_WIDTH - 1),
		10909 => to_unsigned(28356, LUT_AMPL_WIDTH - 1),
		10910 => to_unsigned(28357, LUT_AMPL_WIDTH - 1),
		10911 => to_unsigned(28359, LUT_AMPL_WIDTH - 1),
		10912 => to_unsigned(28360, LUT_AMPL_WIDTH - 1),
		10913 => to_unsigned(28362, LUT_AMPL_WIDTH - 1),
		10914 => to_unsigned(28363, LUT_AMPL_WIDTH - 1),
		10915 => to_unsigned(28365, LUT_AMPL_WIDTH - 1),
		10916 => to_unsigned(28367, LUT_AMPL_WIDTH - 1),
		10917 => to_unsigned(28368, LUT_AMPL_WIDTH - 1),
		10918 => to_unsigned(28370, LUT_AMPL_WIDTH - 1),
		10919 => to_unsigned(28371, LUT_AMPL_WIDTH - 1),
		10920 => to_unsigned(28373, LUT_AMPL_WIDTH - 1),
		10921 => to_unsigned(28374, LUT_AMPL_WIDTH - 1),
		10922 => to_unsigned(28376, LUT_AMPL_WIDTH - 1),
		10923 => to_unsigned(28378, LUT_AMPL_WIDTH - 1),
		10924 => to_unsigned(28379, LUT_AMPL_WIDTH - 1),
		10925 => to_unsigned(28381, LUT_AMPL_WIDTH - 1),
		10926 => to_unsigned(28382, LUT_AMPL_WIDTH - 1),
		10927 => to_unsigned(28384, LUT_AMPL_WIDTH - 1),
		10928 => to_unsigned(28385, LUT_AMPL_WIDTH - 1),
		10929 => to_unsigned(28387, LUT_AMPL_WIDTH - 1),
		10930 => to_unsigned(28389, LUT_AMPL_WIDTH - 1),
		10931 => to_unsigned(28390, LUT_AMPL_WIDTH - 1),
		10932 => to_unsigned(28392, LUT_AMPL_WIDTH - 1),
		10933 => to_unsigned(28393, LUT_AMPL_WIDTH - 1),
		10934 => to_unsigned(28395, LUT_AMPL_WIDTH - 1),
		10935 => to_unsigned(28396, LUT_AMPL_WIDTH - 1),
		10936 => to_unsigned(28398, LUT_AMPL_WIDTH - 1),
		10937 => to_unsigned(28400, LUT_AMPL_WIDTH - 1),
		10938 => to_unsigned(28401, LUT_AMPL_WIDTH - 1),
		10939 => to_unsigned(28403, LUT_AMPL_WIDTH - 1),
		10940 => to_unsigned(28404, LUT_AMPL_WIDTH - 1),
		10941 => to_unsigned(28406, LUT_AMPL_WIDTH - 1),
		10942 => to_unsigned(28407, LUT_AMPL_WIDTH - 1),
		10943 => to_unsigned(28409, LUT_AMPL_WIDTH - 1),
		10944 => to_unsigned(28411, LUT_AMPL_WIDTH - 1),
		10945 => to_unsigned(28412, LUT_AMPL_WIDTH - 1),
		10946 => to_unsigned(28414, LUT_AMPL_WIDTH - 1),
		10947 => to_unsigned(28415, LUT_AMPL_WIDTH - 1),
		10948 => to_unsigned(28417, LUT_AMPL_WIDTH - 1),
		10949 => to_unsigned(28418, LUT_AMPL_WIDTH - 1),
		10950 => to_unsigned(28420, LUT_AMPL_WIDTH - 1),
		10951 => to_unsigned(28421, LUT_AMPL_WIDTH - 1),
		10952 => to_unsigned(28423, LUT_AMPL_WIDTH - 1),
		10953 => to_unsigned(28425, LUT_AMPL_WIDTH - 1),
		10954 => to_unsigned(28426, LUT_AMPL_WIDTH - 1),
		10955 => to_unsigned(28428, LUT_AMPL_WIDTH - 1),
		10956 => to_unsigned(28429, LUT_AMPL_WIDTH - 1),
		10957 => to_unsigned(28431, LUT_AMPL_WIDTH - 1),
		10958 => to_unsigned(28432, LUT_AMPL_WIDTH - 1),
		10959 => to_unsigned(28434, LUT_AMPL_WIDTH - 1),
		10960 => to_unsigned(28436, LUT_AMPL_WIDTH - 1),
		10961 => to_unsigned(28437, LUT_AMPL_WIDTH - 1),
		10962 => to_unsigned(28439, LUT_AMPL_WIDTH - 1),
		10963 => to_unsigned(28440, LUT_AMPL_WIDTH - 1),
		10964 => to_unsigned(28442, LUT_AMPL_WIDTH - 1),
		10965 => to_unsigned(28443, LUT_AMPL_WIDTH - 1),
		10966 => to_unsigned(28445, LUT_AMPL_WIDTH - 1),
		10967 => to_unsigned(28446, LUT_AMPL_WIDTH - 1),
		10968 => to_unsigned(28448, LUT_AMPL_WIDTH - 1),
		10969 => to_unsigned(28450, LUT_AMPL_WIDTH - 1),
		10970 => to_unsigned(28451, LUT_AMPL_WIDTH - 1),
		10971 => to_unsigned(28453, LUT_AMPL_WIDTH - 1),
		10972 => to_unsigned(28454, LUT_AMPL_WIDTH - 1),
		10973 => to_unsigned(28456, LUT_AMPL_WIDTH - 1),
		10974 => to_unsigned(28457, LUT_AMPL_WIDTH - 1),
		10975 => to_unsigned(28459, LUT_AMPL_WIDTH - 1),
		10976 => to_unsigned(28460, LUT_AMPL_WIDTH - 1),
		10977 => to_unsigned(28462, LUT_AMPL_WIDTH - 1),
		10978 => to_unsigned(28464, LUT_AMPL_WIDTH - 1),
		10979 => to_unsigned(28465, LUT_AMPL_WIDTH - 1),
		10980 => to_unsigned(28467, LUT_AMPL_WIDTH - 1),
		10981 => to_unsigned(28468, LUT_AMPL_WIDTH - 1),
		10982 => to_unsigned(28470, LUT_AMPL_WIDTH - 1),
		10983 => to_unsigned(28471, LUT_AMPL_WIDTH - 1),
		10984 => to_unsigned(28473, LUT_AMPL_WIDTH - 1),
		10985 => to_unsigned(28474, LUT_AMPL_WIDTH - 1),
		10986 => to_unsigned(28476, LUT_AMPL_WIDTH - 1),
		10987 => to_unsigned(28478, LUT_AMPL_WIDTH - 1),
		10988 => to_unsigned(28479, LUT_AMPL_WIDTH - 1),
		10989 => to_unsigned(28481, LUT_AMPL_WIDTH - 1),
		10990 => to_unsigned(28482, LUT_AMPL_WIDTH - 1),
		10991 => to_unsigned(28484, LUT_AMPL_WIDTH - 1),
		10992 => to_unsigned(28485, LUT_AMPL_WIDTH - 1),
		10993 => to_unsigned(28487, LUT_AMPL_WIDTH - 1),
		10994 => to_unsigned(28488, LUT_AMPL_WIDTH - 1),
		10995 => to_unsigned(28490, LUT_AMPL_WIDTH - 1),
		10996 => to_unsigned(28492, LUT_AMPL_WIDTH - 1),
		10997 => to_unsigned(28493, LUT_AMPL_WIDTH - 1),
		10998 => to_unsigned(28495, LUT_AMPL_WIDTH - 1),
		10999 => to_unsigned(28496, LUT_AMPL_WIDTH - 1),
		11000 => to_unsigned(28498, LUT_AMPL_WIDTH - 1),
		11001 => to_unsigned(28499, LUT_AMPL_WIDTH - 1),
		11002 => to_unsigned(28501, LUT_AMPL_WIDTH - 1),
		11003 => to_unsigned(28502, LUT_AMPL_WIDTH - 1),
		11004 => to_unsigned(28504, LUT_AMPL_WIDTH - 1),
		11005 => to_unsigned(28505, LUT_AMPL_WIDTH - 1),
		11006 => to_unsigned(28507, LUT_AMPL_WIDTH - 1),
		11007 => to_unsigned(28509, LUT_AMPL_WIDTH - 1),
		11008 => to_unsigned(28510, LUT_AMPL_WIDTH - 1),
		11009 => to_unsigned(28512, LUT_AMPL_WIDTH - 1),
		11010 => to_unsigned(28513, LUT_AMPL_WIDTH - 1),
		11011 => to_unsigned(28515, LUT_AMPL_WIDTH - 1),
		11012 => to_unsigned(28516, LUT_AMPL_WIDTH - 1),
		11013 => to_unsigned(28518, LUT_AMPL_WIDTH - 1),
		11014 => to_unsigned(28519, LUT_AMPL_WIDTH - 1),
		11015 => to_unsigned(28521, LUT_AMPL_WIDTH - 1),
		11016 => to_unsigned(28523, LUT_AMPL_WIDTH - 1),
		11017 => to_unsigned(28524, LUT_AMPL_WIDTH - 1),
		11018 => to_unsigned(28526, LUT_AMPL_WIDTH - 1),
		11019 => to_unsigned(28527, LUT_AMPL_WIDTH - 1),
		11020 => to_unsigned(28529, LUT_AMPL_WIDTH - 1),
		11021 => to_unsigned(28530, LUT_AMPL_WIDTH - 1),
		11022 => to_unsigned(28532, LUT_AMPL_WIDTH - 1),
		11023 => to_unsigned(28533, LUT_AMPL_WIDTH - 1),
		11024 => to_unsigned(28535, LUT_AMPL_WIDTH - 1),
		11025 => to_unsigned(28536, LUT_AMPL_WIDTH - 1),
		11026 => to_unsigned(28538, LUT_AMPL_WIDTH - 1),
		11027 => to_unsigned(28540, LUT_AMPL_WIDTH - 1),
		11028 => to_unsigned(28541, LUT_AMPL_WIDTH - 1),
		11029 => to_unsigned(28543, LUT_AMPL_WIDTH - 1),
		11030 => to_unsigned(28544, LUT_AMPL_WIDTH - 1),
		11031 => to_unsigned(28546, LUT_AMPL_WIDTH - 1),
		11032 => to_unsigned(28547, LUT_AMPL_WIDTH - 1),
		11033 => to_unsigned(28549, LUT_AMPL_WIDTH - 1),
		11034 => to_unsigned(28550, LUT_AMPL_WIDTH - 1),
		11035 => to_unsigned(28552, LUT_AMPL_WIDTH - 1),
		11036 => to_unsigned(28553, LUT_AMPL_WIDTH - 1),
		11037 => to_unsigned(28555, LUT_AMPL_WIDTH - 1),
		11038 => to_unsigned(28556, LUT_AMPL_WIDTH - 1),
		11039 => to_unsigned(28558, LUT_AMPL_WIDTH - 1),
		11040 => to_unsigned(28560, LUT_AMPL_WIDTH - 1),
		11041 => to_unsigned(28561, LUT_AMPL_WIDTH - 1),
		11042 => to_unsigned(28563, LUT_AMPL_WIDTH - 1),
		11043 => to_unsigned(28564, LUT_AMPL_WIDTH - 1),
		11044 => to_unsigned(28566, LUT_AMPL_WIDTH - 1),
		11045 => to_unsigned(28567, LUT_AMPL_WIDTH - 1),
		11046 => to_unsigned(28569, LUT_AMPL_WIDTH - 1),
		11047 => to_unsigned(28570, LUT_AMPL_WIDTH - 1),
		11048 => to_unsigned(28572, LUT_AMPL_WIDTH - 1),
		11049 => to_unsigned(28573, LUT_AMPL_WIDTH - 1),
		11050 => to_unsigned(28575, LUT_AMPL_WIDTH - 1),
		11051 => to_unsigned(28576, LUT_AMPL_WIDTH - 1),
		11052 => to_unsigned(28578, LUT_AMPL_WIDTH - 1),
		11053 => to_unsigned(28580, LUT_AMPL_WIDTH - 1),
		11054 => to_unsigned(28581, LUT_AMPL_WIDTH - 1),
		11055 => to_unsigned(28583, LUT_AMPL_WIDTH - 1),
		11056 => to_unsigned(28584, LUT_AMPL_WIDTH - 1),
		11057 => to_unsigned(28586, LUT_AMPL_WIDTH - 1),
		11058 => to_unsigned(28587, LUT_AMPL_WIDTH - 1),
		11059 => to_unsigned(28589, LUT_AMPL_WIDTH - 1),
		11060 => to_unsigned(28590, LUT_AMPL_WIDTH - 1),
		11061 => to_unsigned(28592, LUT_AMPL_WIDTH - 1),
		11062 => to_unsigned(28593, LUT_AMPL_WIDTH - 1),
		11063 => to_unsigned(28595, LUT_AMPL_WIDTH - 1),
		11064 => to_unsigned(28596, LUT_AMPL_WIDTH - 1),
		11065 => to_unsigned(28598, LUT_AMPL_WIDTH - 1),
		11066 => to_unsigned(28600, LUT_AMPL_WIDTH - 1),
		11067 => to_unsigned(28601, LUT_AMPL_WIDTH - 1),
		11068 => to_unsigned(28603, LUT_AMPL_WIDTH - 1),
		11069 => to_unsigned(28604, LUT_AMPL_WIDTH - 1),
		11070 => to_unsigned(28606, LUT_AMPL_WIDTH - 1),
		11071 => to_unsigned(28607, LUT_AMPL_WIDTH - 1),
		11072 => to_unsigned(28609, LUT_AMPL_WIDTH - 1),
		11073 => to_unsigned(28610, LUT_AMPL_WIDTH - 1),
		11074 => to_unsigned(28612, LUT_AMPL_WIDTH - 1),
		11075 => to_unsigned(28613, LUT_AMPL_WIDTH - 1),
		11076 => to_unsigned(28615, LUT_AMPL_WIDTH - 1),
		11077 => to_unsigned(28616, LUT_AMPL_WIDTH - 1),
		11078 => to_unsigned(28618, LUT_AMPL_WIDTH - 1),
		11079 => to_unsigned(28619, LUT_AMPL_WIDTH - 1),
		11080 => to_unsigned(28621, LUT_AMPL_WIDTH - 1),
		11081 => to_unsigned(28622, LUT_AMPL_WIDTH - 1),
		11082 => to_unsigned(28624, LUT_AMPL_WIDTH - 1),
		11083 => to_unsigned(28626, LUT_AMPL_WIDTH - 1),
		11084 => to_unsigned(28627, LUT_AMPL_WIDTH - 1),
		11085 => to_unsigned(28629, LUT_AMPL_WIDTH - 1),
		11086 => to_unsigned(28630, LUT_AMPL_WIDTH - 1),
		11087 => to_unsigned(28632, LUT_AMPL_WIDTH - 1),
		11088 => to_unsigned(28633, LUT_AMPL_WIDTH - 1),
		11089 => to_unsigned(28635, LUT_AMPL_WIDTH - 1),
		11090 => to_unsigned(28636, LUT_AMPL_WIDTH - 1),
		11091 => to_unsigned(28638, LUT_AMPL_WIDTH - 1),
		11092 => to_unsigned(28639, LUT_AMPL_WIDTH - 1),
		11093 => to_unsigned(28641, LUT_AMPL_WIDTH - 1),
		11094 => to_unsigned(28642, LUT_AMPL_WIDTH - 1),
		11095 => to_unsigned(28644, LUT_AMPL_WIDTH - 1),
		11096 => to_unsigned(28645, LUT_AMPL_WIDTH - 1),
		11097 => to_unsigned(28647, LUT_AMPL_WIDTH - 1),
		11098 => to_unsigned(28648, LUT_AMPL_WIDTH - 1),
		11099 => to_unsigned(28650, LUT_AMPL_WIDTH - 1),
		11100 => to_unsigned(28651, LUT_AMPL_WIDTH - 1),
		11101 => to_unsigned(28653, LUT_AMPL_WIDTH - 1),
		11102 => to_unsigned(28655, LUT_AMPL_WIDTH - 1),
		11103 => to_unsigned(28656, LUT_AMPL_WIDTH - 1),
		11104 => to_unsigned(28658, LUT_AMPL_WIDTH - 1),
		11105 => to_unsigned(28659, LUT_AMPL_WIDTH - 1),
		11106 => to_unsigned(28661, LUT_AMPL_WIDTH - 1),
		11107 => to_unsigned(28662, LUT_AMPL_WIDTH - 1),
		11108 => to_unsigned(28664, LUT_AMPL_WIDTH - 1),
		11109 => to_unsigned(28665, LUT_AMPL_WIDTH - 1),
		11110 => to_unsigned(28667, LUT_AMPL_WIDTH - 1),
		11111 => to_unsigned(28668, LUT_AMPL_WIDTH - 1),
		11112 => to_unsigned(28670, LUT_AMPL_WIDTH - 1),
		11113 => to_unsigned(28671, LUT_AMPL_WIDTH - 1),
		11114 => to_unsigned(28673, LUT_AMPL_WIDTH - 1),
		11115 => to_unsigned(28674, LUT_AMPL_WIDTH - 1),
		11116 => to_unsigned(28676, LUT_AMPL_WIDTH - 1),
		11117 => to_unsigned(28677, LUT_AMPL_WIDTH - 1),
		11118 => to_unsigned(28679, LUT_AMPL_WIDTH - 1),
		11119 => to_unsigned(28680, LUT_AMPL_WIDTH - 1),
		11120 => to_unsigned(28682, LUT_AMPL_WIDTH - 1),
		11121 => to_unsigned(28683, LUT_AMPL_WIDTH - 1),
		11122 => to_unsigned(28685, LUT_AMPL_WIDTH - 1),
		11123 => to_unsigned(28686, LUT_AMPL_WIDTH - 1),
		11124 => to_unsigned(28688, LUT_AMPL_WIDTH - 1),
		11125 => to_unsigned(28690, LUT_AMPL_WIDTH - 1),
		11126 => to_unsigned(28691, LUT_AMPL_WIDTH - 1),
		11127 => to_unsigned(28693, LUT_AMPL_WIDTH - 1),
		11128 => to_unsigned(28694, LUT_AMPL_WIDTH - 1),
		11129 => to_unsigned(28696, LUT_AMPL_WIDTH - 1),
		11130 => to_unsigned(28697, LUT_AMPL_WIDTH - 1),
		11131 => to_unsigned(28699, LUT_AMPL_WIDTH - 1),
		11132 => to_unsigned(28700, LUT_AMPL_WIDTH - 1),
		11133 => to_unsigned(28702, LUT_AMPL_WIDTH - 1),
		11134 => to_unsigned(28703, LUT_AMPL_WIDTH - 1),
		11135 => to_unsigned(28705, LUT_AMPL_WIDTH - 1),
		11136 => to_unsigned(28706, LUT_AMPL_WIDTH - 1),
		11137 => to_unsigned(28708, LUT_AMPL_WIDTH - 1),
		11138 => to_unsigned(28709, LUT_AMPL_WIDTH - 1),
		11139 => to_unsigned(28711, LUT_AMPL_WIDTH - 1),
		11140 => to_unsigned(28712, LUT_AMPL_WIDTH - 1),
		11141 => to_unsigned(28714, LUT_AMPL_WIDTH - 1),
		11142 => to_unsigned(28715, LUT_AMPL_WIDTH - 1),
		11143 => to_unsigned(28717, LUT_AMPL_WIDTH - 1),
		11144 => to_unsigned(28718, LUT_AMPL_WIDTH - 1),
		11145 => to_unsigned(28720, LUT_AMPL_WIDTH - 1),
		11146 => to_unsigned(28721, LUT_AMPL_WIDTH - 1),
		11147 => to_unsigned(28723, LUT_AMPL_WIDTH - 1),
		11148 => to_unsigned(28724, LUT_AMPL_WIDTH - 1),
		11149 => to_unsigned(28726, LUT_AMPL_WIDTH - 1),
		11150 => to_unsigned(28727, LUT_AMPL_WIDTH - 1),
		11151 => to_unsigned(28729, LUT_AMPL_WIDTH - 1),
		11152 => to_unsigned(28730, LUT_AMPL_WIDTH - 1),
		11153 => to_unsigned(28732, LUT_AMPL_WIDTH - 1),
		11154 => to_unsigned(28733, LUT_AMPL_WIDTH - 1),
		11155 => to_unsigned(28735, LUT_AMPL_WIDTH - 1),
		11156 => to_unsigned(28736, LUT_AMPL_WIDTH - 1),
		11157 => to_unsigned(28738, LUT_AMPL_WIDTH - 1),
		11158 => to_unsigned(28739, LUT_AMPL_WIDTH - 1),
		11159 => to_unsigned(28741, LUT_AMPL_WIDTH - 1),
		11160 => to_unsigned(28742, LUT_AMPL_WIDTH - 1),
		11161 => to_unsigned(28744, LUT_AMPL_WIDTH - 1),
		11162 => to_unsigned(28745, LUT_AMPL_WIDTH - 1),
		11163 => to_unsigned(28747, LUT_AMPL_WIDTH - 1),
		11164 => to_unsigned(28748, LUT_AMPL_WIDTH - 1),
		11165 => to_unsigned(28750, LUT_AMPL_WIDTH - 1),
		11166 => to_unsigned(28752, LUT_AMPL_WIDTH - 1),
		11167 => to_unsigned(28753, LUT_AMPL_WIDTH - 1),
		11168 => to_unsigned(28755, LUT_AMPL_WIDTH - 1),
		11169 => to_unsigned(28756, LUT_AMPL_WIDTH - 1),
		11170 => to_unsigned(28758, LUT_AMPL_WIDTH - 1),
		11171 => to_unsigned(28759, LUT_AMPL_WIDTH - 1),
		11172 => to_unsigned(28761, LUT_AMPL_WIDTH - 1),
		11173 => to_unsigned(28762, LUT_AMPL_WIDTH - 1),
		11174 => to_unsigned(28764, LUT_AMPL_WIDTH - 1),
		11175 => to_unsigned(28765, LUT_AMPL_WIDTH - 1),
		11176 => to_unsigned(28767, LUT_AMPL_WIDTH - 1),
		11177 => to_unsigned(28768, LUT_AMPL_WIDTH - 1),
		11178 => to_unsigned(28770, LUT_AMPL_WIDTH - 1),
		11179 => to_unsigned(28771, LUT_AMPL_WIDTH - 1),
		11180 => to_unsigned(28773, LUT_AMPL_WIDTH - 1),
		11181 => to_unsigned(28774, LUT_AMPL_WIDTH - 1),
		11182 => to_unsigned(28776, LUT_AMPL_WIDTH - 1),
		11183 => to_unsigned(28777, LUT_AMPL_WIDTH - 1),
		11184 => to_unsigned(28779, LUT_AMPL_WIDTH - 1),
		11185 => to_unsigned(28780, LUT_AMPL_WIDTH - 1),
		11186 => to_unsigned(28782, LUT_AMPL_WIDTH - 1),
		11187 => to_unsigned(28783, LUT_AMPL_WIDTH - 1),
		11188 => to_unsigned(28785, LUT_AMPL_WIDTH - 1),
		11189 => to_unsigned(28786, LUT_AMPL_WIDTH - 1),
		11190 => to_unsigned(28788, LUT_AMPL_WIDTH - 1),
		11191 => to_unsigned(28789, LUT_AMPL_WIDTH - 1),
		11192 => to_unsigned(28791, LUT_AMPL_WIDTH - 1),
		11193 => to_unsigned(28792, LUT_AMPL_WIDTH - 1),
		11194 => to_unsigned(28794, LUT_AMPL_WIDTH - 1),
		11195 => to_unsigned(28795, LUT_AMPL_WIDTH - 1),
		11196 => to_unsigned(28797, LUT_AMPL_WIDTH - 1),
		11197 => to_unsigned(28798, LUT_AMPL_WIDTH - 1),
		11198 => to_unsigned(28800, LUT_AMPL_WIDTH - 1),
		11199 => to_unsigned(28801, LUT_AMPL_WIDTH - 1),
		11200 => to_unsigned(28803, LUT_AMPL_WIDTH - 1),
		11201 => to_unsigned(28804, LUT_AMPL_WIDTH - 1),
		11202 => to_unsigned(28806, LUT_AMPL_WIDTH - 1),
		11203 => to_unsigned(28807, LUT_AMPL_WIDTH - 1),
		11204 => to_unsigned(28809, LUT_AMPL_WIDTH - 1),
		11205 => to_unsigned(28810, LUT_AMPL_WIDTH - 1),
		11206 => to_unsigned(28812, LUT_AMPL_WIDTH - 1),
		11207 => to_unsigned(28813, LUT_AMPL_WIDTH - 1),
		11208 => to_unsigned(28815, LUT_AMPL_WIDTH - 1),
		11209 => to_unsigned(28816, LUT_AMPL_WIDTH - 1),
		11210 => to_unsigned(28818, LUT_AMPL_WIDTH - 1),
		11211 => to_unsigned(28819, LUT_AMPL_WIDTH - 1),
		11212 => to_unsigned(28821, LUT_AMPL_WIDTH - 1),
		11213 => to_unsigned(28822, LUT_AMPL_WIDTH - 1),
		11214 => to_unsigned(28824, LUT_AMPL_WIDTH - 1),
		11215 => to_unsigned(28825, LUT_AMPL_WIDTH - 1),
		11216 => to_unsigned(28827, LUT_AMPL_WIDTH - 1),
		11217 => to_unsigned(28828, LUT_AMPL_WIDTH - 1),
		11218 => to_unsigned(28830, LUT_AMPL_WIDTH - 1),
		11219 => to_unsigned(28831, LUT_AMPL_WIDTH - 1),
		11220 => to_unsigned(28832, LUT_AMPL_WIDTH - 1),
		11221 => to_unsigned(28834, LUT_AMPL_WIDTH - 1),
		11222 => to_unsigned(28835, LUT_AMPL_WIDTH - 1),
		11223 => to_unsigned(28837, LUT_AMPL_WIDTH - 1),
		11224 => to_unsigned(28838, LUT_AMPL_WIDTH - 1),
		11225 => to_unsigned(28840, LUT_AMPL_WIDTH - 1),
		11226 => to_unsigned(28841, LUT_AMPL_WIDTH - 1),
		11227 => to_unsigned(28843, LUT_AMPL_WIDTH - 1),
		11228 => to_unsigned(28844, LUT_AMPL_WIDTH - 1),
		11229 => to_unsigned(28846, LUT_AMPL_WIDTH - 1),
		11230 => to_unsigned(28847, LUT_AMPL_WIDTH - 1),
		11231 => to_unsigned(28849, LUT_AMPL_WIDTH - 1),
		11232 => to_unsigned(28850, LUT_AMPL_WIDTH - 1),
		11233 => to_unsigned(28852, LUT_AMPL_WIDTH - 1),
		11234 => to_unsigned(28853, LUT_AMPL_WIDTH - 1),
		11235 => to_unsigned(28855, LUT_AMPL_WIDTH - 1),
		11236 => to_unsigned(28856, LUT_AMPL_WIDTH - 1),
		11237 => to_unsigned(28858, LUT_AMPL_WIDTH - 1),
		11238 => to_unsigned(28859, LUT_AMPL_WIDTH - 1),
		11239 => to_unsigned(28861, LUT_AMPL_WIDTH - 1),
		11240 => to_unsigned(28862, LUT_AMPL_WIDTH - 1),
		11241 => to_unsigned(28864, LUT_AMPL_WIDTH - 1),
		11242 => to_unsigned(28865, LUT_AMPL_WIDTH - 1),
		11243 => to_unsigned(28867, LUT_AMPL_WIDTH - 1),
		11244 => to_unsigned(28868, LUT_AMPL_WIDTH - 1),
		11245 => to_unsigned(28870, LUT_AMPL_WIDTH - 1),
		11246 => to_unsigned(28871, LUT_AMPL_WIDTH - 1),
		11247 => to_unsigned(28873, LUT_AMPL_WIDTH - 1),
		11248 => to_unsigned(28874, LUT_AMPL_WIDTH - 1),
		11249 => to_unsigned(28876, LUT_AMPL_WIDTH - 1),
		11250 => to_unsigned(28877, LUT_AMPL_WIDTH - 1),
		11251 => to_unsigned(28879, LUT_AMPL_WIDTH - 1),
		11252 => to_unsigned(28880, LUT_AMPL_WIDTH - 1),
		11253 => to_unsigned(28882, LUT_AMPL_WIDTH - 1),
		11254 => to_unsigned(28883, LUT_AMPL_WIDTH - 1),
		11255 => to_unsigned(28885, LUT_AMPL_WIDTH - 1),
		11256 => to_unsigned(28886, LUT_AMPL_WIDTH - 1),
		11257 => to_unsigned(28888, LUT_AMPL_WIDTH - 1),
		11258 => to_unsigned(28889, LUT_AMPL_WIDTH - 1),
		11259 => to_unsigned(28891, LUT_AMPL_WIDTH - 1),
		11260 => to_unsigned(28892, LUT_AMPL_WIDTH - 1),
		11261 => to_unsigned(28893, LUT_AMPL_WIDTH - 1),
		11262 => to_unsigned(28895, LUT_AMPL_WIDTH - 1),
		11263 => to_unsigned(28896, LUT_AMPL_WIDTH - 1),
		11264 => to_unsigned(28898, LUT_AMPL_WIDTH - 1),
		11265 => to_unsigned(28899, LUT_AMPL_WIDTH - 1),
		11266 => to_unsigned(28901, LUT_AMPL_WIDTH - 1),
		11267 => to_unsigned(28902, LUT_AMPL_WIDTH - 1),
		11268 => to_unsigned(28904, LUT_AMPL_WIDTH - 1),
		11269 => to_unsigned(28905, LUT_AMPL_WIDTH - 1),
		11270 => to_unsigned(28907, LUT_AMPL_WIDTH - 1),
		11271 => to_unsigned(28908, LUT_AMPL_WIDTH - 1),
		11272 => to_unsigned(28910, LUT_AMPL_WIDTH - 1),
		11273 => to_unsigned(28911, LUT_AMPL_WIDTH - 1),
		11274 => to_unsigned(28913, LUT_AMPL_WIDTH - 1),
		11275 => to_unsigned(28914, LUT_AMPL_WIDTH - 1),
		11276 => to_unsigned(28916, LUT_AMPL_WIDTH - 1),
		11277 => to_unsigned(28917, LUT_AMPL_WIDTH - 1),
		11278 => to_unsigned(28919, LUT_AMPL_WIDTH - 1),
		11279 => to_unsigned(28920, LUT_AMPL_WIDTH - 1),
		11280 => to_unsigned(28922, LUT_AMPL_WIDTH - 1),
		11281 => to_unsigned(28923, LUT_AMPL_WIDTH - 1),
		11282 => to_unsigned(28925, LUT_AMPL_WIDTH - 1),
		11283 => to_unsigned(28926, LUT_AMPL_WIDTH - 1),
		11284 => to_unsigned(28927, LUT_AMPL_WIDTH - 1),
		11285 => to_unsigned(28929, LUT_AMPL_WIDTH - 1),
		11286 => to_unsigned(28930, LUT_AMPL_WIDTH - 1),
		11287 => to_unsigned(28932, LUT_AMPL_WIDTH - 1),
		11288 => to_unsigned(28933, LUT_AMPL_WIDTH - 1),
		11289 => to_unsigned(28935, LUT_AMPL_WIDTH - 1),
		11290 => to_unsigned(28936, LUT_AMPL_WIDTH - 1),
		11291 => to_unsigned(28938, LUT_AMPL_WIDTH - 1),
		11292 => to_unsigned(28939, LUT_AMPL_WIDTH - 1),
		11293 => to_unsigned(28941, LUT_AMPL_WIDTH - 1),
		11294 => to_unsigned(28942, LUT_AMPL_WIDTH - 1),
		11295 => to_unsigned(28944, LUT_AMPL_WIDTH - 1),
		11296 => to_unsigned(28945, LUT_AMPL_WIDTH - 1),
		11297 => to_unsigned(28947, LUT_AMPL_WIDTH - 1),
		11298 => to_unsigned(28948, LUT_AMPL_WIDTH - 1),
		11299 => to_unsigned(28950, LUT_AMPL_WIDTH - 1),
		11300 => to_unsigned(28951, LUT_AMPL_WIDTH - 1),
		11301 => to_unsigned(28953, LUT_AMPL_WIDTH - 1),
		11302 => to_unsigned(28954, LUT_AMPL_WIDTH - 1),
		11303 => to_unsigned(28955, LUT_AMPL_WIDTH - 1),
		11304 => to_unsigned(28957, LUT_AMPL_WIDTH - 1),
		11305 => to_unsigned(28958, LUT_AMPL_WIDTH - 1),
		11306 => to_unsigned(28960, LUT_AMPL_WIDTH - 1),
		11307 => to_unsigned(28961, LUT_AMPL_WIDTH - 1),
		11308 => to_unsigned(28963, LUT_AMPL_WIDTH - 1),
		11309 => to_unsigned(28964, LUT_AMPL_WIDTH - 1),
		11310 => to_unsigned(28966, LUT_AMPL_WIDTH - 1),
		11311 => to_unsigned(28967, LUT_AMPL_WIDTH - 1),
		11312 => to_unsigned(28969, LUT_AMPL_WIDTH - 1),
		11313 => to_unsigned(28970, LUT_AMPL_WIDTH - 1),
		11314 => to_unsigned(28972, LUT_AMPL_WIDTH - 1),
		11315 => to_unsigned(28973, LUT_AMPL_WIDTH - 1),
		11316 => to_unsigned(28975, LUT_AMPL_WIDTH - 1),
		11317 => to_unsigned(28976, LUT_AMPL_WIDTH - 1),
		11318 => to_unsigned(28977, LUT_AMPL_WIDTH - 1),
		11319 => to_unsigned(28979, LUT_AMPL_WIDTH - 1),
		11320 => to_unsigned(28980, LUT_AMPL_WIDTH - 1),
		11321 => to_unsigned(28982, LUT_AMPL_WIDTH - 1),
		11322 => to_unsigned(28983, LUT_AMPL_WIDTH - 1),
		11323 => to_unsigned(28985, LUT_AMPL_WIDTH - 1),
		11324 => to_unsigned(28986, LUT_AMPL_WIDTH - 1),
		11325 => to_unsigned(28988, LUT_AMPL_WIDTH - 1),
		11326 => to_unsigned(28989, LUT_AMPL_WIDTH - 1),
		11327 => to_unsigned(28991, LUT_AMPL_WIDTH - 1),
		11328 => to_unsigned(28992, LUT_AMPL_WIDTH - 1),
		11329 => to_unsigned(28994, LUT_AMPL_WIDTH - 1),
		11330 => to_unsigned(28995, LUT_AMPL_WIDTH - 1),
		11331 => to_unsigned(28997, LUT_AMPL_WIDTH - 1),
		11332 => to_unsigned(28998, LUT_AMPL_WIDTH - 1),
		11333 => to_unsigned(28999, LUT_AMPL_WIDTH - 1),
		11334 => to_unsigned(29001, LUT_AMPL_WIDTH - 1),
		11335 => to_unsigned(29002, LUT_AMPL_WIDTH - 1),
		11336 => to_unsigned(29004, LUT_AMPL_WIDTH - 1),
		11337 => to_unsigned(29005, LUT_AMPL_WIDTH - 1),
		11338 => to_unsigned(29007, LUT_AMPL_WIDTH - 1),
		11339 => to_unsigned(29008, LUT_AMPL_WIDTH - 1),
		11340 => to_unsigned(29010, LUT_AMPL_WIDTH - 1),
		11341 => to_unsigned(29011, LUT_AMPL_WIDTH - 1),
		11342 => to_unsigned(29013, LUT_AMPL_WIDTH - 1),
		11343 => to_unsigned(29014, LUT_AMPL_WIDTH - 1),
		11344 => to_unsigned(29016, LUT_AMPL_WIDTH - 1),
		11345 => to_unsigned(29017, LUT_AMPL_WIDTH - 1),
		11346 => to_unsigned(29018, LUT_AMPL_WIDTH - 1),
		11347 => to_unsigned(29020, LUT_AMPL_WIDTH - 1),
		11348 => to_unsigned(29021, LUT_AMPL_WIDTH - 1),
		11349 => to_unsigned(29023, LUT_AMPL_WIDTH - 1),
		11350 => to_unsigned(29024, LUT_AMPL_WIDTH - 1),
		11351 => to_unsigned(29026, LUT_AMPL_WIDTH - 1),
		11352 => to_unsigned(29027, LUT_AMPL_WIDTH - 1),
		11353 => to_unsigned(29029, LUT_AMPL_WIDTH - 1),
		11354 => to_unsigned(29030, LUT_AMPL_WIDTH - 1),
		11355 => to_unsigned(29032, LUT_AMPL_WIDTH - 1),
		11356 => to_unsigned(29033, LUT_AMPL_WIDTH - 1),
		11357 => to_unsigned(29034, LUT_AMPL_WIDTH - 1),
		11358 => to_unsigned(29036, LUT_AMPL_WIDTH - 1),
		11359 => to_unsigned(29037, LUT_AMPL_WIDTH - 1),
		11360 => to_unsigned(29039, LUT_AMPL_WIDTH - 1),
		11361 => to_unsigned(29040, LUT_AMPL_WIDTH - 1),
		11362 => to_unsigned(29042, LUT_AMPL_WIDTH - 1),
		11363 => to_unsigned(29043, LUT_AMPL_WIDTH - 1),
		11364 => to_unsigned(29045, LUT_AMPL_WIDTH - 1),
		11365 => to_unsigned(29046, LUT_AMPL_WIDTH - 1),
		11366 => to_unsigned(29048, LUT_AMPL_WIDTH - 1),
		11367 => to_unsigned(29049, LUT_AMPL_WIDTH - 1),
		11368 => to_unsigned(29050, LUT_AMPL_WIDTH - 1),
		11369 => to_unsigned(29052, LUT_AMPL_WIDTH - 1),
		11370 => to_unsigned(29053, LUT_AMPL_WIDTH - 1),
		11371 => to_unsigned(29055, LUT_AMPL_WIDTH - 1),
		11372 => to_unsigned(29056, LUT_AMPL_WIDTH - 1),
		11373 => to_unsigned(29058, LUT_AMPL_WIDTH - 1),
		11374 => to_unsigned(29059, LUT_AMPL_WIDTH - 1),
		11375 => to_unsigned(29061, LUT_AMPL_WIDTH - 1),
		11376 => to_unsigned(29062, LUT_AMPL_WIDTH - 1),
		11377 => to_unsigned(29064, LUT_AMPL_WIDTH - 1),
		11378 => to_unsigned(29065, LUT_AMPL_WIDTH - 1),
		11379 => to_unsigned(29066, LUT_AMPL_WIDTH - 1),
		11380 => to_unsigned(29068, LUT_AMPL_WIDTH - 1),
		11381 => to_unsigned(29069, LUT_AMPL_WIDTH - 1),
		11382 => to_unsigned(29071, LUT_AMPL_WIDTH - 1),
		11383 => to_unsigned(29072, LUT_AMPL_WIDTH - 1),
		11384 => to_unsigned(29074, LUT_AMPL_WIDTH - 1),
		11385 => to_unsigned(29075, LUT_AMPL_WIDTH - 1),
		11386 => to_unsigned(29077, LUT_AMPL_WIDTH - 1),
		11387 => to_unsigned(29078, LUT_AMPL_WIDTH - 1),
		11388 => to_unsigned(29079, LUT_AMPL_WIDTH - 1),
		11389 => to_unsigned(29081, LUT_AMPL_WIDTH - 1),
		11390 => to_unsigned(29082, LUT_AMPL_WIDTH - 1),
		11391 => to_unsigned(29084, LUT_AMPL_WIDTH - 1),
		11392 => to_unsigned(29085, LUT_AMPL_WIDTH - 1),
		11393 => to_unsigned(29087, LUT_AMPL_WIDTH - 1),
		11394 => to_unsigned(29088, LUT_AMPL_WIDTH - 1),
		11395 => to_unsigned(29090, LUT_AMPL_WIDTH - 1),
		11396 => to_unsigned(29091, LUT_AMPL_WIDTH - 1),
		11397 => to_unsigned(29093, LUT_AMPL_WIDTH - 1),
		11398 => to_unsigned(29094, LUT_AMPL_WIDTH - 1),
		11399 => to_unsigned(29095, LUT_AMPL_WIDTH - 1),
		11400 => to_unsigned(29097, LUT_AMPL_WIDTH - 1),
		11401 => to_unsigned(29098, LUT_AMPL_WIDTH - 1),
		11402 => to_unsigned(29100, LUT_AMPL_WIDTH - 1),
		11403 => to_unsigned(29101, LUT_AMPL_WIDTH - 1),
		11404 => to_unsigned(29103, LUT_AMPL_WIDTH - 1),
		11405 => to_unsigned(29104, LUT_AMPL_WIDTH - 1),
		11406 => to_unsigned(29106, LUT_AMPL_WIDTH - 1),
		11407 => to_unsigned(29107, LUT_AMPL_WIDTH - 1),
		11408 => to_unsigned(29108, LUT_AMPL_WIDTH - 1),
		11409 => to_unsigned(29110, LUT_AMPL_WIDTH - 1),
		11410 => to_unsigned(29111, LUT_AMPL_WIDTH - 1),
		11411 => to_unsigned(29113, LUT_AMPL_WIDTH - 1),
		11412 => to_unsigned(29114, LUT_AMPL_WIDTH - 1),
		11413 => to_unsigned(29116, LUT_AMPL_WIDTH - 1),
		11414 => to_unsigned(29117, LUT_AMPL_WIDTH - 1),
		11415 => to_unsigned(29118, LUT_AMPL_WIDTH - 1),
		11416 => to_unsigned(29120, LUT_AMPL_WIDTH - 1),
		11417 => to_unsigned(29121, LUT_AMPL_WIDTH - 1),
		11418 => to_unsigned(29123, LUT_AMPL_WIDTH - 1),
		11419 => to_unsigned(29124, LUT_AMPL_WIDTH - 1),
		11420 => to_unsigned(29126, LUT_AMPL_WIDTH - 1),
		11421 => to_unsigned(29127, LUT_AMPL_WIDTH - 1),
		11422 => to_unsigned(29129, LUT_AMPL_WIDTH - 1),
		11423 => to_unsigned(29130, LUT_AMPL_WIDTH - 1),
		11424 => to_unsigned(29131, LUT_AMPL_WIDTH - 1),
		11425 => to_unsigned(29133, LUT_AMPL_WIDTH - 1),
		11426 => to_unsigned(29134, LUT_AMPL_WIDTH - 1),
		11427 => to_unsigned(29136, LUT_AMPL_WIDTH - 1),
		11428 => to_unsigned(29137, LUT_AMPL_WIDTH - 1),
		11429 => to_unsigned(29139, LUT_AMPL_WIDTH - 1),
		11430 => to_unsigned(29140, LUT_AMPL_WIDTH - 1),
		11431 => to_unsigned(29142, LUT_AMPL_WIDTH - 1),
		11432 => to_unsigned(29143, LUT_AMPL_WIDTH - 1),
		11433 => to_unsigned(29144, LUT_AMPL_WIDTH - 1),
		11434 => to_unsigned(29146, LUT_AMPL_WIDTH - 1),
		11435 => to_unsigned(29147, LUT_AMPL_WIDTH - 1),
		11436 => to_unsigned(29149, LUT_AMPL_WIDTH - 1),
		11437 => to_unsigned(29150, LUT_AMPL_WIDTH - 1),
		11438 => to_unsigned(29152, LUT_AMPL_WIDTH - 1),
		11439 => to_unsigned(29153, LUT_AMPL_WIDTH - 1),
		11440 => to_unsigned(29154, LUT_AMPL_WIDTH - 1),
		11441 => to_unsigned(29156, LUT_AMPL_WIDTH - 1),
		11442 => to_unsigned(29157, LUT_AMPL_WIDTH - 1),
		11443 => to_unsigned(29159, LUT_AMPL_WIDTH - 1),
		11444 => to_unsigned(29160, LUT_AMPL_WIDTH - 1),
		11445 => to_unsigned(29162, LUT_AMPL_WIDTH - 1),
		11446 => to_unsigned(29163, LUT_AMPL_WIDTH - 1),
		11447 => to_unsigned(29164, LUT_AMPL_WIDTH - 1),
		11448 => to_unsigned(29166, LUT_AMPL_WIDTH - 1),
		11449 => to_unsigned(29167, LUT_AMPL_WIDTH - 1),
		11450 => to_unsigned(29169, LUT_AMPL_WIDTH - 1),
		11451 => to_unsigned(29170, LUT_AMPL_WIDTH - 1),
		11452 => to_unsigned(29172, LUT_AMPL_WIDTH - 1),
		11453 => to_unsigned(29173, LUT_AMPL_WIDTH - 1),
		11454 => to_unsigned(29174, LUT_AMPL_WIDTH - 1),
		11455 => to_unsigned(29176, LUT_AMPL_WIDTH - 1),
		11456 => to_unsigned(29177, LUT_AMPL_WIDTH - 1),
		11457 => to_unsigned(29179, LUT_AMPL_WIDTH - 1),
		11458 => to_unsigned(29180, LUT_AMPL_WIDTH - 1),
		11459 => to_unsigned(29182, LUT_AMPL_WIDTH - 1),
		11460 => to_unsigned(29183, LUT_AMPL_WIDTH - 1),
		11461 => to_unsigned(29184, LUT_AMPL_WIDTH - 1),
		11462 => to_unsigned(29186, LUT_AMPL_WIDTH - 1),
		11463 => to_unsigned(29187, LUT_AMPL_WIDTH - 1),
		11464 => to_unsigned(29189, LUT_AMPL_WIDTH - 1),
		11465 => to_unsigned(29190, LUT_AMPL_WIDTH - 1),
		11466 => to_unsigned(29192, LUT_AMPL_WIDTH - 1),
		11467 => to_unsigned(29193, LUT_AMPL_WIDTH - 1),
		11468 => to_unsigned(29194, LUT_AMPL_WIDTH - 1),
		11469 => to_unsigned(29196, LUT_AMPL_WIDTH - 1),
		11470 => to_unsigned(29197, LUT_AMPL_WIDTH - 1),
		11471 => to_unsigned(29199, LUT_AMPL_WIDTH - 1),
		11472 => to_unsigned(29200, LUT_AMPL_WIDTH - 1),
		11473 => to_unsigned(29202, LUT_AMPL_WIDTH - 1),
		11474 => to_unsigned(29203, LUT_AMPL_WIDTH - 1),
		11475 => to_unsigned(29204, LUT_AMPL_WIDTH - 1),
		11476 => to_unsigned(29206, LUT_AMPL_WIDTH - 1),
		11477 => to_unsigned(29207, LUT_AMPL_WIDTH - 1),
		11478 => to_unsigned(29209, LUT_AMPL_WIDTH - 1),
		11479 => to_unsigned(29210, LUT_AMPL_WIDTH - 1),
		11480 => to_unsigned(29212, LUT_AMPL_WIDTH - 1),
		11481 => to_unsigned(29213, LUT_AMPL_WIDTH - 1),
		11482 => to_unsigned(29214, LUT_AMPL_WIDTH - 1),
		11483 => to_unsigned(29216, LUT_AMPL_WIDTH - 1),
		11484 => to_unsigned(29217, LUT_AMPL_WIDTH - 1),
		11485 => to_unsigned(29219, LUT_AMPL_WIDTH - 1),
		11486 => to_unsigned(29220, LUT_AMPL_WIDTH - 1),
		11487 => to_unsigned(29222, LUT_AMPL_WIDTH - 1),
		11488 => to_unsigned(29223, LUT_AMPL_WIDTH - 1),
		11489 => to_unsigned(29224, LUT_AMPL_WIDTH - 1),
		11490 => to_unsigned(29226, LUT_AMPL_WIDTH - 1),
		11491 => to_unsigned(29227, LUT_AMPL_WIDTH - 1),
		11492 => to_unsigned(29229, LUT_AMPL_WIDTH - 1),
		11493 => to_unsigned(29230, LUT_AMPL_WIDTH - 1),
		11494 => to_unsigned(29231, LUT_AMPL_WIDTH - 1),
		11495 => to_unsigned(29233, LUT_AMPL_WIDTH - 1),
		11496 => to_unsigned(29234, LUT_AMPL_WIDTH - 1),
		11497 => to_unsigned(29236, LUT_AMPL_WIDTH - 1),
		11498 => to_unsigned(29237, LUT_AMPL_WIDTH - 1),
		11499 => to_unsigned(29239, LUT_AMPL_WIDTH - 1),
		11500 => to_unsigned(29240, LUT_AMPL_WIDTH - 1),
		11501 => to_unsigned(29241, LUT_AMPL_WIDTH - 1),
		11502 => to_unsigned(29243, LUT_AMPL_WIDTH - 1),
		11503 => to_unsigned(29244, LUT_AMPL_WIDTH - 1),
		11504 => to_unsigned(29246, LUT_AMPL_WIDTH - 1),
		11505 => to_unsigned(29247, LUT_AMPL_WIDTH - 1),
		11506 => to_unsigned(29248, LUT_AMPL_WIDTH - 1),
		11507 => to_unsigned(29250, LUT_AMPL_WIDTH - 1),
		11508 => to_unsigned(29251, LUT_AMPL_WIDTH - 1),
		11509 => to_unsigned(29253, LUT_AMPL_WIDTH - 1),
		11510 => to_unsigned(29254, LUT_AMPL_WIDTH - 1),
		11511 => to_unsigned(29256, LUT_AMPL_WIDTH - 1),
		11512 => to_unsigned(29257, LUT_AMPL_WIDTH - 1),
		11513 => to_unsigned(29258, LUT_AMPL_WIDTH - 1),
		11514 => to_unsigned(29260, LUT_AMPL_WIDTH - 1),
		11515 => to_unsigned(29261, LUT_AMPL_WIDTH - 1),
		11516 => to_unsigned(29263, LUT_AMPL_WIDTH - 1),
		11517 => to_unsigned(29264, LUT_AMPL_WIDTH - 1),
		11518 => to_unsigned(29265, LUT_AMPL_WIDTH - 1),
		11519 => to_unsigned(29267, LUT_AMPL_WIDTH - 1),
		11520 => to_unsigned(29268, LUT_AMPL_WIDTH - 1),
		11521 => to_unsigned(29270, LUT_AMPL_WIDTH - 1),
		11522 => to_unsigned(29271, LUT_AMPL_WIDTH - 1),
		11523 => to_unsigned(29273, LUT_AMPL_WIDTH - 1),
		11524 => to_unsigned(29274, LUT_AMPL_WIDTH - 1),
		11525 => to_unsigned(29275, LUT_AMPL_WIDTH - 1),
		11526 => to_unsigned(29277, LUT_AMPL_WIDTH - 1),
		11527 => to_unsigned(29278, LUT_AMPL_WIDTH - 1),
		11528 => to_unsigned(29280, LUT_AMPL_WIDTH - 1),
		11529 => to_unsigned(29281, LUT_AMPL_WIDTH - 1),
		11530 => to_unsigned(29282, LUT_AMPL_WIDTH - 1),
		11531 => to_unsigned(29284, LUT_AMPL_WIDTH - 1),
		11532 => to_unsigned(29285, LUT_AMPL_WIDTH - 1),
		11533 => to_unsigned(29287, LUT_AMPL_WIDTH - 1),
		11534 => to_unsigned(29288, LUT_AMPL_WIDTH - 1),
		11535 => to_unsigned(29289, LUT_AMPL_WIDTH - 1),
		11536 => to_unsigned(29291, LUT_AMPL_WIDTH - 1),
		11537 => to_unsigned(29292, LUT_AMPL_WIDTH - 1),
		11538 => to_unsigned(29294, LUT_AMPL_WIDTH - 1),
		11539 => to_unsigned(29295, LUT_AMPL_WIDTH - 1),
		11540 => to_unsigned(29296, LUT_AMPL_WIDTH - 1),
		11541 => to_unsigned(29298, LUT_AMPL_WIDTH - 1),
		11542 => to_unsigned(29299, LUT_AMPL_WIDTH - 1),
		11543 => to_unsigned(29301, LUT_AMPL_WIDTH - 1),
		11544 => to_unsigned(29302, LUT_AMPL_WIDTH - 1),
		11545 => to_unsigned(29304, LUT_AMPL_WIDTH - 1),
		11546 => to_unsigned(29305, LUT_AMPL_WIDTH - 1),
		11547 => to_unsigned(29306, LUT_AMPL_WIDTH - 1),
		11548 => to_unsigned(29308, LUT_AMPL_WIDTH - 1),
		11549 => to_unsigned(29309, LUT_AMPL_WIDTH - 1),
		11550 => to_unsigned(29311, LUT_AMPL_WIDTH - 1),
		11551 => to_unsigned(29312, LUT_AMPL_WIDTH - 1),
		11552 => to_unsigned(29313, LUT_AMPL_WIDTH - 1),
		11553 => to_unsigned(29315, LUT_AMPL_WIDTH - 1),
		11554 => to_unsigned(29316, LUT_AMPL_WIDTH - 1),
		11555 => to_unsigned(29318, LUT_AMPL_WIDTH - 1),
		11556 => to_unsigned(29319, LUT_AMPL_WIDTH - 1),
		11557 => to_unsigned(29320, LUT_AMPL_WIDTH - 1),
		11558 => to_unsigned(29322, LUT_AMPL_WIDTH - 1),
		11559 => to_unsigned(29323, LUT_AMPL_WIDTH - 1),
		11560 => to_unsigned(29325, LUT_AMPL_WIDTH - 1),
		11561 => to_unsigned(29326, LUT_AMPL_WIDTH - 1),
		11562 => to_unsigned(29327, LUT_AMPL_WIDTH - 1),
		11563 => to_unsigned(29329, LUT_AMPL_WIDTH - 1),
		11564 => to_unsigned(29330, LUT_AMPL_WIDTH - 1),
		11565 => to_unsigned(29332, LUT_AMPL_WIDTH - 1),
		11566 => to_unsigned(29333, LUT_AMPL_WIDTH - 1),
		11567 => to_unsigned(29334, LUT_AMPL_WIDTH - 1),
		11568 => to_unsigned(29336, LUT_AMPL_WIDTH - 1),
		11569 => to_unsigned(29337, LUT_AMPL_WIDTH - 1),
		11570 => to_unsigned(29339, LUT_AMPL_WIDTH - 1),
		11571 => to_unsigned(29340, LUT_AMPL_WIDTH - 1),
		11572 => to_unsigned(29341, LUT_AMPL_WIDTH - 1),
		11573 => to_unsigned(29343, LUT_AMPL_WIDTH - 1),
		11574 => to_unsigned(29344, LUT_AMPL_WIDTH - 1),
		11575 => to_unsigned(29346, LUT_AMPL_WIDTH - 1),
		11576 => to_unsigned(29347, LUT_AMPL_WIDTH - 1),
		11577 => to_unsigned(29348, LUT_AMPL_WIDTH - 1),
		11578 => to_unsigned(29350, LUT_AMPL_WIDTH - 1),
		11579 => to_unsigned(29351, LUT_AMPL_WIDTH - 1),
		11580 => to_unsigned(29353, LUT_AMPL_WIDTH - 1),
		11581 => to_unsigned(29354, LUT_AMPL_WIDTH - 1),
		11582 => to_unsigned(29355, LUT_AMPL_WIDTH - 1),
		11583 => to_unsigned(29357, LUT_AMPL_WIDTH - 1),
		11584 => to_unsigned(29358, LUT_AMPL_WIDTH - 1),
		11585 => to_unsigned(29360, LUT_AMPL_WIDTH - 1),
		11586 => to_unsigned(29361, LUT_AMPL_WIDTH - 1),
		11587 => to_unsigned(29362, LUT_AMPL_WIDTH - 1),
		11588 => to_unsigned(29364, LUT_AMPL_WIDTH - 1),
		11589 => to_unsigned(29365, LUT_AMPL_WIDTH - 1),
		11590 => to_unsigned(29366, LUT_AMPL_WIDTH - 1),
		11591 => to_unsigned(29368, LUT_AMPL_WIDTH - 1),
		11592 => to_unsigned(29369, LUT_AMPL_WIDTH - 1),
		11593 => to_unsigned(29371, LUT_AMPL_WIDTH - 1),
		11594 => to_unsigned(29372, LUT_AMPL_WIDTH - 1),
		11595 => to_unsigned(29373, LUT_AMPL_WIDTH - 1),
		11596 => to_unsigned(29375, LUT_AMPL_WIDTH - 1),
		11597 => to_unsigned(29376, LUT_AMPL_WIDTH - 1),
		11598 => to_unsigned(29378, LUT_AMPL_WIDTH - 1),
		11599 => to_unsigned(29379, LUT_AMPL_WIDTH - 1),
		11600 => to_unsigned(29380, LUT_AMPL_WIDTH - 1),
		11601 => to_unsigned(29382, LUT_AMPL_WIDTH - 1),
		11602 => to_unsigned(29383, LUT_AMPL_WIDTH - 1),
		11603 => to_unsigned(29385, LUT_AMPL_WIDTH - 1),
		11604 => to_unsigned(29386, LUT_AMPL_WIDTH - 1),
		11605 => to_unsigned(29387, LUT_AMPL_WIDTH - 1),
		11606 => to_unsigned(29389, LUT_AMPL_WIDTH - 1),
		11607 => to_unsigned(29390, LUT_AMPL_WIDTH - 1),
		11608 => to_unsigned(29392, LUT_AMPL_WIDTH - 1),
		11609 => to_unsigned(29393, LUT_AMPL_WIDTH - 1),
		11610 => to_unsigned(29394, LUT_AMPL_WIDTH - 1),
		11611 => to_unsigned(29396, LUT_AMPL_WIDTH - 1),
		11612 => to_unsigned(29397, LUT_AMPL_WIDTH - 1),
		11613 => to_unsigned(29398, LUT_AMPL_WIDTH - 1),
		11614 => to_unsigned(29400, LUT_AMPL_WIDTH - 1),
		11615 => to_unsigned(29401, LUT_AMPL_WIDTH - 1),
		11616 => to_unsigned(29403, LUT_AMPL_WIDTH - 1),
		11617 => to_unsigned(29404, LUT_AMPL_WIDTH - 1),
		11618 => to_unsigned(29405, LUT_AMPL_WIDTH - 1),
		11619 => to_unsigned(29407, LUT_AMPL_WIDTH - 1),
		11620 => to_unsigned(29408, LUT_AMPL_WIDTH - 1),
		11621 => to_unsigned(29410, LUT_AMPL_WIDTH - 1),
		11622 => to_unsigned(29411, LUT_AMPL_WIDTH - 1),
		11623 => to_unsigned(29412, LUT_AMPL_WIDTH - 1),
		11624 => to_unsigned(29414, LUT_AMPL_WIDTH - 1),
		11625 => to_unsigned(29415, LUT_AMPL_WIDTH - 1),
		11626 => to_unsigned(29416, LUT_AMPL_WIDTH - 1),
		11627 => to_unsigned(29418, LUT_AMPL_WIDTH - 1),
		11628 => to_unsigned(29419, LUT_AMPL_WIDTH - 1),
		11629 => to_unsigned(29421, LUT_AMPL_WIDTH - 1),
		11630 => to_unsigned(29422, LUT_AMPL_WIDTH - 1),
		11631 => to_unsigned(29423, LUT_AMPL_WIDTH - 1),
		11632 => to_unsigned(29425, LUT_AMPL_WIDTH - 1),
		11633 => to_unsigned(29426, LUT_AMPL_WIDTH - 1),
		11634 => to_unsigned(29428, LUT_AMPL_WIDTH - 1),
		11635 => to_unsigned(29429, LUT_AMPL_WIDTH - 1),
		11636 => to_unsigned(29430, LUT_AMPL_WIDTH - 1),
		11637 => to_unsigned(29432, LUT_AMPL_WIDTH - 1),
		11638 => to_unsigned(29433, LUT_AMPL_WIDTH - 1),
		11639 => to_unsigned(29434, LUT_AMPL_WIDTH - 1),
		11640 => to_unsigned(29436, LUT_AMPL_WIDTH - 1),
		11641 => to_unsigned(29437, LUT_AMPL_WIDTH - 1),
		11642 => to_unsigned(29439, LUT_AMPL_WIDTH - 1),
		11643 => to_unsigned(29440, LUT_AMPL_WIDTH - 1),
		11644 => to_unsigned(29441, LUT_AMPL_WIDTH - 1),
		11645 => to_unsigned(29443, LUT_AMPL_WIDTH - 1),
		11646 => to_unsigned(29444, LUT_AMPL_WIDTH - 1),
		11647 => to_unsigned(29445, LUT_AMPL_WIDTH - 1),
		11648 => to_unsigned(29447, LUT_AMPL_WIDTH - 1),
		11649 => to_unsigned(29448, LUT_AMPL_WIDTH - 1),
		11650 => to_unsigned(29450, LUT_AMPL_WIDTH - 1),
		11651 => to_unsigned(29451, LUT_AMPL_WIDTH - 1),
		11652 => to_unsigned(29452, LUT_AMPL_WIDTH - 1),
		11653 => to_unsigned(29454, LUT_AMPL_WIDTH - 1),
		11654 => to_unsigned(29455, LUT_AMPL_WIDTH - 1),
		11655 => to_unsigned(29457, LUT_AMPL_WIDTH - 1),
		11656 => to_unsigned(29458, LUT_AMPL_WIDTH - 1),
		11657 => to_unsigned(29459, LUT_AMPL_WIDTH - 1),
		11658 => to_unsigned(29461, LUT_AMPL_WIDTH - 1),
		11659 => to_unsigned(29462, LUT_AMPL_WIDTH - 1),
		11660 => to_unsigned(29463, LUT_AMPL_WIDTH - 1),
		11661 => to_unsigned(29465, LUT_AMPL_WIDTH - 1),
		11662 => to_unsigned(29466, LUT_AMPL_WIDTH - 1),
		11663 => to_unsigned(29468, LUT_AMPL_WIDTH - 1),
		11664 => to_unsigned(29469, LUT_AMPL_WIDTH - 1),
		11665 => to_unsigned(29470, LUT_AMPL_WIDTH - 1),
		11666 => to_unsigned(29472, LUT_AMPL_WIDTH - 1),
		11667 => to_unsigned(29473, LUT_AMPL_WIDTH - 1),
		11668 => to_unsigned(29474, LUT_AMPL_WIDTH - 1),
		11669 => to_unsigned(29476, LUT_AMPL_WIDTH - 1),
		11670 => to_unsigned(29477, LUT_AMPL_WIDTH - 1),
		11671 => to_unsigned(29478, LUT_AMPL_WIDTH - 1),
		11672 => to_unsigned(29480, LUT_AMPL_WIDTH - 1),
		11673 => to_unsigned(29481, LUT_AMPL_WIDTH - 1),
		11674 => to_unsigned(29483, LUT_AMPL_WIDTH - 1),
		11675 => to_unsigned(29484, LUT_AMPL_WIDTH - 1),
		11676 => to_unsigned(29485, LUT_AMPL_WIDTH - 1),
		11677 => to_unsigned(29487, LUT_AMPL_WIDTH - 1),
		11678 => to_unsigned(29488, LUT_AMPL_WIDTH - 1),
		11679 => to_unsigned(29489, LUT_AMPL_WIDTH - 1),
		11680 => to_unsigned(29491, LUT_AMPL_WIDTH - 1),
		11681 => to_unsigned(29492, LUT_AMPL_WIDTH - 1),
		11682 => to_unsigned(29494, LUT_AMPL_WIDTH - 1),
		11683 => to_unsigned(29495, LUT_AMPL_WIDTH - 1),
		11684 => to_unsigned(29496, LUT_AMPL_WIDTH - 1),
		11685 => to_unsigned(29498, LUT_AMPL_WIDTH - 1),
		11686 => to_unsigned(29499, LUT_AMPL_WIDTH - 1),
		11687 => to_unsigned(29500, LUT_AMPL_WIDTH - 1),
		11688 => to_unsigned(29502, LUT_AMPL_WIDTH - 1),
		11689 => to_unsigned(29503, LUT_AMPL_WIDTH - 1),
		11690 => to_unsigned(29504, LUT_AMPL_WIDTH - 1),
		11691 => to_unsigned(29506, LUT_AMPL_WIDTH - 1),
		11692 => to_unsigned(29507, LUT_AMPL_WIDTH - 1),
		11693 => to_unsigned(29509, LUT_AMPL_WIDTH - 1),
		11694 => to_unsigned(29510, LUT_AMPL_WIDTH - 1),
		11695 => to_unsigned(29511, LUT_AMPL_WIDTH - 1),
		11696 => to_unsigned(29513, LUT_AMPL_WIDTH - 1),
		11697 => to_unsigned(29514, LUT_AMPL_WIDTH - 1),
		11698 => to_unsigned(29515, LUT_AMPL_WIDTH - 1),
		11699 => to_unsigned(29517, LUT_AMPL_WIDTH - 1),
		11700 => to_unsigned(29518, LUT_AMPL_WIDTH - 1),
		11701 => to_unsigned(29520, LUT_AMPL_WIDTH - 1),
		11702 => to_unsigned(29521, LUT_AMPL_WIDTH - 1),
		11703 => to_unsigned(29522, LUT_AMPL_WIDTH - 1),
		11704 => to_unsigned(29524, LUT_AMPL_WIDTH - 1),
		11705 => to_unsigned(29525, LUT_AMPL_WIDTH - 1),
		11706 => to_unsigned(29526, LUT_AMPL_WIDTH - 1),
		11707 => to_unsigned(29528, LUT_AMPL_WIDTH - 1),
		11708 => to_unsigned(29529, LUT_AMPL_WIDTH - 1),
		11709 => to_unsigned(29530, LUT_AMPL_WIDTH - 1),
		11710 => to_unsigned(29532, LUT_AMPL_WIDTH - 1),
		11711 => to_unsigned(29533, LUT_AMPL_WIDTH - 1),
		11712 => to_unsigned(29534, LUT_AMPL_WIDTH - 1),
		11713 => to_unsigned(29536, LUT_AMPL_WIDTH - 1),
		11714 => to_unsigned(29537, LUT_AMPL_WIDTH - 1),
		11715 => to_unsigned(29539, LUT_AMPL_WIDTH - 1),
		11716 => to_unsigned(29540, LUT_AMPL_WIDTH - 1),
		11717 => to_unsigned(29541, LUT_AMPL_WIDTH - 1),
		11718 => to_unsigned(29543, LUT_AMPL_WIDTH - 1),
		11719 => to_unsigned(29544, LUT_AMPL_WIDTH - 1),
		11720 => to_unsigned(29545, LUT_AMPL_WIDTH - 1),
		11721 => to_unsigned(29547, LUT_AMPL_WIDTH - 1),
		11722 => to_unsigned(29548, LUT_AMPL_WIDTH - 1),
		11723 => to_unsigned(29549, LUT_AMPL_WIDTH - 1),
		11724 => to_unsigned(29551, LUT_AMPL_WIDTH - 1),
		11725 => to_unsigned(29552, LUT_AMPL_WIDTH - 1),
		11726 => to_unsigned(29554, LUT_AMPL_WIDTH - 1),
		11727 => to_unsigned(29555, LUT_AMPL_WIDTH - 1),
		11728 => to_unsigned(29556, LUT_AMPL_WIDTH - 1),
		11729 => to_unsigned(29558, LUT_AMPL_WIDTH - 1),
		11730 => to_unsigned(29559, LUT_AMPL_WIDTH - 1),
		11731 => to_unsigned(29560, LUT_AMPL_WIDTH - 1),
		11732 => to_unsigned(29562, LUT_AMPL_WIDTH - 1),
		11733 => to_unsigned(29563, LUT_AMPL_WIDTH - 1),
		11734 => to_unsigned(29564, LUT_AMPL_WIDTH - 1),
		11735 => to_unsigned(29566, LUT_AMPL_WIDTH - 1),
		11736 => to_unsigned(29567, LUT_AMPL_WIDTH - 1),
		11737 => to_unsigned(29568, LUT_AMPL_WIDTH - 1),
		11738 => to_unsigned(29570, LUT_AMPL_WIDTH - 1),
		11739 => to_unsigned(29571, LUT_AMPL_WIDTH - 1),
		11740 => to_unsigned(29572, LUT_AMPL_WIDTH - 1),
		11741 => to_unsigned(29574, LUT_AMPL_WIDTH - 1),
		11742 => to_unsigned(29575, LUT_AMPL_WIDTH - 1),
		11743 => to_unsigned(29577, LUT_AMPL_WIDTH - 1),
		11744 => to_unsigned(29578, LUT_AMPL_WIDTH - 1),
		11745 => to_unsigned(29579, LUT_AMPL_WIDTH - 1),
		11746 => to_unsigned(29581, LUT_AMPL_WIDTH - 1),
		11747 => to_unsigned(29582, LUT_AMPL_WIDTH - 1),
		11748 => to_unsigned(29583, LUT_AMPL_WIDTH - 1),
		11749 => to_unsigned(29585, LUT_AMPL_WIDTH - 1),
		11750 => to_unsigned(29586, LUT_AMPL_WIDTH - 1),
		11751 => to_unsigned(29587, LUT_AMPL_WIDTH - 1),
		11752 => to_unsigned(29589, LUT_AMPL_WIDTH - 1),
		11753 => to_unsigned(29590, LUT_AMPL_WIDTH - 1),
		11754 => to_unsigned(29591, LUT_AMPL_WIDTH - 1),
		11755 => to_unsigned(29593, LUT_AMPL_WIDTH - 1),
		11756 => to_unsigned(29594, LUT_AMPL_WIDTH - 1),
		11757 => to_unsigned(29595, LUT_AMPL_WIDTH - 1),
		11758 => to_unsigned(29597, LUT_AMPL_WIDTH - 1),
		11759 => to_unsigned(29598, LUT_AMPL_WIDTH - 1),
		11760 => to_unsigned(29599, LUT_AMPL_WIDTH - 1),
		11761 => to_unsigned(29601, LUT_AMPL_WIDTH - 1),
		11762 => to_unsigned(29602, LUT_AMPL_WIDTH - 1),
		11763 => to_unsigned(29604, LUT_AMPL_WIDTH - 1),
		11764 => to_unsigned(29605, LUT_AMPL_WIDTH - 1),
		11765 => to_unsigned(29606, LUT_AMPL_WIDTH - 1),
		11766 => to_unsigned(29608, LUT_AMPL_WIDTH - 1),
		11767 => to_unsigned(29609, LUT_AMPL_WIDTH - 1),
		11768 => to_unsigned(29610, LUT_AMPL_WIDTH - 1),
		11769 => to_unsigned(29612, LUT_AMPL_WIDTH - 1),
		11770 => to_unsigned(29613, LUT_AMPL_WIDTH - 1),
		11771 => to_unsigned(29614, LUT_AMPL_WIDTH - 1),
		11772 => to_unsigned(29616, LUT_AMPL_WIDTH - 1),
		11773 => to_unsigned(29617, LUT_AMPL_WIDTH - 1),
		11774 => to_unsigned(29618, LUT_AMPL_WIDTH - 1),
		11775 => to_unsigned(29620, LUT_AMPL_WIDTH - 1),
		11776 => to_unsigned(29621, LUT_AMPL_WIDTH - 1),
		11777 => to_unsigned(29622, LUT_AMPL_WIDTH - 1),
		11778 => to_unsigned(29624, LUT_AMPL_WIDTH - 1),
		11779 => to_unsigned(29625, LUT_AMPL_WIDTH - 1),
		11780 => to_unsigned(29626, LUT_AMPL_WIDTH - 1),
		11781 => to_unsigned(29628, LUT_AMPL_WIDTH - 1),
		11782 => to_unsigned(29629, LUT_AMPL_WIDTH - 1),
		11783 => to_unsigned(29630, LUT_AMPL_WIDTH - 1),
		11784 => to_unsigned(29632, LUT_AMPL_WIDTH - 1),
		11785 => to_unsigned(29633, LUT_AMPL_WIDTH - 1),
		11786 => to_unsigned(29634, LUT_AMPL_WIDTH - 1),
		11787 => to_unsigned(29636, LUT_AMPL_WIDTH - 1),
		11788 => to_unsigned(29637, LUT_AMPL_WIDTH - 1),
		11789 => to_unsigned(29638, LUT_AMPL_WIDTH - 1),
		11790 => to_unsigned(29640, LUT_AMPL_WIDTH - 1),
		11791 => to_unsigned(29641, LUT_AMPL_WIDTH - 1),
		11792 => to_unsigned(29642, LUT_AMPL_WIDTH - 1),
		11793 => to_unsigned(29644, LUT_AMPL_WIDTH - 1),
		11794 => to_unsigned(29645, LUT_AMPL_WIDTH - 1),
		11795 => to_unsigned(29646, LUT_AMPL_WIDTH - 1),
		11796 => to_unsigned(29648, LUT_AMPL_WIDTH - 1),
		11797 => to_unsigned(29649, LUT_AMPL_WIDTH - 1),
		11798 => to_unsigned(29651, LUT_AMPL_WIDTH - 1),
		11799 => to_unsigned(29652, LUT_AMPL_WIDTH - 1),
		11800 => to_unsigned(29653, LUT_AMPL_WIDTH - 1),
		11801 => to_unsigned(29655, LUT_AMPL_WIDTH - 1),
		11802 => to_unsigned(29656, LUT_AMPL_WIDTH - 1),
		11803 => to_unsigned(29657, LUT_AMPL_WIDTH - 1),
		11804 => to_unsigned(29659, LUT_AMPL_WIDTH - 1),
		11805 => to_unsigned(29660, LUT_AMPL_WIDTH - 1),
		11806 => to_unsigned(29661, LUT_AMPL_WIDTH - 1),
		11807 => to_unsigned(29663, LUT_AMPL_WIDTH - 1),
		11808 => to_unsigned(29664, LUT_AMPL_WIDTH - 1),
		11809 => to_unsigned(29665, LUT_AMPL_WIDTH - 1),
		11810 => to_unsigned(29667, LUT_AMPL_WIDTH - 1),
		11811 => to_unsigned(29668, LUT_AMPL_WIDTH - 1),
		11812 => to_unsigned(29669, LUT_AMPL_WIDTH - 1),
		11813 => to_unsigned(29671, LUT_AMPL_WIDTH - 1),
		11814 => to_unsigned(29672, LUT_AMPL_WIDTH - 1),
		11815 => to_unsigned(29673, LUT_AMPL_WIDTH - 1),
		11816 => to_unsigned(29675, LUT_AMPL_WIDTH - 1),
		11817 => to_unsigned(29676, LUT_AMPL_WIDTH - 1),
		11818 => to_unsigned(29677, LUT_AMPL_WIDTH - 1),
		11819 => to_unsigned(29679, LUT_AMPL_WIDTH - 1),
		11820 => to_unsigned(29680, LUT_AMPL_WIDTH - 1),
		11821 => to_unsigned(29681, LUT_AMPL_WIDTH - 1),
		11822 => to_unsigned(29683, LUT_AMPL_WIDTH - 1),
		11823 => to_unsigned(29684, LUT_AMPL_WIDTH - 1),
		11824 => to_unsigned(29685, LUT_AMPL_WIDTH - 1),
		11825 => to_unsigned(29687, LUT_AMPL_WIDTH - 1),
		11826 => to_unsigned(29688, LUT_AMPL_WIDTH - 1),
		11827 => to_unsigned(29689, LUT_AMPL_WIDTH - 1),
		11828 => to_unsigned(29690, LUT_AMPL_WIDTH - 1),
		11829 => to_unsigned(29692, LUT_AMPL_WIDTH - 1),
		11830 => to_unsigned(29693, LUT_AMPL_WIDTH - 1),
		11831 => to_unsigned(29694, LUT_AMPL_WIDTH - 1),
		11832 => to_unsigned(29696, LUT_AMPL_WIDTH - 1),
		11833 => to_unsigned(29697, LUT_AMPL_WIDTH - 1),
		11834 => to_unsigned(29698, LUT_AMPL_WIDTH - 1),
		11835 => to_unsigned(29700, LUT_AMPL_WIDTH - 1),
		11836 => to_unsigned(29701, LUT_AMPL_WIDTH - 1),
		11837 => to_unsigned(29702, LUT_AMPL_WIDTH - 1),
		11838 => to_unsigned(29704, LUT_AMPL_WIDTH - 1),
		11839 => to_unsigned(29705, LUT_AMPL_WIDTH - 1),
		11840 => to_unsigned(29706, LUT_AMPL_WIDTH - 1),
		11841 => to_unsigned(29708, LUT_AMPL_WIDTH - 1),
		11842 => to_unsigned(29709, LUT_AMPL_WIDTH - 1),
		11843 => to_unsigned(29710, LUT_AMPL_WIDTH - 1),
		11844 => to_unsigned(29712, LUT_AMPL_WIDTH - 1),
		11845 => to_unsigned(29713, LUT_AMPL_WIDTH - 1),
		11846 => to_unsigned(29714, LUT_AMPL_WIDTH - 1),
		11847 => to_unsigned(29716, LUT_AMPL_WIDTH - 1),
		11848 => to_unsigned(29717, LUT_AMPL_WIDTH - 1),
		11849 => to_unsigned(29718, LUT_AMPL_WIDTH - 1),
		11850 => to_unsigned(29720, LUT_AMPL_WIDTH - 1),
		11851 => to_unsigned(29721, LUT_AMPL_WIDTH - 1),
		11852 => to_unsigned(29722, LUT_AMPL_WIDTH - 1),
		11853 => to_unsigned(29724, LUT_AMPL_WIDTH - 1),
		11854 => to_unsigned(29725, LUT_AMPL_WIDTH - 1),
		11855 => to_unsigned(29726, LUT_AMPL_WIDTH - 1),
		11856 => to_unsigned(29728, LUT_AMPL_WIDTH - 1),
		11857 => to_unsigned(29729, LUT_AMPL_WIDTH - 1),
		11858 => to_unsigned(29730, LUT_AMPL_WIDTH - 1),
		11859 => to_unsigned(29732, LUT_AMPL_WIDTH - 1),
		11860 => to_unsigned(29733, LUT_AMPL_WIDTH - 1),
		11861 => to_unsigned(29734, LUT_AMPL_WIDTH - 1),
		11862 => to_unsigned(29736, LUT_AMPL_WIDTH - 1),
		11863 => to_unsigned(29737, LUT_AMPL_WIDTH - 1),
		11864 => to_unsigned(29738, LUT_AMPL_WIDTH - 1),
		11865 => to_unsigned(29739, LUT_AMPL_WIDTH - 1),
		11866 => to_unsigned(29741, LUT_AMPL_WIDTH - 1),
		11867 => to_unsigned(29742, LUT_AMPL_WIDTH - 1),
		11868 => to_unsigned(29743, LUT_AMPL_WIDTH - 1),
		11869 => to_unsigned(29745, LUT_AMPL_WIDTH - 1),
		11870 => to_unsigned(29746, LUT_AMPL_WIDTH - 1),
		11871 => to_unsigned(29747, LUT_AMPL_WIDTH - 1),
		11872 => to_unsigned(29749, LUT_AMPL_WIDTH - 1),
		11873 => to_unsigned(29750, LUT_AMPL_WIDTH - 1),
		11874 => to_unsigned(29751, LUT_AMPL_WIDTH - 1),
		11875 => to_unsigned(29753, LUT_AMPL_WIDTH - 1),
		11876 => to_unsigned(29754, LUT_AMPL_WIDTH - 1),
		11877 => to_unsigned(29755, LUT_AMPL_WIDTH - 1),
		11878 => to_unsigned(29757, LUT_AMPL_WIDTH - 1),
		11879 => to_unsigned(29758, LUT_AMPL_WIDTH - 1),
		11880 => to_unsigned(29759, LUT_AMPL_WIDTH - 1),
		11881 => to_unsigned(29761, LUT_AMPL_WIDTH - 1),
		11882 => to_unsigned(29762, LUT_AMPL_WIDTH - 1),
		11883 => to_unsigned(29763, LUT_AMPL_WIDTH - 1),
		11884 => to_unsigned(29764, LUT_AMPL_WIDTH - 1),
		11885 => to_unsigned(29766, LUT_AMPL_WIDTH - 1),
		11886 => to_unsigned(29767, LUT_AMPL_WIDTH - 1),
		11887 => to_unsigned(29768, LUT_AMPL_WIDTH - 1),
		11888 => to_unsigned(29770, LUT_AMPL_WIDTH - 1),
		11889 => to_unsigned(29771, LUT_AMPL_WIDTH - 1),
		11890 => to_unsigned(29772, LUT_AMPL_WIDTH - 1),
		11891 => to_unsigned(29774, LUT_AMPL_WIDTH - 1),
		11892 => to_unsigned(29775, LUT_AMPL_WIDTH - 1),
		11893 => to_unsigned(29776, LUT_AMPL_WIDTH - 1),
		11894 => to_unsigned(29778, LUT_AMPL_WIDTH - 1),
		11895 => to_unsigned(29779, LUT_AMPL_WIDTH - 1),
		11896 => to_unsigned(29780, LUT_AMPL_WIDTH - 1),
		11897 => to_unsigned(29782, LUT_AMPL_WIDTH - 1),
		11898 => to_unsigned(29783, LUT_AMPL_WIDTH - 1),
		11899 => to_unsigned(29784, LUT_AMPL_WIDTH - 1),
		11900 => to_unsigned(29785, LUT_AMPL_WIDTH - 1),
		11901 => to_unsigned(29787, LUT_AMPL_WIDTH - 1),
		11902 => to_unsigned(29788, LUT_AMPL_WIDTH - 1),
		11903 => to_unsigned(29789, LUT_AMPL_WIDTH - 1),
		11904 => to_unsigned(29791, LUT_AMPL_WIDTH - 1),
		11905 => to_unsigned(29792, LUT_AMPL_WIDTH - 1),
		11906 => to_unsigned(29793, LUT_AMPL_WIDTH - 1),
		11907 => to_unsigned(29795, LUT_AMPL_WIDTH - 1),
		11908 => to_unsigned(29796, LUT_AMPL_WIDTH - 1),
		11909 => to_unsigned(29797, LUT_AMPL_WIDTH - 1),
		11910 => to_unsigned(29799, LUT_AMPL_WIDTH - 1),
		11911 => to_unsigned(29800, LUT_AMPL_WIDTH - 1),
		11912 => to_unsigned(29801, LUT_AMPL_WIDTH - 1),
		11913 => to_unsigned(29802, LUT_AMPL_WIDTH - 1),
		11914 => to_unsigned(29804, LUT_AMPL_WIDTH - 1),
		11915 => to_unsigned(29805, LUT_AMPL_WIDTH - 1),
		11916 => to_unsigned(29806, LUT_AMPL_WIDTH - 1),
		11917 => to_unsigned(29808, LUT_AMPL_WIDTH - 1),
		11918 => to_unsigned(29809, LUT_AMPL_WIDTH - 1),
		11919 => to_unsigned(29810, LUT_AMPL_WIDTH - 1),
		11920 => to_unsigned(29812, LUT_AMPL_WIDTH - 1),
		11921 => to_unsigned(29813, LUT_AMPL_WIDTH - 1),
		11922 => to_unsigned(29814, LUT_AMPL_WIDTH - 1),
		11923 => to_unsigned(29816, LUT_AMPL_WIDTH - 1),
		11924 => to_unsigned(29817, LUT_AMPL_WIDTH - 1),
		11925 => to_unsigned(29818, LUT_AMPL_WIDTH - 1),
		11926 => to_unsigned(29819, LUT_AMPL_WIDTH - 1),
		11927 => to_unsigned(29821, LUT_AMPL_WIDTH - 1),
		11928 => to_unsigned(29822, LUT_AMPL_WIDTH - 1),
		11929 => to_unsigned(29823, LUT_AMPL_WIDTH - 1),
		11930 => to_unsigned(29825, LUT_AMPL_WIDTH - 1),
		11931 => to_unsigned(29826, LUT_AMPL_WIDTH - 1),
		11932 => to_unsigned(29827, LUT_AMPL_WIDTH - 1),
		11933 => to_unsigned(29829, LUT_AMPL_WIDTH - 1),
		11934 => to_unsigned(29830, LUT_AMPL_WIDTH - 1),
		11935 => to_unsigned(29831, LUT_AMPL_WIDTH - 1),
		11936 => to_unsigned(29832, LUT_AMPL_WIDTH - 1),
		11937 => to_unsigned(29834, LUT_AMPL_WIDTH - 1),
		11938 => to_unsigned(29835, LUT_AMPL_WIDTH - 1),
		11939 => to_unsigned(29836, LUT_AMPL_WIDTH - 1),
		11940 => to_unsigned(29838, LUT_AMPL_WIDTH - 1),
		11941 => to_unsigned(29839, LUT_AMPL_WIDTH - 1),
		11942 => to_unsigned(29840, LUT_AMPL_WIDTH - 1),
		11943 => to_unsigned(29842, LUT_AMPL_WIDTH - 1),
		11944 => to_unsigned(29843, LUT_AMPL_WIDTH - 1),
		11945 => to_unsigned(29844, LUT_AMPL_WIDTH - 1),
		11946 => to_unsigned(29845, LUT_AMPL_WIDTH - 1),
		11947 => to_unsigned(29847, LUT_AMPL_WIDTH - 1),
		11948 => to_unsigned(29848, LUT_AMPL_WIDTH - 1),
		11949 => to_unsigned(29849, LUT_AMPL_WIDTH - 1),
		11950 => to_unsigned(29851, LUT_AMPL_WIDTH - 1),
		11951 => to_unsigned(29852, LUT_AMPL_WIDTH - 1),
		11952 => to_unsigned(29853, LUT_AMPL_WIDTH - 1),
		11953 => to_unsigned(29854, LUT_AMPL_WIDTH - 1),
		11954 => to_unsigned(29856, LUT_AMPL_WIDTH - 1),
		11955 => to_unsigned(29857, LUT_AMPL_WIDTH - 1),
		11956 => to_unsigned(29858, LUT_AMPL_WIDTH - 1),
		11957 => to_unsigned(29860, LUT_AMPL_WIDTH - 1),
		11958 => to_unsigned(29861, LUT_AMPL_WIDTH - 1),
		11959 => to_unsigned(29862, LUT_AMPL_WIDTH - 1),
		11960 => to_unsigned(29864, LUT_AMPL_WIDTH - 1),
		11961 => to_unsigned(29865, LUT_AMPL_WIDTH - 1),
		11962 => to_unsigned(29866, LUT_AMPL_WIDTH - 1),
		11963 => to_unsigned(29867, LUT_AMPL_WIDTH - 1),
		11964 => to_unsigned(29869, LUT_AMPL_WIDTH - 1),
		11965 => to_unsigned(29870, LUT_AMPL_WIDTH - 1),
		11966 => to_unsigned(29871, LUT_AMPL_WIDTH - 1),
		11967 => to_unsigned(29873, LUT_AMPL_WIDTH - 1),
		11968 => to_unsigned(29874, LUT_AMPL_WIDTH - 1),
		11969 => to_unsigned(29875, LUT_AMPL_WIDTH - 1),
		11970 => to_unsigned(29876, LUT_AMPL_WIDTH - 1),
		11971 => to_unsigned(29878, LUT_AMPL_WIDTH - 1),
		11972 => to_unsigned(29879, LUT_AMPL_WIDTH - 1),
		11973 => to_unsigned(29880, LUT_AMPL_WIDTH - 1),
		11974 => to_unsigned(29882, LUT_AMPL_WIDTH - 1),
		11975 => to_unsigned(29883, LUT_AMPL_WIDTH - 1),
		11976 => to_unsigned(29884, LUT_AMPL_WIDTH - 1),
		11977 => to_unsigned(29885, LUT_AMPL_WIDTH - 1),
		11978 => to_unsigned(29887, LUT_AMPL_WIDTH - 1),
		11979 => to_unsigned(29888, LUT_AMPL_WIDTH - 1),
		11980 => to_unsigned(29889, LUT_AMPL_WIDTH - 1),
		11981 => to_unsigned(29891, LUT_AMPL_WIDTH - 1),
		11982 => to_unsigned(29892, LUT_AMPL_WIDTH - 1),
		11983 => to_unsigned(29893, LUT_AMPL_WIDTH - 1),
		11984 => to_unsigned(29894, LUT_AMPL_WIDTH - 1),
		11985 => to_unsigned(29896, LUT_AMPL_WIDTH - 1),
		11986 => to_unsigned(29897, LUT_AMPL_WIDTH - 1),
		11987 => to_unsigned(29898, LUT_AMPL_WIDTH - 1),
		11988 => to_unsigned(29900, LUT_AMPL_WIDTH - 1),
		11989 => to_unsigned(29901, LUT_AMPL_WIDTH - 1),
		11990 => to_unsigned(29902, LUT_AMPL_WIDTH - 1),
		11991 => to_unsigned(29903, LUT_AMPL_WIDTH - 1),
		11992 => to_unsigned(29905, LUT_AMPL_WIDTH - 1),
		11993 => to_unsigned(29906, LUT_AMPL_WIDTH - 1),
		11994 => to_unsigned(29907, LUT_AMPL_WIDTH - 1),
		11995 => to_unsigned(29909, LUT_AMPL_WIDTH - 1),
		11996 => to_unsigned(29910, LUT_AMPL_WIDTH - 1),
		11997 => to_unsigned(29911, LUT_AMPL_WIDTH - 1),
		11998 => to_unsigned(29912, LUT_AMPL_WIDTH - 1),
		11999 => to_unsigned(29914, LUT_AMPL_WIDTH - 1),
		12000 => to_unsigned(29915, LUT_AMPL_WIDTH - 1),
		12001 => to_unsigned(29916, LUT_AMPL_WIDTH - 1),
		12002 => to_unsigned(29918, LUT_AMPL_WIDTH - 1),
		12003 => to_unsigned(29919, LUT_AMPL_WIDTH - 1),
		12004 => to_unsigned(29920, LUT_AMPL_WIDTH - 1),
		12005 => to_unsigned(29921, LUT_AMPL_WIDTH - 1),
		12006 => to_unsigned(29923, LUT_AMPL_WIDTH - 1),
		12007 => to_unsigned(29924, LUT_AMPL_WIDTH - 1),
		12008 => to_unsigned(29925, LUT_AMPL_WIDTH - 1),
		12009 => to_unsigned(29927, LUT_AMPL_WIDTH - 1),
		12010 => to_unsigned(29928, LUT_AMPL_WIDTH - 1),
		12011 => to_unsigned(29929, LUT_AMPL_WIDTH - 1),
		12012 => to_unsigned(29930, LUT_AMPL_WIDTH - 1),
		12013 => to_unsigned(29932, LUT_AMPL_WIDTH - 1),
		12014 => to_unsigned(29933, LUT_AMPL_WIDTH - 1),
		12015 => to_unsigned(29934, LUT_AMPL_WIDTH - 1),
		12016 => to_unsigned(29936, LUT_AMPL_WIDTH - 1),
		12017 => to_unsigned(29937, LUT_AMPL_WIDTH - 1),
		12018 => to_unsigned(29938, LUT_AMPL_WIDTH - 1),
		12019 => to_unsigned(29939, LUT_AMPL_WIDTH - 1),
		12020 => to_unsigned(29941, LUT_AMPL_WIDTH - 1),
		12021 => to_unsigned(29942, LUT_AMPL_WIDTH - 1),
		12022 => to_unsigned(29943, LUT_AMPL_WIDTH - 1),
		12023 => to_unsigned(29944, LUT_AMPL_WIDTH - 1),
		12024 => to_unsigned(29946, LUT_AMPL_WIDTH - 1),
		12025 => to_unsigned(29947, LUT_AMPL_WIDTH - 1),
		12026 => to_unsigned(29948, LUT_AMPL_WIDTH - 1),
		12027 => to_unsigned(29950, LUT_AMPL_WIDTH - 1),
		12028 => to_unsigned(29951, LUT_AMPL_WIDTH - 1),
		12029 => to_unsigned(29952, LUT_AMPL_WIDTH - 1),
		12030 => to_unsigned(29953, LUT_AMPL_WIDTH - 1),
		12031 => to_unsigned(29955, LUT_AMPL_WIDTH - 1),
		12032 => to_unsigned(29956, LUT_AMPL_WIDTH - 1),
		12033 => to_unsigned(29957, LUT_AMPL_WIDTH - 1),
		12034 => to_unsigned(29958, LUT_AMPL_WIDTH - 1),
		12035 => to_unsigned(29960, LUT_AMPL_WIDTH - 1),
		12036 => to_unsigned(29961, LUT_AMPL_WIDTH - 1),
		12037 => to_unsigned(29962, LUT_AMPL_WIDTH - 1),
		12038 => to_unsigned(29964, LUT_AMPL_WIDTH - 1),
		12039 => to_unsigned(29965, LUT_AMPL_WIDTH - 1),
		12040 => to_unsigned(29966, LUT_AMPL_WIDTH - 1),
		12041 => to_unsigned(29967, LUT_AMPL_WIDTH - 1),
		12042 => to_unsigned(29969, LUT_AMPL_WIDTH - 1),
		12043 => to_unsigned(29970, LUT_AMPL_WIDTH - 1),
		12044 => to_unsigned(29971, LUT_AMPL_WIDTH - 1),
		12045 => to_unsigned(29972, LUT_AMPL_WIDTH - 1),
		12046 => to_unsigned(29974, LUT_AMPL_WIDTH - 1),
		12047 => to_unsigned(29975, LUT_AMPL_WIDTH - 1),
		12048 => to_unsigned(29976, LUT_AMPL_WIDTH - 1),
		12049 => to_unsigned(29978, LUT_AMPL_WIDTH - 1),
		12050 => to_unsigned(29979, LUT_AMPL_WIDTH - 1),
		12051 => to_unsigned(29980, LUT_AMPL_WIDTH - 1),
		12052 => to_unsigned(29981, LUT_AMPL_WIDTH - 1),
		12053 => to_unsigned(29983, LUT_AMPL_WIDTH - 1),
		12054 => to_unsigned(29984, LUT_AMPL_WIDTH - 1),
		12055 => to_unsigned(29985, LUT_AMPL_WIDTH - 1),
		12056 => to_unsigned(29986, LUT_AMPL_WIDTH - 1),
		12057 => to_unsigned(29988, LUT_AMPL_WIDTH - 1),
		12058 => to_unsigned(29989, LUT_AMPL_WIDTH - 1),
		12059 => to_unsigned(29990, LUT_AMPL_WIDTH - 1),
		12060 => to_unsigned(29991, LUT_AMPL_WIDTH - 1),
		12061 => to_unsigned(29993, LUT_AMPL_WIDTH - 1),
		12062 => to_unsigned(29994, LUT_AMPL_WIDTH - 1),
		12063 => to_unsigned(29995, LUT_AMPL_WIDTH - 1),
		12064 => to_unsigned(29997, LUT_AMPL_WIDTH - 1),
		12065 => to_unsigned(29998, LUT_AMPL_WIDTH - 1),
		12066 => to_unsigned(29999, LUT_AMPL_WIDTH - 1),
		12067 => to_unsigned(30000, LUT_AMPL_WIDTH - 1),
		12068 => to_unsigned(30002, LUT_AMPL_WIDTH - 1),
		12069 => to_unsigned(30003, LUT_AMPL_WIDTH - 1),
		12070 => to_unsigned(30004, LUT_AMPL_WIDTH - 1),
		12071 => to_unsigned(30005, LUT_AMPL_WIDTH - 1),
		12072 => to_unsigned(30007, LUT_AMPL_WIDTH - 1),
		12073 => to_unsigned(30008, LUT_AMPL_WIDTH - 1),
		12074 => to_unsigned(30009, LUT_AMPL_WIDTH - 1),
		12075 => to_unsigned(30010, LUT_AMPL_WIDTH - 1),
		12076 => to_unsigned(30012, LUT_AMPL_WIDTH - 1),
		12077 => to_unsigned(30013, LUT_AMPL_WIDTH - 1),
		12078 => to_unsigned(30014, LUT_AMPL_WIDTH - 1),
		12079 => to_unsigned(30015, LUT_AMPL_WIDTH - 1),
		12080 => to_unsigned(30017, LUT_AMPL_WIDTH - 1),
		12081 => to_unsigned(30018, LUT_AMPL_WIDTH - 1),
		12082 => to_unsigned(30019, LUT_AMPL_WIDTH - 1),
		12083 => to_unsigned(30020, LUT_AMPL_WIDTH - 1),
		12084 => to_unsigned(30022, LUT_AMPL_WIDTH - 1),
		12085 => to_unsigned(30023, LUT_AMPL_WIDTH - 1),
		12086 => to_unsigned(30024, LUT_AMPL_WIDTH - 1),
		12087 => to_unsigned(30026, LUT_AMPL_WIDTH - 1),
		12088 => to_unsigned(30027, LUT_AMPL_WIDTH - 1),
		12089 => to_unsigned(30028, LUT_AMPL_WIDTH - 1),
		12090 => to_unsigned(30029, LUT_AMPL_WIDTH - 1),
		12091 => to_unsigned(30031, LUT_AMPL_WIDTH - 1),
		12092 => to_unsigned(30032, LUT_AMPL_WIDTH - 1),
		12093 => to_unsigned(30033, LUT_AMPL_WIDTH - 1),
		12094 => to_unsigned(30034, LUT_AMPL_WIDTH - 1),
		12095 => to_unsigned(30036, LUT_AMPL_WIDTH - 1),
		12096 => to_unsigned(30037, LUT_AMPL_WIDTH - 1),
		12097 => to_unsigned(30038, LUT_AMPL_WIDTH - 1),
		12098 => to_unsigned(30039, LUT_AMPL_WIDTH - 1),
		12099 => to_unsigned(30041, LUT_AMPL_WIDTH - 1),
		12100 => to_unsigned(30042, LUT_AMPL_WIDTH - 1),
		12101 => to_unsigned(30043, LUT_AMPL_WIDTH - 1),
		12102 => to_unsigned(30044, LUT_AMPL_WIDTH - 1),
		12103 => to_unsigned(30046, LUT_AMPL_WIDTH - 1),
		12104 => to_unsigned(30047, LUT_AMPL_WIDTH - 1),
		12105 => to_unsigned(30048, LUT_AMPL_WIDTH - 1),
		12106 => to_unsigned(30049, LUT_AMPL_WIDTH - 1),
		12107 => to_unsigned(30051, LUT_AMPL_WIDTH - 1),
		12108 => to_unsigned(30052, LUT_AMPL_WIDTH - 1),
		12109 => to_unsigned(30053, LUT_AMPL_WIDTH - 1),
		12110 => to_unsigned(30054, LUT_AMPL_WIDTH - 1),
		12111 => to_unsigned(30056, LUT_AMPL_WIDTH - 1),
		12112 => to_unsigned(30057, LUT_AMPL_WIDTH - 1),
		12113 => to_unsigned(30058, LUT_AMPL_WIDTH - 1),
		12114 => to_unsigned(30059, LUT_AMPL_WIDTH - 1),
		12115 => to_unsigned(30061, LUT_AMPL_WIDTH - 1),
		12116 => to_unsigned(30062, LUT_AMPL_WIDTH - 1),
		12117 => to_unsigned(30063, LUT_AMPL_WIDTH - 1),
		12118 => to_unsigned(30064, LUT_AMPL_WIDTH - 1),
		12119 => to_unsigned(30066, LUT_AMPL_WIDTH - 1),
		12120 => to_unsigned(30067, LUT_AMPL_WIDTH - 1),
		12121 => to_unsigned(30068, LUT_AMPL_WIDTH - 1),
		12122 => to_unsigned(30069, LUT_AMPL_WIDTH - 1),
		12123 => to_unsigned(30071, LUT_AMPL_WIDTH - 1),
		12124 => to_unsigned(30072, LUT_AMPL_WIDTH - 1),
		12125 => to_unsigned(30073, LUT_AMPL_WIDTH - 1),
		12126 => to_unsigned(30074, LUT_AMPL_WIDTH - 1),
		12127 => to_unsigned(30076, LUT_AMPL_WIDTH - 1),
		12128 => to_unsigned(30077, LUT_AMPL_WIDTH - 1),
		12129 => to_unsigned(30078, LUT_AMPL_WIDTH - 1),
		12130 => to_unsigned(30079, LUT_AMPL_WIDTH - 1),
		12131 => to_unsigned(30081, LUT_AMPL_WIDTH - 1),
		12132 => to_unsigned(30082, LUT_AMPL_WIDTH - 1),
		12133 => to_unsigned(30083, LUT_AMPL_WIDTH - 1),
		12134 => to_unsigned(30084, LUT_AMPL_WIDTH - 1),
		12135 => to_unsigned(30086, LUT_AMPL_WIDTH - 1),
		12136 => to_unsigned(30087, LUT_AMPL_WIDTH - 1),
		12137 => to_unsigned(30088, LUT_AMPL_WIDTH - 1),
		12138 => to_unsigned(30089, LUT_AMPL_WIDTH - 1),
		12139 => to_unsigned(30091, LUT_AMPL_WIDTH - 1),
		12140 => to_unsigned(30092, LUT_AMPL_WIDTH - 1),
		12141 => to_unsigned(30093, LUT_AMPL_WIDTH - 1),
		12142 => to_unsigned(30094, LUT_AMPL_WIDTH - 1),
		12143 => to_unsigned(30096, LUT_AMPL_WIDTH - 1),
		12144 => to_unsigned(30097, LUT_AMPL_WIDTH - 1),
		12145 => to_unsigned(30098, LUT_AMPL_WIDTH - 1),
		12146 => to_unsigned(30099, LUT_AMPL_WIDTH - 1),
		12147 => to_unsigned(30100, LUT_AMPL_WIDTH - 1),
		12148 => to_unsigned(30102, LUT_AMPL_WIDTH - 1),
		12149 => to_unsigned(30103, LUT_AMPL_WIDTH - 1),
		12150 => to_unsigned(30104, LUT_AMPL_WIDTH - 1),
		12151 => to_unsigned(30105, LUT_AMPL_WIDTH - 1),
		12152 => to_unsigned(30107, LUT_AMPL_WIDTH - 1),
		12153 => to_unsigned(30108, LUT_AMPL_WIDTH - 1),
		12154 => to_unsigned(30109, LUT_AMPL_WIDTH - 1),
		12155 => to_unsigned(30110, LUT_AMPL_WIDTH - 1),
		12156 => to_unsigned(30112, LUT_AMPL_WIDTH - 1),
		12157 => to_unsigned(30113, LUT_AMPL_WIDTH - 1),
		12158 => to_unsigned(30114, LUT_AMPL_WIDTH - 1),
		12159 => to_unsigned(30115, LUT_AMPL_WIDTH - 1),
		12160 => to_unsigned(30117, LUT_AMPL_WIDTH - 1),
		12161 => to_unsigned(30118, LUT_AMPL_WIDTH - 1),
		12162 => to_unsigned(30119, LUT_AMPL_WIDTH - 1),
		12163 => to_unsigned(30120, LUT_AMPL_WIDTH - 1),
		12164 => to_unsigned(30122, LUT_AMPL_WIDTH - 1),
		12165 => to_unsigned(30123, LUT_AMPL_WIDTH - 1),
		12166 => to_unsigned(30124, LUT_AMPL_WIDTH - 1),
		12167 => to_unsigned(30125, LUT_AMPL_WIDTH - 1),
		12168 => to_unsigned(30126, LUT_AMPL_WIDTH - 1),
		12169 => to_unsigned(30128, LUT_AMPL_WIDTH - 1),
		12170 => to_unsigned(30129, LUT_AMPL_WIDTH - 1),
		12171 => to_unsigned(30130, LUT_AMPL_WIDTH - 1),
		12172 => to_unsigned(30131, LUT_AMPL_WIDTH - 1),
		12173 => to_unsigned(30133, LUT_AMPL_WIDTH - 1),
		12174 => to_unsigned(30134, LUT_AMPL_WIDTH - 1),
		12175 => to_unsigned(30135, LUT_AMPL_WIDTH - 1),
		12176 => to_unsigned(30136, LUT_AMPL_WIDTH - 1),
		12177 => to_unsigned(30138, LUT_AMPL_WIDTH - 1),
		12178 => to_unsigned(30139, LUT_AMPL_WIDTH - 1),
		12179 => to_unsigned(30140, LUT_AMPL_WIDTH - 1),
		12180 => to_unsigned(30141, LUT_AMPL_WIDTH - 1),
		12181 => to_unsigned(30143, LUT_AMPL_WIDTH - 1),
		12182 => to_unsigned(30144, LUT_AMPL_WIDTH - 1),
		12183 => to_unsigned(30145, LUT_AMPL_WIDTH - 1),
		12184 => to_unsigned(30146, LUT_AMPL_WIDTH - 1),
		12185 => to_unsigned(30147, LUT_AMPL_WIDTH - 1),
		12186 => to_unsigned(30149, LUT_AMPL_WIDTH - 1),
		12187 => to_unsigned(30150, LUT_AMPL_WIDTH - 1),
		12188 => to_unsigned(30151, LUT_AMPL_WIDTH - 1),
		12189 => to_unsigned(30152, LUT_AMPL_WIDTH - 1),
		12190 => to_unsigned(30154, LUT_AMPL_WIDTH - 1),
		12191 => to_unsigned(30155, LUT_AMPL_WIDTH - 1),
		12192 => to_unsigned(30156, LUT_AMPL_WIDTH - 1),
		12193 => to_unsigned(30157, LUT_AMPL_WIDTH - 1),
		12194 => to_unsigned(30159, LUT_AMPL_WIDTH - 1),
		12195 => to_unsigned(30160, LUT_AMPL_WIDTH - 1),
		12196 => to_unsigned(30161, LUT_AMPL_WIDTH - 1),
		12197 => to_unsigned(30162, LUT_AMPL_WIDTH - 1),
		12198 => to_unsigned(30163, LUT_AMPL_WIDTH - 1),
		12199 => to_unsigned(30165, LUT_AMPL_WIDTH - 1),
		12200 => to_unsigned(30166, LUT_AMPL_WIDTH - 1),
		12201 => to_unsigned(30167, LUT_AMPL_WIDTH - 1),
		12202 => to_unsigned(30168, LUT_AMPL_WIDTH - 1),
		12203 => to_unsigned(30170, LUT_AMPL_WIDTH - 1),
		12204 => to_unsigned(30171, LUT_AMPL_WIDTH - 1),
		12205 => to_unsigned(30172, LUT_AMPL_WIDTH - 1),
		12206 => to_unsigned(30173, LUT_AMPL_WIDTH - 1),
		12207 => to_unsigned(30174, LUT_AMPL_WIDTH - 1),
		12208 => to_unsigned(30176, LUT_AMPL_WIDTH - 1),
		12209 => to_unsigned(30177, LUT_AMPL_WIDTH - 1),
		12210 => to_unsigned(30178, LUT_AMPL_WIDTH - 1),
		12211 => to_unsigned(30179, LUT_AMPL_WIDTH - 1),
		12212 => to_unsigned(30181, LUT_AMPL_WIDTH - 1),
		12213 => to_unsigned(30182, LUT_AMPL_WIDTH - 1),
		12214 => to_unsigned(30183, LUT_AMPL_WIDTH - 1),
		12215 => to_unsigned(30184, LUT_AMPL_WIDTH - 1),
		12216 => to_unsigned(30185, LUT_AMPL_WIDTH - 1),
		12217 => to_unsigned(30187, LUT_AMPL_WIDTH - 1),
		12218 => to_unsigned(30188, LUT_AMPL_WIDTH - 1),
		12219 => to_unsigned(30189, LUT_AMPL_WIDTH - 1),
		12220 => to_unsigned(30190, LUT_AMPL_WIDTH - 1),
		12221 => to_unsigned(30192, LUT_AMPL_WIDTH - 1),
		12222 => to_unsigned(30193, LUT_AMPL_WIDTH - 1),
		12223 => to_unsigned(30194, LUT_AMPL_WIDTH - 1),
		12224 => to_unsigned(30195, LUT_AMPL_WIDTH - 1),
		12225 => to_unsigned(30196, LUT_AMPL_WIDTH - 1),
		12226 => to_unsigned(30198, LUT_AMPL_WIDTH - 1),
		12227 => to_unsigned(30199, LUT_AMPL_WIDTH - 1),
		12228 => to_unsigned(30200, LUT_AMPL_WIDTH - 1),
		12229 => to_unsigned(30201, LUT_AMPL_WIDTH - 1),
		12230 => to_unsigned(30203, LUT_AMPL_WIDTH - 1),
		12231 => to_unsigned(30204, LUT_AMPL_WIDTH - 1),
		12232 => to_unsigned(30205, LUT_AMPL_WIDTH - 1),
		12233 => to_unsigned(30206, LUT_AMPL_WIDTH - 1),
		12234 => to_unsigned(30207, LUT_AMPL_WIDTH - 1),
		12235 => to_unsigned(30209, LUT_AMPL_WIDTH - 1),
		12236 => to_unsigned(30210, LUT_AMPL_WIDTH - 1),
		12237 => to_unsigned(30211, LUT_AMPL_WIDTH - 1),
		12238 => to_unsigned(30212, LUT_AMPL_WIDTH - 1),
		12239 => to_unsigned(30214, LUT_AMPL_WIDTH - 1),
		12240 => to_unsigned(30215, LUT_AMPL_WIDTH - 1),
		12241 => to_unsigned(30216, LUT_AMPL_WIDTH - 1),
		12242 => to_unsigned(30217, LUT_AMPL_WIDTH - 1),
		12243 => to_unsigned(30218, LUT_AMPL_WIDTH - 1),
		12244 => to_unsigned(30220, LUT_AMPL_WIDTH - 1),
		12245 => to_unsigned(30221, LUT_AMPL_WIDTH - 1),
		12246 => to_unsigned(30222, LUT_AMPL_WIDTH - 1),
		12247 => to_unsigned(30223, LUT_AMPL_WIDTH - 1),
		12248 => to_unsigned(30224, LUT_AMPL_WIDTH - 1),
		12249 => to_unsigned(30226, LUT_AMPL_WIDTH - 1),
		12250 => to_unsigned(30227, LUT_AMPL_WIDTH - 1),
		12251 => to_unsigned(30228, LUT_AMPL_WIDTH - 1),
		12252 => to_unsigned(30229, LUT_AMPL_WIDTH - 1),
		12253 => to_unsigned(30231, LUT_AMPL_WIDTH - 1),
		12254 => to_unsigned(30232, LUT_AMPL_WIDTH - 1),
		12255 => to_unsigned(30233, LUT_AMPL_WIDTH - 1),
		12256 => to_unsigned(30234, LUT_AMPL_WIDTH - 1),
		12257 => to_unsigned(30235, LUT_AMPL_WIDTH - 1),
		12258 => to_unsigned(30237, LUT_AMPL_WIDTH - 1),
		12259 => to_unsigned(30238, LUT_AMPL_WIDTH - 1),
		12260 => to_unsigned(30239, LUT_AMPL_WIDTH - 1),
		12261 => to_unsigned(30240, LUT_AMPL_WIDTH - 1),
		12262 => to_unsigned(30241, LUT_AMPL_WIDTH - 1),
		12263 => to_unsigned(30243, LUT_AMPL_WIDTH - 1),
		12264 => to_unsigned(30244, LUT_AMPL_WIDTH - 1),
		12265 => to_unsigned(30245, LUT_AMPL_WIDTH - 1),
		12266 => to_unsigned(30246, LUT_AMPL_WIDTH - 1),
		12267 => to_unsigned(30247, LUT_AMPL_WIDTH - 1),
		12268 => to_unsigned(30249, LUT_AMPL_WIDTH - 1),
		12269 => to_unsigned(30250, LUT_AMPL_WIDTH - 1),
		12270 => to_unsigned(30251, LUT_AMPL_WIDTH - 1),
		12271 => to_unsigned(30252, LUT_AMPL_WIDTH - 1),
		12272 => to_unsigned(30253, LUT_AMPL_WIDTH - 1),
		12273 => to_unsigned(30255, LUT_AMPL_WIDTH - 1),
		12274 => to_unsigned(30256, LUT_AMPL_WIDTH - 1),
		12275 => to_unsigned(30257, LUT_AMPL_WIDTH - 1),
		12276 => to_unsigned(30258, LUT_AMPL_WIDTH - 1),
		12277 => to_unsigned(30260, LUT_AMPL_WIDTH - 1),
		12278 => to_unsigned(30261, LUT_AMPL_WIDTH - 1),
		12279 => to_unsigned(30262, LUT_AMPL_WIDTH - 1),
		12280 => to_unsigned(30263, LUT_AMPL_WIDTH - 1),
		12281 => to_unsigned(30264, LUT_AMPL_WIDTH - 1),
		12282 => to_unsigned(30266, LUT_AMPL_WIDTH - 1),
		12283 => to_unsigned(30267, LUT_AMPL_WIDTH - 1),
		12284 => to_unsigned(30268, LUT_AMPL_WIDTH - 1),
		12285 => to_unsigned(30269, LUT_AMPL_WIDTH - 1),
		12286 => to_unsigned(30270, LUT_AMPL_WIDTH - 1),
		12287 => to_unsigned(30272, LUT_AMPL_WIDTH - 1),
		12288 => to_unsigned(30273, LUT_AMPL_WIDTH - 1),
		12289 => to_unsigned(30274, LUT_AMPL_WIDTH - 1),
		12290 => to_unsigned(30275, LUT_AMPL_WIDTH - 1),
		12291 => to_unsigned(30276, LUT_AMPL_WIDTH - 1),
		12292 => to_unsigned(30278, LUT_AMPL_WIDTH - 1),
		12293 => to_unsigned(30279, LUT_AMPL_WIDTH - 1),
		12294 => to_unsigned(30280, LUT_AMPL_WIDTH - 1),
		12295 => to_unsigned(30281, LUT_AMPL_WIDTH - 1),
		12296 => to_unsigned(30282, LUT_AMPL_WIDTH - 1),
		12297 => to_unsigned(30284, LUT_AMPL_WIDTH - 1),
		12298 => to_unsigned(30285, LUT_AMPL_WIDTH - 1),
		12299 => to_unsigned(30286, LUT_AMPL_WIDTH - 1),
		12300 => to_unsigned(30287, LUT_AMPL_WIDTH - 1),
		12301 => to_unsigned(30288, LUT_AMPL_WIDTH - 1),
		12302 => to_unsigned(30290, LUT_AMPL_WIDTH - 1),
		12303 => to_unsigned(30291, LUT_AMPL_WIDTH - 1),
		12304 => to_unsigned(30292, LUT_AMPL_WIDTH - 1),
		12305 => to_unsigned(30293, LUT_AMPL_WIDTH - 1),
		12306 => to_unsigned(30294, LUT_AMPL_WIDTH - 1),
		12307 => to_unsigned(30296, LUT_AMPL_WIDTH - 1),
		12308 => to_unsigned(30297, LUT_AMPL_WIDTH - 1),
		12309 => to_unsigned(30298, LUT_AMPL_WIDTH - 1),
		12310 => to_unsigned(30299, LUT_AMPL_WIDTH - 1),
		12311 => to_unsigned(30300, LUT_AMPL_WIDTH - 1),
		12312 => to_unsigned(30302, LUT_AMPL_WIDTH - 1),
		12313 => to_unsigned(30303, LUT_AMPL_WIDTH - 1),
		12314 => to_unsigned(30304, LUT_AMPL_WIDTH - 1),
		12315 => to_unsigned(30305, LUT_AMPL_WIDTH - 1),
		12316 => to_unsigned(30306, LUT_AMPL_WIDTH - 1),
		12317 => to_unsigned(30308, LUT_AMPL_WIDTH - 1),
		12318 => to_unsigned(30309, LUT_AMPL_WIDTH - 1),
		12319 => to_unsigned(30310, LUT_AMPL_WIDTH - 1),
		12320 => to_unsigned(30311, LUT_AMPL_WIDTH - 1),
		12321 => to_unsigned(30312, LUT_AMPL_WIDTH - 1),
		12322 => to_unsigned(30313, LUT_AMPL_WIDTH - 1),
		12323 => to_unsigned(30315, LUT_AMPL_WIDTH - 1),
		12324 => to_unsigned(30316, LUT_AMPL_WIDTH - 1),
		12325 => to_unsigned(30317, LUT_AMPL_WIDTH - 1),
		12326 => to_unsigned(30318, LUT_AMPL_WIDTH - 1),
		12327 => to_unsigned(30319, LUT_AMPL_WIDTH - 1),
		12328 => to_unsigned(30321, LUT_AMPL_WIDTH - 1),
		12329 => to_unsigned(30322, LUT_AMPL_WIDTH - 1),
		12330 => to_unsigned(30323, LUT_AMPL_WIDTH - 1),
		12331 => to_unsigned(30324, LUT_AMPL_WIDTH - 1),
		12332 => to_unsigned(30325, LUT_AMPL_WIDTH - 1),
		12333 => to_unsigned(30327, LUT_AMPL_WIDTH - 1),
		12334 => to_unsigned(30328, LUT_AMPL_WIDTH - 1),
		12335 => to_unsigned(30329, LUT_AMPL_WIDTH - 1),
		12336 => to_unsigned(30330, LUT_AMPL_WIDTH - 1),
		12337 => to_unsigned(30331, LUT_AMPL_WIDTH - 1),
		12338 => to_unsigned(30333, LUT_AMPL_WIDTH - 1),
		12339 => to_unsigned(30334, LUT_AMPL_WIDTH - 1),
		12340 => to_unsigned(30335, LUT_AMPL_WIDTH - 1),
		12341 => to_unsigned(30336, LUT_AMPL_WIDTH - 1),
		12342 => to_unsigned(30337, LUT_AMPL_WIDTH - 1),
		12343 => to_unsigned(30338, LUT_AMPL_WIDTH - 1),
		12344 => to_unsigned(30340, LUT_AMPL_WIDTH - 1),
		12345 => to_unsigned(30341, LUT_AMPL_WIDTH - 1),
		12346 => to_unsigned(30342, LUT_AMPL_WIDTH - 1),
		12347 => to_unsigned(30343, LUT_AMPL_WIDTH - 1),
		12348 => to_unsigned(30344, LUT_AMPL_WIDTH - 1),
		12349 => to_unsigned(30346, LUT_AMPL_WIDTH - 1),
		12350 => to_unsigned(30347, LUT_AMPL_WIDTH - 1),
		12351 => to_unsigned(30348, LUT_AMPL_WIDTH - 1),
		12352 => to_unsigned(30349, LUT_AMPL_WIDTH - 1),
		12353 => to_unsigned(30350, LUT_AMPL_WIDTH - 1),
		12354 => to_unsigned(30351, LUT_AMPL_WIDTH - 1),
		12355 => to_unsigned(30353, LUT_AMPL_WIDTH - 1),
		12356 => to_unsigned(30354, LUT_AMPL_WIDTH - 1),
		12357 => to_unsigned(30355, LUT_AMPL_WIDTH - 1),
		12358 => to_unsigned(30356, LUT_AMPL_WIDTH - 1),
		12359 => to_unsigned(30357, LUT_AMPL_WIDTH - 1),
		12360 => to_unsigned(30359, LUT_AMPL_WIDTH - 1),
		12361 => to_unsigned(30360, LUT_AMPL_WIDTH - 1),
		12362 => to_unsigned(30361, LUT_AMPL_WIDTH - 1),
		12363 => to_unsigned(30362, LUT_AMPL_WIDTH - 1),
		12364 => to_unsigned(30363, LUT_AMPL_WIDTH - 1),
		12365 => to_unsigned(30365, LUT_AMPL_WIDTH - 1),
		12366 => to_unsigned(30366, LUT_AMPL_WIDTH - 1),
		12367 => to_unsigned(30367, LUT_AMPL_WIDTH - 1),
		12368 => to_unsigned(30368, LUT_AMPL_WIDTH - 1),
		12369 => to_unsigned(30369, LUT_AMPL_WIDTH - 1),
		12370 => to_unsigned(30370, LUT_AMPL_WIDTH - 1),
		12371 => to_unsigned(30372, LUT_AMPL_WIDTH - 1),
		12372 => to_unsigned(30373, LUT_AMPL_WIDTH - 1),
		12373 => to_unsigned(30374, LUT_AMPL_WIDTH - 1),
		12374 => to_unsigned(30375, LUT_AMPL_WIDTH - 1),
		12375 => to_unsigned(30376, LUT_AMPL_WIDTH - 1),
		12376 => to_unsigned(30377, LUT_AMPL_WIDTH - 1),
		12377 => to_unsigned(30379, LUT_AMPL_WIDTH - 1),
		12378 => to_unsigned(30380, LUT_AMPL_WIDTH - 1),
		12379 => to_unsigned(30381, LUT_AMPL_WIDTH - 1),
		12380 => to_unsigned(30382, LUT_AMPL_WIDTH - 1),
		12381 => to_unsigned(30383, LUT_AMPL_WIDTH - 1),
		12382 => to_unsigned(30385, LUT_AMPL_WIDTH - 1),
		12383 => to_unsigned(30386, LUT_AMPL_WIDTH - 1),
		12384 => to_unsigned(30387, LUT_AMPL_WIDTH - 1),
		12385 => to_unsigned(30388, LUT_AMPL_WIDTH - 1),
		12386 => to_unsigned(30389, LUT_AMPL_WIDTH - 1),
		12387 => to_unsigned(30390, LUT_AMPL_WIDTH - 1),
		12388 => to_unsigned(30392, LUT_AMPL_WIDTH - 1),
		12389 => to_unsigned(30393, LUT_AMPL_WIDTH - 1),
		12390 => to_unsigned(30394, LUT_AMPL_WIDTH - 1),
		12391 => to_unsigned(30395, LUT_AMPL_WIDTH - 1),
		12392 => to_unsigned(30396, LUT_AMPL_WIDTH - 1),
		12393 => to_unsigned(30397, LUT_AMPL_WIDTH - 1),
		12394 => to_unsigned(30399, LUT_AMPL_WIDTH - 1),
		12395 => to_unsigned(30400, LUT_AMPL_WIDTH - 1),
		12396 => to_unsigned(30401, LUT_AMPL_WIDTH - 1),
		12397 => to_unsigned(30402, LUT_AMPL_WIDTH - 1),
		12398 => to_unsigned(30403, LUT_AMPL_WIDTH - 1),
		12399 => to_unsigned(30404, LUT_AMPL_WIDTH - 1),
		12400 => to_unsigned(30406, LUT_AMPL_WIDTH - 1),
		12401 => to_unsigned(30407, LUT_AMPL_WIDTH - 1),
		12402 => to_unsigned(30408, LUT_AMPL_WIDTH - 1),
		12403 => to_unsigned(30409, LUT_AMPL_WIDTH - 1),
		12404 => to_unsigned(30410, LUT_AMPL_WIDTH - 1),
		12405 => to_unsigned(30412, LUT_AMPL_WIDTH - 1),
		12406 => to_unsigned(30413, LUT_AMPL_WIDTH - 1),
		12407 => to_unsigned(30414, LUT_AMPL_WIDTH - 1),
		12408 => to_unsigned(30415, LUT_AMPL_WIDTH - 1),
		12409 => to_unsigned(30416, LUT_AMPL_WIDTH - 1),
		12410 => to_unsigned(30417, LUT_AMPL_WIDTH - 1),
		12411 => to_unsigned(30419, LUT_AMPL_WIDTH - 1),
		12412 => to_unsigned(30420, LUT_AMPL_WIDTH - 1),
		12413 => to_unsigned(30421, LUT_AMPL_WIDTH - 1),
		12414 => to_unsigned(30422, LUT_AMPL_WIDTH - 1),
		12415 => to_unsigned(30423, LUT_AMPL_WIDTH - 1),
		12416 => to_unsigned(30424, LUT_AMPL_WIDTH - 1),
		12417 => to_unsigned(30426, LUT_AMPL_WIDTH - 1),
		12418 => to_unsigned(30427, LUT_AMPL_WIDTH - 1),
		12419 => to_unsigned(30428, LUT_AMPL_WIDTH - 1),
		12420 => to_unsigned(30429, LUT_AMPL_WIDTH - 1),
		12421 => to_unsigned(30430, LUT_AMPL_WIDTH - 1),
		12422 => to_unsigned(30431, LUT_AMPL_WIDTH - 1),
		12423 => to_unsigned(30433, LUT_AMPL_WIDTH - 1),
		12424 => to_unsigned(30434, LUT_AMPL_WIDTH - 1),
		12425 => to_unsigned(30435, LUT_AMPL_WIDTH - 1),
		12426 => to_unsigned(30436, LUT_AMPL_WIDTH - 1),
		12427 => to_unsigned(30437, LUT_AMPL_WIDTH - 1),
		12428 => to_unsigned(30438, LUT_AMPL_WIDTH - 1),
		12429 => to_unsigned(30439, LUT_AMPL_WIDTH - 1),
		12430 => to_unsigned(30441, LUT_AMPL_WIDTH - 1),
		12431 => to_unsigned(30442, LUT_AMPL_WIDTH - 1),
		12432 => to_unsigned(30443, LUT_AMPL_WIDTH - 1),
		12433 => to_unsigned(30444, LUT_AMPL_WIDTH - 1),
		12434 => to_unsigned(30445, LUT_AMPL_WIDTH - 1),
		12435 => to_unsigned(30446, LUT_AMPL_WIDTH - 1),
		12436 => to_unsigned(30448, LUT_AMPL_WIDTH - 1),
		12437 => to_unsigned(30449, LUT_AMPL_WIDTH - 1),
		12438 => to_unsigned(30450, LUT_AMPL_WIDTH - 1),
		12439 => to_unsigned(30451, LUT_AMPL_WIDTH - 1),
		12440 => to_unsigned(30452, LUT_AMPL_WIDTH - 1),
		12441 => to_unsigned(30453, LUT_AMPL_WIDTH - 1),
		12442 => to_unsigned(30455, LUT_AMPL_WIDTH - 1),
		12443 => to_unsigned(30456, LUT_AMPL_WIDTH - 1),
		12444 => to_unsigned(30457, LUT_AMPL_WIDTH - 1),
		12445 => to_unsigned(30458, LUT_AMPL_WIDTH - 1),
		12446 => to_unsigned(30459, LUT_AMPL_WIDTH - 1),
		12447 => to_unsigned(30460, LUT_AMPL_WIDTH - 1),
		12448 => to_unsigned(30462, LUT_AMPL_WIDTH - 1),
		12449 => to_unsigned(30463, LUT_AMPL_WIDTH - 1),
		12450 => to_unsigned(30464, LUT_AMPL_WIDTH - 1),
		12451 => to_unsigned(30465, LUT_AMPL_WIDTH - 1),
		12452 => to_unsigned(30466, LUT_AMPL_WIDTH - 1),
		12453 => to_unsigned(30467, LUT_AMPL_WIDTH - 1),
		12454 => to_unsigned(30468, LUT_AMPL_WIDTH - 1),
		12455 => to_unsigned(30470, LUT_AMPL_WIDTH - 1),
		12456 => to_unsigned(30471, LUT_AMPL_WIDTH - 1),
		12457 => to_unsigned(30472, LUT_AMPL_WIDTH - 1),
		12458 => to_unsigned(30473, LUT_AMPL_WIDTH - 1),
		12459 => to_unsigned(30474, LUT_AMPL_WIDTH - 1),
		12460 => to_unsigned(30475, LUT_AMPL_WIDTH - 1),
		12461 => to_unsigned(30477, LUT_AMPL_WIDTH - 1),
		12462 => to_unsigned(30478, LUT_AMPL_WIDTH - 1),
		12463 => to_unsigned(30479, LUT_AMPL_WIDTH - 1),
		12464 => to_unsigned(30480, LUT_AMPL_WIDTH - 1),
		12465 => to_unsigned(30481, LUT_AMPL_WIDTH - 1),
		12466 => to_unsigned(30482, LUT_AMPL_WIDTH - 1),
		12467 => to_unsigned(30483, LUT_AMPL_WIDTH - 1),
		12468 => to_unsigned(30485, LUT_AMPL_WIDTH - 1),
		12469 => to_unsigned(30486, LUT_AMPL_WIDTH - 1),
		12470 => to_unsigned(30487, LUT_AMPL_WIDTH - 1),
		12471 => to_unsigned(30488, LUT_AMPL_WIDTH - 1),
		12472 => to_unsigned(30489, LUT_AMPL_WIDTH - 1),
		12473 => to_unsigned(30490, LUT_AMPL_WIDTH - 1),
		12474 => to_unsigned(30492, LUT_AMPL_WIDTH - 1),
		12475 => to_unsigned(30493, LUT_AMPL_WIDTH - 1),
		12476 => to_unsigned(30494, LUT_AMPL_WIDTH - 1),
		12477 => to_unsigned(30495, LUT_AMPL_WIDTH - 1),
		12478 => to_unsigned(30496, LUT_AMPL_WIDTH - 1),
		12479 => to_unsigned(30497, LUT_AMPL_WIDTH - 1),
		12480 => to_unsigned(30498, LUT_AMPL_WIDTH - 1),
		12481 => to_unsigned(30500, LUT_AMPL_WIDTH - 1),
		12482 => to_unsigned(30501, LUT_AMPL_WIDTH - 1),
		12483 => to_unsigned(30502, LUT_AMPL_WIDTH - 1),
		12484 => to_unsigned(30503, LUT_AMPL_WIDTH - 1),
		12485 => to_unsigned(30504, LUT_AMPL_WIDTH - 1),
		12486 => to_unsigned(30505, LUT_AMPL_WIDTH - 1),
		12487 => to_unsigned(30506, LUT_AMPL_WIDTH - 1),
		12488 => to_unsigned(30508, LUT_AMPL_WIDTH - 1),
		12489 => to_unsigned(30509, LUT_AMPL_WIDTH - 1),
		12490 => to_unsigned(30510, LUT_AMPL_WIDTH - 1),
		12491 => to_unsigned(30511, LUT_AMPL_WIDTH - 1),
		12492 => to_unsigned(30512, LUT_AMPL_WIDTH - 1),
		12493 => to_unsigned(30513, LUT_AMPL_WIDTH - 1),
		12494 => to_unsigned(30514, LUT_AMPL_WIDTH - 1),
		12495 => to_unsigned(30516, LUT_AMPL_WIDTH - 1),
		12496 => to_unsigned(30517, LUT_AMPL_WIDTH - 1),
		12497 => to_unsigned(30518, LUT_AMPL_WIDTH - 1),
		12498 => to_unsigned(30519, LUT_AMPL_WIDTH - 1),
		12499 => to_unsigned(30520, LUT_AMPL_WIDTH - 1),
		12500 => to_unsigned(30521, LUT_AMPL_WIDTH - 1),
		12501 => to_unsigned(30522, LUT_AMPL_WIDTH - 1),
		12502 => to_unsigned(30524, LUT_AMPL_WIDTH - 1),
		12503 => to_unsigned(30525, LUT_AMPL_WIDTH - 1),
		12504 => to_unsigned(30526, LUT_AMPL_WIDTH - 1),
		12505 => to_unsigned(30527, LUT_AMPL_WIDTH - 1),
		12506 => to_unsigned(30528, LUT_AMPL_WIDTH - 1),
		12507 => to_unsigned(30529, LUT_AMPL_WIDTH - 1),
		12508 => to_unsigned(30530, LUT_AMPL_WIDTH - 1),
		12509 => to_unsigned(30532, LUT_AMPL_WIDTH - 1),
		12510 => to_unsigned(30533, LUT_AMPL_WIDTH - 1),
		12511 => to_unsigned(30534, LUT_AMPL_WIDTH - 1),
		12512 => to_unsigned(30535, LUT_AMPL_WIDTH - 1),
		12513 => to_unsigned(30536, LUT_AMPL_WIDTH - 1),
		12514 => to_unsigned(30537, LUT_AMPL_WIDTH - 1),
		12515 => to_unsigned(30538, LUT_AMPL_WIDTH - 1),
		12516 => to_unsigned(30540, LUT_AMPL_WIDTH - 1),
		12517 => to_unsigned(30541, LUT_AMPL_WIDTH - 1),
		12518 => to_unsigned(30542, LUT_AMPL_WIDTH - 1),
		12519 => to_unsigned(30543, LUT_AMPL_WIDTH - 1),
		12520 => to_unsigned(30544, LUT_AMPL_WIDTH - 1),
		12521 => to_unsigned(30545, LUT_AMPL_WIDTH - 1),
		12522 => to_unsigned(30546, LUT_AMPL_WIDTH - 1),
		12523 => to_unsigned(30548, LUT_AMPL_WIDTH - 1),
		12524 => to_unsigned(30549, LUT_AMPL_WIDTH - 1),
		12525 => to_unsigned(30550, LUT_AMPL_WIDTH - 1),
		12526 => to_unsigned(30551, LUT_AMPL_WIDTH - 1),
		12527 => to_unsigned(30552, LUT_AMPL_WIDTH - 1),
		12528 => to_unsigned(30553, LUT_AMPL_WIDTH - 1),
		12529 => to_unsigned(30554, LUT_AMPL_WIDTH - 1),
		12530 => to_unsigned(30556, LUT_AMPL_WIDTH - 1),
		12531 => to_unsigned(30557, LUT_AMPL_WIDTH - 1),
		12532 => to_unsigned(30558, LUT_AMPL_WIDTH - 1),
		12533 => to_unsigned(30559, LUT_AMPL_WIDTH - 1),
		12534 => to_unsigned(30560, LUT_AMPL_WIDTH - 1),
		12535 => to_unsigned(30561, LUT_AMPL_WIDTH - 1),
		12536 => to_unsigned(30562, LUT_AMPL_WIDTH - 1),
		12537 => to_unsigned(30563, LUT_AMPL_WIDTH - 1),
		12538 => to_unsigned(30565, LUT_AMPL_WIDTH - 1),
		12539 => to_unsigned(30566, LUT_AMPL_WIDTH - 1),
		12540 => to_unsigned(30567, LUT_AMPL_WIDTH - 1),
		12541 => to_unsigned(30568, LUT_AMPL_WIDTH - 1),
		12542 => to_unsigned(30569, LUT_AMPL_WIDTH - 1),
		12543 => to_unsigned(30570, LUT_AMPL_WIDTH - 1),
		12544 => to_unsigned(30571, LUT_AMPL_WIDTH - 1),
		12545 => to_unsigned(30573, LUT_AMPL_WIDTH - 1),
		12546 => to_unsigned(30574, LUT_AMPL_WIDTH - 1),
		12547 => to_unsigned(30575, LUT_AMPL_WIDTH - 1),
		12548 => to_unsigned(30576, LUT_AMPL_WIDTH - 1),
		12549 => to_unsigned(30577, LUT_AMPL_WIDTH - 1),
		12550 => to_unsigned(30578, LUT_AMPL_WIDTH - 1),
		12551 => to_unsigned(30579, LUT_AMPL_WIDTH - 1),
		12552 => to_unsigned(30580, LUT_AMPL_WIDTH - 1),
		12553 => to_unsigned(30582, LUT_AMPL_WIDTH - 1),
		12554 => to_unsigned(30583, LUT_AMPL_WIDTH - 1),
		12555 => to_unsigned(30584, LUT_AMPL_WIDTH - 1),
		12556 => to_unsigned(30585, LUT_AMPL_WIDTH - 1),
		12557 => to_unsigned(30586, LUT_AMPL_WIDTH - 1),
		12558 => to_unsigned(30587, LUT_AMPL_WIDTH - 1),
		12559 => to_unsigned(30588, LUT_AMPL_WIDTH - 1),
		12560 => to_unsigned(30589, LUT_AMPL_WIDTH - 1),
		12561 => to_unsigned(30591, LUT_AMPL_WIDTH - 1),
		12562 => to_unsigned(30592, LUT_AMPL_WIDTH - 1),
		12563 => to_unsigned(30593, LUT_AMPL_WIDTH - 1),
		12564 => to_unsigned(30594, LUT_AMPL_WIDTH - 1),
		12565 => to_unsigned(30595, LUT_AMPL_WIDTH - 1),
		12566 => to_unsigned(30596, LUT_AMPL_WIDTH - 1),
		12567 => to_unsigned(30597, LUT_AMPL_WIDTH - 1),
		12568 => to_unsigned(30598, LUT_AMPL_WIDTH - 1),
		12569 => to_unsigned(30600, LUT_AMPL_WIDTH - 1),
		12570 => to_unsigned(30601, LUT_AMPL_WIDTH - 1),
		12571 => to_unsigned(30602, LUT_AMPL_WIDTH - 1),
		12572 => to_unsigned(30603, LUT_AMPL_WIDTH - 1),
		12573 => to_unsigned(30604, LUT_AMPL_WIDTH - 1),
		12574 => to_unsigned(30605, LUT_AMPL_WIDTH - 1),
		12575 => to_unsigned(30606, LUT_AMPL_WIDTH - 1),
		12576 => to_unsigned(30607, LUT_AMPL_WIDTH - 1),
		12577 => to_unsigned(30609, LUT_AMPL_WIDTH - 1),
		12578 => to_unsigned(30610, LUT_AMPL_WIDTH - 1),
		12579 => to_unsigned(30611, LUT_AMPL_WIDTH - 1),
		12580 => to_unsigned(30612, LUT_AMPL_WIDTH - 1),
		12581 => to_unsigned(30613, LUT_AMPL_WIDTH - 1),
		12582 => to_unsigned(30614, LUT_AMPL_WIDTH - 1),
		12583 => to_unsigned(30615, LUT_AMPL_WIDTH - 1),
		12584 => to_unsigned(30616, LUT_AMPL_WIDTH - 1),
		12585 => to_unsigned(30617, LUT_AMPL_WIDTH - 1),
		12586 => to_unsigned(30619, LUT_AMPL_WIDTH - 1),
		12587 => to_unsigned(30620, LUT_AMPL_WIDTH - 1),
		12588 => to_unsigned(30621, LUT_AMPL_WIDTH - 1),
		12589 => to_unsigned(30622, LUT_AMPL_WIDTH - 1),
		12590 => to_unsigned(30623, LUT_AMPL_WIDTH - 1),
		12591 => to_unsigned(30624, LUT_AMPL_WIDTH - 1),
		12592 => to_unsigned(30625, LUT_AMPL_WIDTH - 1),
		12593 => to_unsigned(30626, LUT_AMPL_WIDTH - 1),
		12594 => to_unsigned(30628, LUT_AMPL_WIDTH - 1),
		12595 => to_unsigned(30629, LUT_AMPL_WIDTH - 1),
		12596 => to_unsigned(30630, LUT_AMPL_WIDTH - 1),
		12597 => to_unsigned(30631, LUT_AMPL_WIDTH - 1),
		12598 => to_unsigned(30632, LUT_AMPL_WIDTH - 1),
		12599 => to_unsigned(30633, LUT_AMPL_WIDTH - 1),
		12600 => to_unsigned(30634, LUT_AMPL_WIDTH - 1),
		12601 => to_unsigned(30635, LUT_AMPL_WIDTH - 1),
		12602 => to_unsigned(30636, LUT_AMPL_WIDTH - 1),
		12603 => to_unsigned(30638, LUT_AMPL_WIDTH - 1),
		12604 => to_unsigned(30639, LUT_AMPL_WIDTH - 1),
		12605 => to_unsigned(30640, LUT_AMPL_WIDTH - 1),
		12606 => to_unsigned(30641, LUT_AMPL_WIDTH - 1),
		12607 => to_unsigned(30642, LUT_AMPL_WIDTH - 1),
		12608 => to_unsigned(30643, LUT_AMPL_WIDTH - 1),
		12609 => to_unsigned(30644, LUT_AMPL_WIDTH - 1),
		12610 => to_unsigned(30645, LUT_AMPL_WIDTH - 1),
		12611 => to_unsigned(30646, LUT_AMPL_WIDTH - 1),
		12612 => to_unsigned(30648, LUT_AMPL_WIDTH - 1),
		12613 => to_unsigned(30649, LUT_AMPL_WIDTH - 1),
		12614 => to_unsigned(30650, LUT_AMPL_WIDTH - 1),
		12615 => to_unsigned(30651, LUT_AMPL_WIDTH - 1),
		12616 => to_unsigned(30652, LUT_AMPL_WIDTH - 1),
		12617 => to_unsigned(30653, LUT_AMPL_WIDTH - 1),
		12618 => to_unsigned(30654, LUT_AMPL_WIDTH - 1),
		12619 => to_unsigned(30655, LUT_AMPL_WIDTH - 1),
		12620 => to_unsigned(30656, LUT_AMPL_WIDTH - 1),
		12621 => to_unsigned(30658, LUT_AMPL_WIDTH - 1),
		12622 => to_unsigned(30659, LUT_AMPL_WIDTH - 1),
		12623 => to_unsigned(30660, LUT_AMPL_WIDTH - 1),
		12624 => to_unsigned(30661, LUT_AMPL_WIDTH - 1),
		12625 => to_unsigned(30662, LUT_AMPL_WIDTH - 1),
		12626 => to_unsigned(30663, LUT_AMPL_WIDTH - 1),
		12627 => to_unsigned(30664, LUT_AMPL_WIDTH - 1),
		12628 => to_unsigned(30665, LUT_AMPL_WIDTH - 1),
		12629 => to_unsigned(30666, LUT_AMPL_WIDTH - 1),
		12630 => to_unsigned(30668, LUT_AMPL_WIDTH - 1),
		12631 => to_unsigned(30669, LUT_AMPL_WIDTH - 1),
		12632 => to_unsigned(30670, LUT_AMPL_WIDTH - 1),
		12633 => to_unsigned(30671, LUT_AMPL_WIDTH - 1),
		12634 => to_unsigned(30672, LUT_AMPL_WIDTH - 1),
		12635 => to_unsigned(30673, LUT_AMPL_WIDTH - 1),
		12636 => to_unsigned(30674, LUT_AMPL_WIDTH - 1),
		12637 => to_unsigned(30675, LUT_AMPL_WIDTH - 1),
		12638 => to_unsigned(30676, LUT_AMPL_WIDTH - 1),
		12639 => to_unsigned(30678, LUT_AMPL_WIDTH - 1),
		12640 => to_unsigned(30679, LUT_AMPL_WIDTH - 1),
		12641 => to_unsigned(30680, LUT_AMPL_WIDTH - 1),
		12642 => to_unsigned(30681, LUT_AMPL_WIDTH - 1),
		12643 => to_unsigned(30682, LUT_AMPL_WIDTH - 1),
		12644 => to_unsigned(30683, LUT_AMPL_WIDTH - 1),
		12645 => to_unsigned(30684, LUT_AMPL_WIDTH - 1),
		12646 => to_unsigned(30685, LUT_AMPL_WIDTH - 1),
		12647 => to_unsigned(30686, LUT_AMPL_WIDTH - 1),
		12648 => to_unsigned(30687, LUT_AMPL_WIDTH - 1),
		12649 => to_unsigned(30689, LUT_AMPL_WIDTH - 1),
		12650 => to_unsigned(30690, LUT_AMPL_WIDTH - 1),
		12651 => to_unsigned(30691, LUT_AMPL_WIDTH - 1),
		12652 => to_unsigned(30692, LUT_AMPL_WIDTH - 1),
		12653 => to_unsigned(30693, LUT_AMPL_WIDTH - 1),
		12654 => to_unsigned(30694, LUT_AMPL_WIDTH - 1),
		12655 => to_unsigned(30695, LUT_AMPL_WIDTH - 1),
		12656 => to_unsigned(30696, LUT_AMPL_WIDTH - 1),
		12657 => to_unsigned(30697, LUT_AMPL_WIDTH - 1),
		12658 => to_unsigned(30698, LUT_AMPL_WIDTH - 1),
		12659 => to_unsigned(30700, LUT_AMPL_WIDTH - 1),
		12660 => to_unsigned(30701, LUT_AMPL_WIDTH - 1),
		12661 => to_unsigned(30702, LUT_AMPL_WIDTH - 1),
		12662 => to_unsigned(30703, LUT_AMPL_WIDTH - 1),
		12663 => to_unsigned(30704, LUT_AMPL_WIDTH - 1),
		12664 => to_unsigned(30705, LUT_AMPL_WIDTH - 1),
		12665 => to_unsigned(30706, LUT_AMPL_WIDTH - 1),
		12666 => to_unsigned(30707, LUT_AMPL_WIDTH - 1),
		12667 => to_unsigned(30708, LUT_AMPL_WIDTH - 1),
		12668 => to_unsigned(30709, LUT_AMPL_WIDTH - 1),
		12669 => to_unsigned(30711, LUT_AMPL_WIDTH - 1),
		12670 => to_unsigned(30712, LUT_AMPL_WIDTH - 1),
		12671 => to_unsigned(30713, LUT_AMPL_WIDTH - 1),
		12672 => to_unsigned(30714, LUT_AMPL_WIDTH - 1),
		12673 => to_unsigned(30715, LUT_AMPL_WIDTH - 1),
		12674 => to_unsigned(30716, LUT_AMPL_WIDTH - 1),
		12675 => to_unsigned(30717, LUT_AMPL_WIDTH - 1),
		12676 => to_unsigned(30718, LUT_AMPL_WIDTH - 1),
		12677 => to_unsigned(30719, LUT_AMPL_WIDTH - 1),
		12678 => to_unsigned(30720, LUT_AMPL_WIDTH - 1),
		12679 => to_unsigned(30721, LUT_AMPL_WIDTH - 1),
		12680 => to_unsigned(30723, LUT_AMPL_WIDTH - 1),
		12681 => to_unsigned(30724, LUT_AMPL_WIDTH - 1),
		12682 => to_unsigned(30725, LUT_AMPL_WIDTH - 1),
		12683 => to_unsigned(30726, LUT_AMPL_WIDTH - 1),
		12684 => to_unsigned(30727, LUT_AMPL_WIDTH - 1),
		12685 => to_unsigned(30728, LUT_AMPL_WIDTH - 1),
		12686 => to_unsigned(30729, LUT_AMPL_WIDTH - 1),
		12687 => to_unsigned(30730, LUT_AMPL_WIDTH - 1),
		12688 => to_unsigned(30731, LUT_AMPL_WIDTH - 1),
		12689 => to_unsigned(30732, LUT_AMPL_WIDTH - 1),
		12690 => to_unsigned(30733, LUT_AMPL_WIDTH - 1),
		12691 => to_unsigned(30735, LUT_AMPL_WIDTH - 1),
		12692 => to_unsigned(30736, LUT_AMPL_WIDTH - 1),
		12693 => to_unsigned(30737, LUT_AMPL_WIDTH - 1),
		12694 => to_unsigned(30738, LUT_AMPL_WIDTH - 1),
		12695 => to_unsigned(30739, LUT_AMPL_WIDTH - 1),
		12696 => to_unsigned(30740, LUT_AMPL_WIDTH - 1),
		12697 => to_unsigned(30741, LUT_AMPL_WIDTH - 1),
		12698 => to_unsigned(30742, LUT_AMPL_WIDTH - 1),
		12699 => to_unsigned(30743, LUT_AMPL_WIDTH - 1),
		12700 => to_unsigned(30744, LUT_AMPL_WIDTH - 1),
		12701 => to_unsigned(30745, LUT_AMPL_WIDTH - 1),
		12702 => to_unsigned(30746, LUT_AMPL_WIDTH - 1),
		12703 => to_unsigned(30748, LUT_AMPL_WIDTH - 1),
		12704 => to_unsigned(30749, LUT_AMPL_WIDTH - 1),
		12705 => to_unsigned(30750, LUT_AMPL_WIDTH - 1),
		12706 => to_unsigned(30751, LUT_AMPL_WIDTH - 1),
		12707 => to_unsigned(30752, LUT_AMPL_WIDTH - 1),
		12708 => to_unsigned(30753, LUT_AMPL_WIDTH - 1),
		12709 => to_unsigned(30754, LUT_AMPL_WIDTH - 1),
		12710 => to_unsigned(30755, LUT_AMPL_WIDTH - 1),
		12711 => to_unsigned(30756, LUT_AMPL_WIDTH - 1),
		12712 => to_unsigned(30757, LUT_AMPL_WIDTH - 1),
		12713 => to_unsigned(30758, LUT_AMPL_WIDTH - 1),
		12714 => to_unsigned(30760, LUT_AMPL_WIDTH - 1),
		12715 => to_unsigned(30761, LUT_AMPL_WIDTH - 1),
		12716 => to_unsigned(30762, LUT_AMPL_WIDTH - 1),
		12717 => to_unsigned(30763, LUT_AMPL_WIDTH - 1),
		12718 => to_unsigned(30764, LUT_AMPL_WIDTH - 1),
		12719 => to_unsigned(30765, LUT_AMPL_WIDTH - 1),
		12720 => to_unsigned(30766, LUT_AMPL_WIDTH - 1),
		12721 => to_unsigned(30767, LUT_AMPL_WIDTH - 1),
		12722 => to_unsigned(30768, LUT_AMPL_WIDTH - 1),
		12723 => to_unsigned(30769, LUT_AMPL_WIDTH - 1),
		12724 => to_unsigned(30770, LUT_AMPL_WIDTH - 1),
		12725 => to_unsigned(30771, LUT_AMPL_WIDTH - 1),
		12726 => to_unsigned(30772, LUT_AMPL_WIDTH - 1),
		12727 => to_unsigned(30774, LUT_AMPL_WIDTH - 1),
		12728 => to_unsigned(30775, LUT_AMPL_WIDTH - 1),
		12729 => to_unsigned(30776, LUT_AMPL_WIDTH - 1),
		12730 => to_unsigned(30777, LUT_AMPL_WIDTH - 1),
		12731 => to_unsigned(30778, LUT_AMPL_WIDTH - 1),
		12732 => to_unsigned(30779, LUT_AMPL_WIDTH - 1),
		12733 => to_unsigned(30780, LUT_AMPL_WIDTH - 1),
		12734 => to_unsigned(30781, LUT_AMPL_WIDTH - 1),
		12735 => to_unsigned(30782, LUT_AMPL_WIDTH - 1),
		12736 => to_unsigned(30783, LUT_AMPL_WIDTH - 1),
		12737 => to_unsigned(30784, LUT_AMPL_WIDTH - 1),
		12738 => to_unsigned(30785, LUT_AMPL_WIDTH - 1),
		12739 => to_unsigned(30786, LUT_AMPL_WIDTH - 1),
		12740 => to_unsigned(30788, LUT_AMPL_WIDTH - 1),
		12741 => to_unsigned(30789, LUT_AMPL_WIDTH - 1),
		12742 => to_unsigned(30790, LUT_AMPL_WIDTH - 1),
		12743 => to_unsigned(30791, LUT_AMPL_WIDTH - 1),
		12744 => to_unsigned(30792, LUT_AMPL_WIDTH - 1),
		12745 => to_unsigned(30793, LUT_AMPL_WIDTH - 1),
		12746 => to_unsigned(30794, LUT_AMPL_WIDTH - 1),
		12747 => to_unsigned(30795, LUT_AMPL_WIDTH - 1),
		12748 => to_unsigned(30796, LUT_AMPL_WIDTH - 1),
		12749 => to_unsigned(30797, LUT_AMPL_WIDTH - 1),
		12750 => to_unsigned(30798, LUT_AMPL_WIDTH - 1),
		12751 => to_unsigned(30799, LUT_AMPL_WIDTH - 1),
		12752 => to_unsigned(30800, LUT_AMPL_WIDTH - 1),
		12753 => to_unsigned(30802, LUT_AMPL_WIDTH - 1),
		12754 => to_unsigned(30803, LUT_AMPL_WIDTH - 1),
		12755 => to_unsigned(30804, LUT_AMPL_WIDTH - 1),
		12756 => to_unsigned(30805, LUT_AMPL_WIDTH - 1),
		12757 => to_unsigned(30806, LUT_AMPL_WIDTH - 1),
		12758 => to_unsigned(30807, LUT_AMPL_WIDTH - 1),
		12759 => to_unsigned(30808, LUT_AMPL_WIDTH - 1),
		12760 => to_unsigned(30809, LUT_AMPL_WIDTH - 1),
		12761 => to_unsigned(30810, LUT_AMPL_WIDTH - 1),
		12762 => to_unsigned(30811, LUT_AMPL_WIDTH - 1),
		12763 => to_unsigned(30812, LUT_AMPL_WIDTH - 1),
		12764 => to_unsigned(30813, LUT_AMPL_WIDTH - 1),
		12765 => to_unsigned(30814, LUT_AMPL_WIDTH - 1),
		12766 => to_unsigned(30815, LUT_AMPL_WIDTH - 1),
		12767 => to_unsigned(30816, LUT_AMPL_WIDTH - 1),
		12768 => to_unsigned(30818, LUT_AMPL_WIDTH - 1),
		12769 => to_unsigned(30819, LUT_AMPL_WIDTH - 1),
		12770 => to_unsigned(30820, LUT_AMPL_WIDTH - 1),
		12771 => to_unsigned(30821, LUT_AMPL_WIDTH - 1),
		12772 => to_unsigned(30822, LUT_AMPL_WIDTH - 1),
		12773 => to_unsigned(30823, LUT_AMPL_WIDTH - 1),
		12774 => to_unsigned(30824, LUT_AMPL_WIDTH - 1),
		12775 => to_unsigned(30825, LUT_AMPL_WIDTH - 1),
		12776 => to_unsigned(30826, LUT_AMPL_WIDTH - 1),
		12777 => to_unsigned(30827, LUT_AMPL_WIDTH - 1),
		12778 => to_unsigned(30828, LUT_AMPL_WIDTH - 1),
		12779 => to_unsigned(30829, LUT_AMPL_WIDTH - 1),
		12780 => to_unsigned(30830, LUT_AMPL_WIDTH - 1),
		12781 => to_unsigned(30831, LUT_AMPL_WIDTH - 1),
		12782 => to_unsigned(30832, LUT_AMPL_WIDTH - 1),
		12783 => to_unsigned(30834, LUT_AMPL_WIDTH - 1),
		12784 => to_unsigned(30835, LUT_AMPL_WIDTH - 1),
		12785 => to_unsigned(30836, LUT_AMPL_WIDTH - 1),
		12786 => to_unsigned(30837, LUT_AMPL_WIDTH - 1),
		12787 => to_unsigned(30838, LUT_AMPL_WIDTH - 1),
		12788 => to_unsigned(30839, LUT_AMPL_WIDTH - 1),
		12789 => to_unsigned(30840, LUT_AMPL_WIDTH - 1),
		12790 => to_unsigned(30841, LUT_AMPL_WIDTH - 1),
		12791 => to_unsigned(30842, LUT_AMPL_WIDTH - 1),
		12792 => to_unsigned(30843, LUT_AMPL_WIDTH - 1),
		12793 => to_unsigned(30844, LUT_AMPL_WIDTH - 1),
		12794 => to_unsigned(30845, LUT_AMPL_WIDTH - 1),
		12795 => to_unsigned(30846, LUT_AMPL_WIDTH - 1),
		12796 => to_unsigned(30847, LUT_AMPL_WIDTH - 1),
		12797 => to_unsigned(30848, LUT_AMPL_WIDTH - 1),
		12798 => to_unsigned(30849, LUT_AMPL_WIDTH - 1),
		12799 => to_unsigned(30851, LUT_AMPL_WIDTH - 1),
		12800 => to_unsigned(30852, LUT_AMPL_WIDTH - 1),
		12801 => to_unsigned(30853, LUT_AMPL_WIDTH - 1),
		12802 => to_unsigned(30854, LUT_AMPL_WIDTH - 1),
		12803 => to_unsigned(30855, LUT_AMPL_WIDTH - 1),
		12804 => to_unsigned(30856, LUT_AMPL_WIDTH - 1),
		12805 => to_unsigned(30857, LUT_AMPL_WIDTH - 1),
		12806 => to_unsigned(30858, LUT_AMPL_WIDTH - 1),
		12807 => to_unsigned(30859, LUT_AMPL_WIDTH - 1),
		12808 => to_unsigned(30860, LUT_AMPL_WIDTH - 1),
		12809 => to_unsigned(30861, LUT_AMPL_WIDTH - 1),
		12810 => to_unsigned(30862, LUT_AMPL_WIDTH - 1),
		12811 => to_unsigned(30863, LUT_AMPL_WIDTH - 1),
		12812 => to_unsigned(30864, LUT_AMPL_WIDTH - 1),
		12813 => to_unsigned(30865, LUT_AMPL_WIDTH - 1),
		12814 => to_unsigned(30866, LUT_AMPL_WIDTH - 1),
		12815 => to_unsigned(30867, LUT_AMPL_WIDTH - 1),
		12816 => to_unsigned(30868, LUT_AMPL_WIDTH - 1),
		12817 => to_unsigned(30870, LUT_AMPL_WIDTH - 1),
		12818 => to_unsigned(30871, LUT_AMPL_WIDTH - 1),
		12819 => to_unsigned(30872, LUT_AMPL_WIDTH - 1),
		12820 => to_unsigned(30873, LUT_AMPL_WIDTH - 1),
		12821 => to_unsigned(30874, LUT_AMPL_WIDTH - 1),
		12822 => to_unsigned(30875, LUT_AMPL_WIDTH - 1),
		12823 => to_unsigned(30876, LUT_AMPL_WIDTH - 1),
		12824 => to_unsigned(30877, LUT_AMPL_WIDTH - 1),
		12825 => to_unsigned(30878, LUT_AMPL_WIDTH - 1),
		12826 => to_unsigned(30879, LUT_AMPL_WIDTH - 1),
		12827 => to_unsigned(30880, LUT_AMPL_WIDTH - 1),
		12828 => to_unsigned(30881, LUT_AMPL_WIDTH - 1),
		12829 => to_unsigned(30882, LUT_AMPL_WIDTH - 1),
		12830 => to_unsigned(30883, LUT_AMPL_WIDTH - 1),
		12831 => to_unsigned(30884, LUT_AMPL_WIDTH - 1),
		12832 => to_unsigned(30885, LUT_AMPL_WIDTH - 1),
		12833 => to_unsigned(30886, LUT_AMPL_WIDTH - 1),
		12834 => to_unsigned(30887, LUT_AMPL_WIDTH - 1),
		12835 => to_unsigned(30888, LUT_AMPL_WIDTH - 1),
		12836 => to_unsigned(30889, LUT_AMPL_WIDTH - 1),
		12837 => to_unsigned(30891, LUT_AMPL_WIDTH - 1),
		12838 => to_unsigned(30892, LUT_AMPL_WIDTH - 1),
		12839 => to_unsigned(30893, LUT_AMPL_WIDTH - 1),
		12840 => to_unsigned(30894, LUT_AMPL_WIDTH - 1),
		12841 => to_unsigned(30895, LUT_AMPL_WIDTH - 1),
		12842 => to_unsigned(30896, LUT_AMPL_WIDTH - 1),
		12843 => to_unsigned(30897, LUT_AMPL_WIDTH - 1),
		12844 => to_unsigned(30898, LUT_AMPL_WIDTH - 1),
		12845 => to_unsigned(30899, LUT_AMPL_WIDTH - 1),
		12846 => to_unsigned(30900, LUT_AMPL_WIDTH - 1),
		12847 => to_unsigned(30901, LUT_AMPL_WIDTH - 1),
		12848 => to_unsigned(30902, LUT_AMPL_WIDTH - 1),
		12849 => to_unsigned(30903, LUT_AMPL_WIDTH - 1),
		12850 => to_unsigned(30904, LUT_AMPL_WIDTH - 1),
		12851 => to_unsigned(30905, LUT_AMPL_WIDTH - 1),
		12852 => to_unsigned(30906, LUT_AMPL_WIDTH - 1),
		12853 => to_unsigned(30907, LUT_AMPL_WIDTH - 1),
		12854 => to_unsigned(30908, LUT_AMPL_WIDTH - 1),
		12855 => to_unsigned(30909, LUT_AMPL_WIDTH - 1),
		12856 => to_unsigned(30910, LUT_AMPL_WIDTH - 1),
		12857 => to_unsigned(30911, LUT_AMPL_WIDTH - 1),
		12858 => to_unsigned(30912, LUT_AMPL_WIDTH - 1),
		12859 => to_unsigned(30914, LUT_AMPL_WIDTH - 1),
		12860 => to_unsigned(30915, LUT_AMPL_WIDTH - 1),
		12861 => to_unsigned(30916, LUT_AMPL_WIDTH - 1),
		12862 => to_unsigned(30917, LUT_AMPL_WIDTH - 1),
		12863 => to_unsigned(30918, LUT_AMPL_WIDTH - 1),
		12864 => to_unsigned(30919, LUT_AMPL_WIDTH - 1),
		12865 => to_unsigned(30920, LUT_AMPL_WIDTH - 1),
		12866 => to_unsigned(30921, LUT_AMPL_WIDTH - 1),
		12867 => to_unsigned(30922, LUT_AMPL_WIDTH - 1),
		12868 => to_unsigned(30923, LUT_AMPL_WIDTH - 1),
		12869 => to_unsigned(30924, LUT_AMPL_WIDTH - 1),
		12870 => to_unsigned(30925, LUT_AMPL_WIDTH - 1),
		12871 => to_unsigned(30926, LUT_AMPL_WIDTH - 1),
		12872 => to_unsigned(30927, LUT_AMPL_WIDTH - 1),
		12873 => to_unsigned(30928, LUT_AMPL_WIDTH - 1),
		12874 => to_unsigned(30929, LUT_AMPL_WIDTH - 1),
		12875 => to_unsigned(30930, LUT_AMPL_WIDTH - 1),
		12876 => to_unsigned(30931, LUT_AMPL_WIDTH - 1),
		12877 => to_unsigned(30932, LUT_AMPL_WIDTH - 1),
		12878 => to_unsigned(30933, LUT_AMPL_WIDTH - 1),
		12879 => to_unsigned(30934, LUT_AMPL_WIDTH - 1),
		12880 => to_unsigned(30935, LUT_AMPL_WIDTH - 1),
		12881 => to_unsigned(30936, LUT_AMPL_WIDTH - 1),
		12882 => to_unsigned(30937, LUT_AMPL_WIDTH - 1),
		12883 => to_unsigned(30938, LUT_AMPL_WIDTH - 1),
		12884 => to_unsigned(30939, LUT_AMPL_WIDTH - 1),
		12885 => to_unsigned(30941, LUT_AMPL_WIDTH - 1),
		12886 => to_unsigned(30942, LUT_AMPL_WIDTH - 1),
		12887 => to_unsigned(30943, LUT_AMPL_WIDTH - 1),
		12888 => to_unsigned(30944, LUT_AMPL_WIDTH - 1),
		12889 => to_unsigned(30945, LUT_AMPL_WIDTH - 1),
		12890 => to_unsigned(30946, LUT_AMPL_WIDTH - 1),
		12891 => to_unsigned(30947, LUT_AMPL_WIDTH - 1),
		12892 => to_unsigned(30948, LUT_AMPL_WIDTH - 1),
		12893 => to_unsigned(30949, LUT_AMPL_WIDTH - 1),
		12894 => to_unsigned(30950, LUT_AMPL_WIDTH - 1),
		12895 => to_unsigned(30951, LUT_AMPL_WIDTH - 1),
		12896 => to_unsigned(30952, LUT_AMPL_WIDTH - 1),
		12897 => to_unsigned(30953, LUT_AMPL_WIDTH - 1),
		12898 => to_unsigned(30954, LUT_AMPL_WIDTH - 1),
		12899 => to_unsigned(30955, LUT_AMPL_WIDTH - 1),
		12900 => to_unsigned(30956, LUT_AMPL_WIDTH - 1),
		12901 => to_unsigned(30957, LUT_AMPL_WIDTH - 1),
		12902 => to_unsigned(30958, LUT_AMPL_WIDTH - 1),
		12903 => to_unsigned(30959, LUT_AMPL_WIDTH - 1),
		12904 => to_unsigned(30960, LUT_AMPL_WIDTH - 1),
		12905 => to_unsigned(30961, LUT_AMPL_WIDTH - 1),
		12906 => to_unsigned(30962, LUT_AMPL_WIDTH - 1),
		12907 => to_unsigned(30963, LUT_AMPL_WIDTH - 1),
		12908 => to_unsigned(30964, LUT_AMPL_WIDTH - 1),
		12909 => to_unsigned(30965, LUT_AMPL_WIDTH - 1),
		12910 => to_unsigned(30966, LUT_AMPL_WIDTH - 1),
		12911 => to_unsigned(30967, LUT_AMPL_WIDTH - 1),
		12912 => to_unsigned(30968, LUT_AMPL_WIDTH - 1),
		12913 => to_unsigned(30969, LUT_AMPL_WIDTH - 1),
		12914 => to_unsigned(30970, LUT_AMPL_WIDTH - 1),
		12915 => to_unsigned(30971, LUT_AMPL_WIDTH - 1),
		12916 => to_unsigned(30972, LUT_AMPL_WIDTH - 1),
		12917 => to_unsigned(30973, LUT_AMPL_WIDTH - 1),
		12918 => to_unsigned(30974, LUT_AMPL_WIDTH - 1),
		12919 => to_unsigned(30976, LUT_AMPL_WIDTH - 1),
		12920 => to_unsigned(30977, LUT_AMPL_WIDTH - 1),
		12921 => to_unsigned(30978, LUT_AMPL_WIDTH - 1),
		12922 => to_unsigned(30979, LUT_AMPL_WIDTH - 1),
		12923 => to_unsigned(30980, LUT_AMPL_WIDTH - 1),
		12924 => to_unsigned(30981, LUT_AMPL_WIDTH - 1),
		12925 => to_unsigned(30982, LUT_AMPL_WIDTH - 1),
		12926 => to_unsigned(30983, LUT_AMPL_WIDTH - 1),
		12927 => to_unsigned(30984, LUT_AMPL_WIDTH - 1),
		12928 => to_unsigned(30985, LUT_AMPL_WIDTH - 1),
		12929 => to_unsigned(30986, LUT_AMPL_WIDTH - 1),
		12930 => to_unsigned(30987, LUT_AMPL_WIDTH - 1),
		12931 => to_unsigned(30988, LUT_AMPL_WIDTH - 1),
		12932 => to_unsigned(30989, LUT_AMPL_WIDTH - 1),
		12933 => to_unsigned(30990, LUT_AMPL_WIDTH - 1),
		12934 => to_unsigned(30991, LUT_AMPL_WIDTH - 1),
		12935 => to_unsigned(30992, LUT_AMPL_WIDTH - 1),
		12936 => to_unsigned(30993, LUT_AMPL_WIDTH - 1),
		12937 => to_unsigned(30994, LUT_AMPL_WIDTH - 1),
		12938 => to_unsigned(30995, LUT_AMPL_WIDTH - 1),
		12939 => to_unsigned(30996, LUT_AMPL_WIDTH - 1),
		12940 => to_unsigned(30997, LUT_AMPL_WIDTH - 1),
		12941 => to_unsigned(30998, LUT_AMPL_WIDTH - 1),
		12942 => to_unsigned(30999, LUT_AMPL_WIDTH - 1),
		12943 => to_unsigned(31000, LUT_AMPL_WIDTH - 1),
		12944 => to_unsigned(31001, LUT_AMPL_WIDTH - 1),
		12945 => to_unsigned(31002, LUT_AMPL_WIDTH - 1),
		12946 => to_unsigned(31003, LUT_AMPL_WIDTH - 1),
		12947 => to_unsigned(31004, LUT_AMPL_WIDTH - 1),
		12948 => to_unsigned(31005, LUT_AMPL_WIDTH - 1),
		12949 => to_unsigned(31006, LUT_AMPL_WIDTH - 1),
		12950 => to_unsigned(31007, LUT_AMPL_WIDTH - 1),
		12951 => to_unsigned(31008, LUT_AMPL_WIDTH - 1),
		12952 => to_unsigned(31009, LUT_AMPL_WIDTH - 1),
		12953 => to_unsigned(31010, LUT_AMPL_WIDTH - 1),
		12954 => to_unsigned(31011, LUT_AMPL_WIDTH - 1),
		12955 => to_unsigned(31012, LUT_AMPL_WIDTH - 1),
		12956 => to_unsigned(31013, LUT_AMPL_WIDTH - 1),
		12957 => to_unsigned(31014, LUT_AMPL_WIDTH - 1),
		12958 => to_unsigned(31015, LUT_AMPL_WIDTH - 1),
		12959 => to_unsigned(31016, LUT_AMPL_WIDTH - 1),
		12960 => to_unsigned(31017, LUT_AMPL_WIDTH - 1),
		12961 => to_unsigned(31018, LUT_AMPL_WIDTH - 1),
		12962 => to_unsigned(31019, LUT_AMPL_WIDTH - 1),
		12963 => to_unsigned(31020, LUT_AMPL_WIDTH - 1),
		12964 => to_unsigned(31021, LUT_AMPL_WIDTH - 1),
		12965 => to_unsigned(31022, LUT_AMPL_WIDTH - 1),
		12966 => to_unsigned(31023, LUT_AMPL_WIDTH - 1),
		12967 => to_unsigned(31024, LUT_AMPL_WIDTH - 1),
		12968 => to_unsigned(31025, LUT_AMPL_WIDTH - 1),
		12969 => to_unsigned(31026, LUT_AMPL_WIDTH - 1),
		12970 => to_unsigned(31027, LUT_AMPL_WIDTH - 1),
		12971 => to_unsigned(31028, LUT_AMPL_WIDTH - 1),
		12972 => to_unsigned(31029, LUT_AMPL_WIDTH - 1),
		12973 => to_unsigned(31030, LUT_AMPL_WIDTH - 1),
		12974 => to_unsigned(31031, LUT_AMPL_WIDTH - 1),
		12975 => to_unsigned(31032, LUT_AMPL_WIDTH - 1),
		12976 => to_unsigned(31033, LUT_AMPL_WIDTH - 1),
		12977 => to_unsigned(31034, LUT_AMPL_WIDTH - 1),
		12978 => to_unsigned(31035, LUT_AMPL_WIDTH - 1),
		12979 => to_unsigned(31036, LUT_AMPL_WIDTH - 1),
		12980 => to_unsigned(31037, LUT_AMPL_WIDTH - 1),
		12981 => to_unsigned(31038, LUT_AMPL_WIDTH - 1),
		12982 => to_unsigned(31039, LUT_AMPL_WIDTH - 1),
		12983 => to_unsigned(31040, LUT_AMPL_WIDTH - 1),
		12984 => to_unsigned(31041, LUT_AMPL_WIDTH - 1),
		12985 => to_unsigned(31043, LUT_AMPL_WIDTH - 1),
		12986 => to_unsigned(31044, LUT_AMPL_WIDTH - 1),
		12987 => to_unsigned(31045, LUT_AMPL_WIDTH - 1),
		12988 => to_unsigned(31046, LUT_AMPL_WIDTH - 1),
		12989 => to_unsigned(31047, LUT_AMPL_WIDTH - 1),
		12990 => to_unsigned(31048, LUT_AMPL_WIDTH - 1),
		12991 => to_unsigned(31049, LUT_AMPL_WIDTH - 1),
		12992 => to_unsigned(31050, LUT_AMPL_WIDTH - 1),
		12993 => to_unsigned(31051, LUT_AMPL_WIDTH - 1),
		12994 => to_unsigned(31052, LUT_AMPL_WIDTH - 1),
		12995 => to_unsigned(31053, LUT_AMPL_WIDTH - 1),
		12996 => to_unsigned(31054, LUT_AMPL_WIDTH - 1),
		12997 => to_unsigned(31055, LUT_AMPL_WIDTH - 1),
		12998 => to_unsigned(31056, LUT_AMPL_WIDTH - 1),
		12999 => to_unsigned(31057, LUT_AMPL_WIDTH - 1),
		13000 => to_unsigned(31058, LUT_AMPL_WIDTH - 1),
		13001 => to_unsigned(31059, LUT_AMPL_WIDTH - 1),
		13002 => to_unsigned(31060, LUT_AMPL_WIDTH - 1),
		13003 => to_unsigned(31061, LUT_AMPL_WIDTH - 1),
		13004 => to_unsigned(31062, LUT_AMPL_WIDTH - 1),
		13005 => to_unsigned(31063, LUT_AMPL_WIDTH - 1),
		13006 => to_unsigned(31064, LUT_AMPL_WIDTH - 1),
		13007 => to_unsigned(31065, LUT_AMPL_WIDTH - 1),
		13008 => to_unsigned(31066, LUT_AMPL_WIDTH - 1),
		13009 => to_unsigned(31067, LUT_AMPL_WIDTH - 1),
		13010 => to_unsigned(31068, LUT_AMPL_WIDTH - 1),
		13011 => to_unsigned(31069, LUT_AMPL_WIDTH - 1),
		13012 => to_unsigned(31070, LUT_AMPL_WIDTH - 1),
		13013 => to_unsigned(31071, LUT_AMPL_WIDTH - 1),
		13014 => to_unsigned(31072, LUT_AMPL_WIDTH - 1),
		13015 => to_unsigned(31073, LUT_AMPL_WIDTH - 1),
		13016 => to_unsigned(31074, LUT_AMPL_WIDTH - 1),
		13017 => to_unsigned(31075, LUT_AMPL_WIDTH - 1),
		13018 => to_unsigned(31076, LUT_AMPL_WIDTH - 1),
		13019 => to_unsigned(31077, LUT_AMPL_WIDTH - 1),
		13020 => to_unsigned(31078, LUT_AMPL_WIDTH - 1),
		13021 => to_unsigned(31079, LUT_AMPL_WIDTH - 1),
		13022 => to_unsigned(31080, LUT_AMPL_WIDTH - 1),
		13023 => to_unsigned(31081, LUT_AMPL_WIDTH - 1),
		13024 => to_unsigned(31082, LUT_AMPL_WIDTH - 1),
		13025 => to_unsigned(31083, LUT_AMPL_WIDTH - 1),
		13026 => to_unsigned(31083, LUT_AMPL_WIDTH - 1),
		13027 => to_unsigned(31084, LUT_AMPL_WIDTH - 1),
		13028 => to_unsigned(31085, LUT_AMPL_WIDTH - 1),
		13029 => to_unsigned(31086, LUT_AMPL_WIDTH - 1),
		13030 => to_unsigned(31087, LUT_AMPL_WIDTH - 1),
		13031 => to_unsigned(31088, LUT_AMPL_WIDTH - 1),
		13032 => to_unsigned(31089, LUT_AMPL_WIDTH - 1),
		13033 => to_unsigned(31090, LUT_AMPL_WIDTH - 1),
		13034 => to_unsigned(31091, LUT_AMPL_WIDTH - 1),
		13035 => to_unsigned(31092, LUT_AMPL_WIDTH - 1),
		13036 => to_unsigned(31093, LUT_AMPL_WIDTH - 1),
		13037 => to_unsigned(31094, LUT_AMPL_WIDTH - 1),
		13038 => to_unsigned(31095, LUT_AMPL_WIDTH - 1),
		13039 => to_unsigned(31096, LUT_AMPL_WIDTH - 1),
		13040 => to_unsigned(31097, LUT_AMPL_WIDTH - 1),
		13041 => to_unsigned(31098, LUT_AMPL_WIDTH - 1),
		13042 => to_unsigned(31099, LUT_AMPL_WIDTH - 1),
		13043 => to_unsigned(31100, LUT_AMPL_WIDTH - 1),
		13044 => to_unsigned(31101, LUT_AMPL_WIDTH - 1),
		13045 => to_unsigned(31102, LUT_AMPL_WIDTH - 1),
		13046 => to_unsigned(31103, LUT_AMPL_WIDTH - 1),
		13047 => to_unsigned(31104, LUT_AMPL_WIDTH - 1),
		13048 => to_unsigned(31105, LUT_AMPL_WIDTH - 1),
		13049 => to_unsigned(31106, LUT_AMPL_WIDTH - 1),
		13050 => to_unsigned(31107, LUT_AMPL_WIDTH - 1),
		13051 => to_unsigned(31108, LUT_AMPL_WIDTH - 1),
		13052 => to_unsigned(31109, LUT_AMPL_WIDTH - 1),
		13053 => to_unsigned(31110, LUT_AMPL_WIDTH - 1),
		13054 => to_unsigned(31111, LUT_AMPL_WIDTH - 1),
		13055 => to_unsigned(31112, LUT_AMPL_WIDTH - 1),
		13056 => to_unsigned(31113, LUT_AMPL_WIDTH - 1),
		13057 => to_unsigned(31114, LUT_AMPL_WIDTH - 1),
		13058 => to_unsigned(31115, LUT_AMPL_WIDTH - 1),
		13059 => to_unsigned(31116, LUT_AMPL_WIDTH - 1),
		13060 => to_unsigned(31117, LUT_AMPL_WIDTH - 1),
		13061 => to_unsigned(31118, LUT_AMPL_WIDTH - 1),
		13062 => to_unsigned(31119, LUT_AMPL_WIDTH - 1),
		13063 => to_unsigned(31120, LUT_AMPL_WIDTH - 1),
		13064 => to_unsigned(31121, LUT_AMPL_WIDTH - 1),
		13065 => to_unsigned(31122, LUT_AMPL_WIDTH - 1),
		13066 => to_unsigned(31123, LUT_AMPL_WIDTH - 1),
		13067 => to_unsigned(31124, LUT_AMPL_WIDTH - 1),
		13068 => to_unsigned(31125, LUT_AMPL_WIDTH - 1),
		13069 => to_unsigned(31126, LUT_AMPL_WIDTH - 1),
		13070 => to_unsigned(31127, LUT_AMPL_WIDTH - 1),
		13071 => to_unsigned(31128, LUT_AMPL_WIDTH - 1),
		13072 => to_unsigned(31129, LUT_AMPL_WIDTH - 1),
		13073 => to_unsigned(31130, LUT_AMPL_WIDTH - 1),
		13074 => to_unsigned(31131, LUT_AMPL_WIDTH - 1),
		13075 => to_unsigned(31132, LUT_AMPL_WIDTH - 1),
		13076 => to_unsigned(31133, LUT_AMPL_WIDTH - 1),
		13077 => to_unsigned(31134, LUT_AMPL_WIDTH - 1),
		13078 => to_unsigned(31135, LUT_AMPL_WIDTH - 1),
		13079 => to_unsigned(31136, LUT_AMPL_WIDTH - 1),
		13080 => to_unsigned(31137, LUT_AMPL_WIDTH - 1),
		13081 => to_unsigned(31138, LUT_AMPL_WIDTH - 1),
		13082 => to_unsigned(31139, LUT_AMPL_WIDTH - 1),
		13083 => to_unsigned(31140, LUT_AMPL_WIDTH - 1),
		13084 => to_unsigned(31141, LUT_AMPL_WIDTH - 1),
		13085 => to_unsigned(31142, LUT_AMPL_WIDTH - 1),
		13086 => to_unsigned(31143, LUT_AMPL_WIDTH - 1),
		13087 => to_unsigned(31144, LUT_AMPL_WIDTH - 1),
		13088 => to_unsigned(31145, LUT_AMPL_WIDTH - 1),
		13089 => to_unsigned(31146, LUT_AMPL_WIDTH - 1),
		13090 => to_unsigned(31147, LUT_AMPL_WIDTH - 1),
		13091 => to_unsigned(31148, LUT_AMPL_WIDTH - 1),
		13092 => to_unsigned(31148, LUT_AMPL_WIDTH - 1),
		13093 => to_unsigned(31149, LUT_AMPL_WIDTH - 1),
		13094 => to_unsigned(31150, LUT_AMPL_WIDTH - 1),
		13095 => to_unsigned(31151, LUT_AMPL_WIDTH - 1),
		13096 => to_unsigned(31152, LUT_AMPL_WIDTH - 1),
		13097 => to_unsigned(31153, LUT_AMPL_WIDTH - 1),
		13098 => to_unsigned(31154, LUT_AMPL_WIDTH - 1),
		13099 => to_unsigned(31155, LUT_AMPL_WIDTH - 1),
		13100 => to_unsigned(31156, LUT_AMPL_WIDTH - 1),
		13101 => to_unsigned(31157, LUT_AMPL_WIDTH - 1),
		13102 => to_unsigned(31158, LUT_AMPL_WIDTH - 1),
		13103 => to_unsigned(31159, LUT_AMPL_WIDTH - 1),
		13104 => to_unsigned(31160, LUT_AMPL_WIDTH - 1),
		13105 => to_unsigned(31161, LUT_AMPL_WIDTH - 1),
		13106 => to_unsigned(31162, LUT_AMPL_WIDTH - 1),
		13107 => to_unsigned(31163, LUT_AMPL_WIDTH - 1),
		13108 => to_unsigned(31164, LUT_AMPL_WIDTH - 1),
		13109 => to_unsigned(31165, LUT_AMPL_WIDTH - 1),
		13110 => to_unsigned(31166, LUT_AMPL_WIDTH - 1),
		13111 => to_unsigned(31167, LUT_AMPL_WIDTH - 1),
		13112 => to_unsigned(31168, LUT_AMPL_WIDTH - 1),
		13113 => to_unsigned(31169, LUT_AMPL_WIDTH - 1),
		13114 => to_unsigned(31170, LUT_AMPL_WIDTH - 1),
		13115 => to_unsigned(31171, LUT_AMPL_WIDTH - 1),
		13116 => to_unsigned(31172, LUT_AMPL_WIDTH - 1),
		13117 => to_unsigned(31173, LUT_AMPL_WIDTH - 1),
		13118 => to_unsigned(31174, LUT_AMPL_WIDTH - 1),
		13119 => to_unsigned(31175, LUT_AMPL_WIDTH - 1),
		13120 => to_unsigned(31176, LUT_AMPL_WIDTH - 1),
		13121 => to_unsigned(31177, LUT_AMPL_WIDTH - 1),
		13122 => to_unsigned(31178, LUT_AMPL_WIDTH - 1),
		13123 => to_unsigned(31179, LUT_AMPL_WIDTH - 1),
		13124 => to_unsigned(31180, LUT_AMPL_WIDTH - 1),
		13125 => to_unsigned(31181, LUT_AMPL_WIDTH - 1),
		13126 => to_unsigned(31181, LUT_AMPL_WIDTH - 1),
		13127 => to_unsigned(31182, LUT_AMPL_WIDTH - 1),
		13128 => to_unsigned(31183, LUT_AMPL_WIDTH - 1),
		13129 => to_unsigned(31184, LUT_AMPL_WIDTH - 1),
		13130 => to_unsigned(31185, LUT_AMPL_WIDTH - 1),
		13131 => to_unsigned(31186, LUT_AMPL_WIDTH - 1),
		13132 => to_unsigned(31187, LUT_AMPL_WIDTH - 1),
		13133 => to_unsigned(31188, LUT_AMPL_WIDTH - 1),
		13134 => to_unsigned(31189, LUT_AMPL_WIDTH - 1),
		13135 => to_unsigned(31190, LUT_AMPL_WIDTH - 1),
		13136 => to_unsigned(31191, LUT_AMPL_WIDTH - 1),
		13137 => to_unsigned(31192, LUT_AMPL_WIDTH - 1),
		13138 => to_unsigned(31193, LUT_AMPL_WIDTH - 1),
		13139 => to_unsigned(31194, LUT_AMPL_WIDTH - 1),
		13140 => to_unsigned(31195, LUT_AMPL_WIDTH - 1),
		13141 => to_unsigned(31196, LUT_AMPL_WIDTH - 1),
		13142 => to_unsigned(31197, LUT_AMPL_WIDTH - 1),
		13143 => to_unsigned(31198, LUT_AMPL_WIDTH - 1),
		13144 => to_unsigned(31199, LUT_AMPL_WIDTH - 1),
		13145 => to_unsigned(31200, LUT_AMPL_WIDTH - 1),
		13146 => to_unsigned(31201, LUT_AMPL_WIDTH - 1),
		13147 => to_unsigned(31202, LUT_AMPL_WIDTH - 1),
		13148 => to_unsigned(31203, LUT_AMPL_WIDTH - 1),
		13149 => to_unsigned(31204, LUT_AMPL_WIDTH - 1),
		13150 => to_unsigned(31205, LUT_AMPL_WIDTH - 1),
		13151 => to_unsigned(31206, LUT_AMPL_WIDTH - 1),
		13152 => to_unsigned(31206, LUT_AMPL_WIDTH - 1),
		13153 => to_unsigned(31207, LUT_AMPL_WIDTH - 1),
		13154 => to_unsigned(31208, LUT_AMPL_WIDTH - 1),
		13155 => to_unsigned(31209, LUT_AMPL_WIDTH - 1),
		13156 => to_unsigned(31210, LUT_AMPL_WIDTH - 1),
		13157 => to_unsigned(31211, LUT_AMPL_WIDTH - 1),
		13158 => to_unsigned(31212, LUT_AMPL_WIDTH - 1),
		13159 => to_unsigned(31213, LUT_AMPL_WIDTH - 1),
		13160 => to_unsigned(31214, LUT_AMPL_WIDTH - 1),
		13161 => to_unsigned(31215, LUT_AMPL_WIDTH - 1),
		13162 => to_unsigned(31216, LUT_AMPL_WIDTH - 1),
		13163 => to_unsigned(31217, LUT_AMPL_WIDTH - 1),
		13164 => to_unsigned(31218, LUT_AMPL_WIDTH - 1),
		13165 => to_unsigned(31219, LUT_AMPL_WIDTH - 1),
		13166 => to_unsigned(31220, LUT_AMPL_WIDTH - 1),
		13167 => to_unsigned(31221, LUT_AMPL_WIDTH - 1),
		13168 => to_unsigned(31222, LUT_AMPL_WIDTH - 1),
		13169 => to_unsigned(31223, LUT_AMPL_WIDTH - 1),
		13170 => to_unsigned(31224, LUT_AMPL_WIDTH - 1),
		13171 => to_unsigned(31225, LUT_AMPL_WIDTH - 1),
		13172 => to_unsigned(31226, LUT_AMPL_WIDTH - 1),
		13173 => to_unsigned(31227, LUT_AMPL_WIDTH - 1),
		13174 => to_unsigned(31227, LUT_AMPL_WIDTH - 1),
		13175 => to_unsigned(31228, LUT_AMPL_WIDTH - 1),
		13176 => to_unsigned(31229, LUT_AMPL_WIDTH - 1),
		13177 => to_unsigned(31230, LUT_AMPL_WIDTH - 1),
		13178 => to_unsigned(31231, LUT_AMPL_WIDTH - 1),
		13179 => to_unsigned(31232, LUT_AMPL_WIDTH - 1),
		13180 => to_unsigned(31233, LUT_AMPL_WIDTH - 1),
		13181 => to_unsigned(31234, LUT_AMPL_WIDTH - 1),
		13182 => to_unsigned(31235, LUT_AMPL_WIDTH - 1),
		13183 => to_unsigned(31236, LUT_AMPL_WIDTH - 1),
		13184 => to_unsigned(31237, LUT_AMPL_WIDTH - 1),
		13185 => to_unsigned(31238, LUT_AMPL_WIDTH - 1),
		13186 => to_unsigned(31239, LUT_AMPL_WIDTH - 1),
		13187 => to_unsigned(31240, LUT_AMPL_WIDTH - 1),
		13188 => to_unsigned(31241, LUT_AMPL_WIDTH - 1),
		13189 => to_unsigned(31242, LUT_AMPL_WIDTH - 1),
		13190 => to_unsigned(31243, LUT_AMPL_WIDTH - 1),
		13191 => to_unsigned(31244, LUT_AMPL_WIDTH - 1),
		13192 => to_unsigned(31245, LUT_AMPL_WIDTH - 1),
		13193 => to_unsigned(31246, LUT_AMPL_WIDTH - 1),
		13194 => to_unsigned(31246, LUT_AMPL_WIDTH - 1),
		13195 => to_unsigned(31247, LUT_AMPL_WIDTH - 1),
		13196 => to_unsigned(31248, LUT_AMPL_WIDTH - 1),
		13197 => to_unsigned(31249, LUT_AMPL_WIDTH - 1),
		13198 => to_unsigned(31250, LUT_AMPL_WIDTH - 1),
		13199 => to_unsigned(31251, LUT_AMPL_WIDTH - 1),
		13200 => to_unsigned(31252, LUT_AMPL_WIDTH - 1),
		13201 => to_unsigned(31253, LUT_AMPL_WIDTH - 1),
		13202 => to_unsigned(31254, LUT_AMPL_WIDTH - 1),
		13203 => to_unsigned(31255, LUT_AMPL_WIDTH - 1),
		13204 => to_unsigned(31256, LUT_AMPL_WIDTH - 1),
		13205 => to_unsigned(31257, LUT_AMPL_WIDTH - 1),
		13206 => to_unsigned(31258, LUT_AMPL_WIDTH - 1),
		13207 => to_unsigned(31259, LUT_AMPL_WIDTH - 1),
		13208 => to_unsigned(31260, LUT_AMPL_WIDTH - 1),
		13209 => to_unsigned(31261, LUT_AMPL_WIDTH - 1),
		13210 => to_unsigned(31262, LUT_AMPL_WIDTH - 1),
		13211 => to_unsigned(31262, LUT_AMPL_WIDTH - 1),
		13212 => to_unsigned(31263, LUT_AMPL_WIDTH - 1),
		13213 => to_unsigned(31264, LUT_AMPL_WIDTH - 1),
		13214 => to_unsigned(31265, LUT_AMPL_WIDTH - 1),
		13215 => to_unsigned(31266, LUT_AMPL_WIDTH - 1),
		13216 => to_unsigned(31267, LUT_AMPL_WIDTH - 1),
		13217 => to_unsigned(31268, LUT_AMPL_WIDTH - 1),
		13218 => to_unsigned(31269, LUT_AMPL_WIDTH - 1),
		13219 => to_unsigned(31270, LUT_AMPL_WIDTH - 1),
		13220 => to_unsigned(31271, LUT_AMPL_WIDTH - 1),
		13221 => to_unsigned(31272, LUT_AMPL_WIDTH - 1),
		13222 => to_unsigned(31273, LUT_AMPL_WIDTH - 1),
		13223 => to_unsigned(31274, LUT_AMPL_WIDTH - 1),
		13224 => to_unsigned(31275, LUT_AMPL_WIDTH - 1),
		13225 => to_unsigned(31276, LUT_AMPL_WIDTH - 1),
		13226 => to_unsigned(31277, LUT_AMPL_WIDTH - 1),
		13227 => to_unsigned(31278, LUT_AMPL_WIDTH - 1),
		13228 => to_unsigned(31278, LUT_AMPL_WIDTH - 1),
		13229 => to_unsigned(31279, LUT_AMPL_WIDTH - 1),
		13230 => to_unsigned(31280, LUT_AMPL_WIDTH - 1),
		13231 => to_unsigned(31281, LUT_AMPL_WIDTH - 1),
		13232 => to_unsigned(31282, LUT_AMPL_WIDTH - 1),
		13233 => to_unsigned(31283, LUT_AMPL_WIDTH - 1),
		13234 => to_unsigned(31284, LUT_AMPL_WIDTH - 1),
		13235 => to_unsigned(31285, LUT_AMPL_WIDTH - 1),
		13236 => to_unsigned(31286, LUT_AMPL_WIDTH - 1),
		13237 => to_unsigned(31287, LUT_AMPL_WIDTH - 1),
		13238 => to_unsigned(31288, LUT_AMPL_WIDTH - 1),
		13239 => to_unsigned(31289, LUT_AMPL_WIDTH - 1),
		13240 => to_unsigned(31290, LUT_AMPL_WIDTH - 1),
		13241 => to_unsigned(31291, LUT_AMPL_WIDTH - 1),
		13242 => to_unsigned(31292, LUT_AMPL_WIDTH - 1),
		13243 => to_unsigned(31292, LUT_AMPL_WIDTH - 1),
		13244 => to_unsigned(31293, LUT_AMPL_WIDTH - 1),
		13245 => to_unsigned(31294, LUT_AMPL_WIDTH - 1),
		13246 => to_unsigned(31295, LUT_AMPL_WIDTH - 1),
		13247 => to_unsigned(31296, LUT_AMPL_WIDTH - 1),
		13248 => to_unsigned(31297, LUT_AMPL_WIDTH - 1),
		13249 => to_unsigned(31298, LUT_AMPL_WIDTH - 1),
		13250 => to_unsigned(31299, LUT_AMPL_WIDTH - 1),
		13251 => to_unsigned(31300, LUT_AMPL_WIDTH - 1),
		13252 => to_unsigned(31301, LUT_AMPL_WIDTH - 1),
		13253 => to_unsigned(31302, LUT_AMPL_WIDTH - 1),
		13254 => to_unsigned(31303, LUT_AMPL_WIDTH - 1),
		13255 => to_unsigned(31304, LUT_AMPL_WIDTH - 1),
		13256 => to_unsigned(31305, LUT_AMPL_WIDTH - 1),
		13257 => to_unsigned(31305, LUT_AMPL_WIDTH - 1),
		13258 => to_unsigned(31306, LUT_AMPL_WIDTH - 1),
		13259 => to_unsigned(31307, LUT_AMPL_WIDTH - 1),
		13260 => to_unsigned(31308, LUT_AMPL_WIDTH - 1),
		13261 => to_unsigned(31309, LUT_AMPL_WIDTH - 1),
		13262 => to_unsigned(31310, LUT_AMPL_WIDTH - 1),
		13263 => to_unsigned(31311, LUT_AMPL_WIDTH - 1),
		13264 => to_unsigned(31312, LUT_AMPL_WIDTH - 1),
		13265 => to_unsigned(31313, LUT_AMPL_WIDTH - 1),
		13266 => to_unsigned(31314, LUT_AMPL_WIDTH - 1),
		13267 => to_unsigned(31315, LUT_AMPL_WIDTH - 1),
		13268 => to_unsigned(31316, LUT_AMPL_WIDTH - 1),
		13269 => to_unsigned(31317, LUT_AMPL_WIDTH - 1),
		13270 => to_unsigned(31318, LUT_AMPL_WIDTH - 1),
		13271 => to_unsigned(31318, LUT_AMPL_WIDTH - 1),
		13272 => to_unsigned(31319, LUT_AMPL_WIDTH - 1),
		13273 => to_unsigned(31320, LUT_AMPL_WIDTH - 1),
		13274 => to_unsigned(31321, LUT_AMPL_WIDTH - 1),
		13275 => to_unsigned(31322, LUT_AMPL_WIDTH - 1),
		13276 => to_unsigned(31323, LUT_AMPL_WIDTH - 1),
		13277 => to_unsigned(31324, LUT_AMPL_WIDTH - 1),
		13278 => to_unsigned(31325, LUT_AMPL_WIDTH - 1),
		13279 => to_unsigned(31326, LUT_AMPL_WIDTH - 1),
		13280 => to_unsigned(31327, LUT_AMPL_WIDTH - 1),
		13281 => to_unsigned(31328, LUT_AMPL_WIDTH - 1),
		13282 => to_unsigned(31329, LUT_AMPL_WIDTH - 1),
		13283 => to_unsigned(31329, LUT_AMPL_WIDTH - 1),
		13284 => to_unsigned(31330, LUT_AMPL_WIDTH - 1),
		13285 => to_unsigned(31331, LUT_AMPL_WIDTH - 1),
		13286 => to_unsigned(31332, LUT_AMPL_WIDTH - 1),
		13287 => to_unsigned(31333, LUT_AMPL_WIDTH - 1),
		13288 => to_unsigned(31334, LUT_AMPL_WIDTH - 1),
		13289 => to_unsigned(31335, LUT_AMPL_WIDTH - 1),
		13290 => to_unsigned(31336, LUT_AMPL_WIDTH - 1),
		13291 => to_unsigned(31337, LUT_AMPL_WIDTH - 1),
		13292 => to_unsigned(31338, LUT_AMPL_WIDTH - 1),
		13293 => to_unsigned(31339, LUT_AMPL_WIDTH - 1),
		13294 => to_unsigned(31340, LUT_AMPL_WIDTH - 1),
		13295 => to_unsigned(31341, LUT_AMPL_WIDTH - 1),
		13296 => to_unsigned(31341, LUT_AMPL_WIDTH - 1),
		13297 => to_unsigned(31342, LUT_AMPL_WIDTH - 1),
		13298 => to_unsigned(31343, LUT_AMPL_WIDTH - 1),
		13299 => to_unsigned(31344, LUT_AMPL_WIDTH - 1),
		13300 => to_unsigned(31345, LUT_AMPL_WIDTH - 1),
		13301 => to_unsigned(31346, LUT_AMPL_WIDTH - 1),
		13302 => to_unsigned(31347, LUT_AMPL_WIDTH - 1),
		13303 => to_unsigned(31348, LUT_AMPL_WIDTH - 1),
		13304 => to_unsigned(31349, LUT_AMPL_WIDTH - 1),
		13305 => to_unsigned(31350, LUT_AMPL_WIDTH - 1),
		13306 => to_unsigned(31351, LUT_AMPL_WIDTH - 1),
		13307 => to_unsigned(31352, LUT_AMPL_WIDTH - 1),
		13308 => to_unsigned(31352, LUT_AMPL_WIDTH - 1),
		13309 => to_unsigned(31353, LUT_AMPL_WIDTH - 1),
		13310 => to_unsigned(31354, LUT_AMPL_WIDTH - 1),
		13311 => to_unsigned(31355, LUT_AMPL_WIDTH - 1),
		13312 => to_unsigned(31356, LUT_AMPL_WIDTH - 1),
		13313 => to_unsigned(31357, LUT_AMPL_WIDTH - 1),
		13314 => to_unsigned(31358, LUT_AMPL_WIDTH - 1),
		13315 => to_unsigned(31359, LUT_AMPL_WIDTH - 1),
		13316 => to_unsigned(31360, LUT_AMPL_WIDTH - 1),
		13317 => to_unsigned(31361, LUT_AMPL_WIDTH - 1),
		13318 => to_unsigned(31362, LUT_AMPL_WIDTH - 1),
		13319 => to_unsigned(31362, LUT_AMPL_WIDTH - 1),
		13320 => to_unsigned(31363, LUT_AMPL_WIDTH - 1),
		13321 => to_unsigned(31364, LUT_AMPL_WIDTH - 1),
		13322 => to_unsigned(31365, LUT_AMPL_WIDTH - 1),
		13323 => to_unsigned(31366, LUT_AMPL_WIDTH - 1),
		13324 => to_unsigned(31367, LUT_AMPL_WIDTH - 1),
		13325 => to_unsigned(31368, LUT_AMPL_WIDTH - 1),
		13326 => to_unsigned(31369, LUT_AMPL_WIDTH - 1),
		13327 => to_unsigned(31370, LUT_AMPL_WIDTH - 1),
		13328 => to_unsigned(31371, LUT_AMPL_WIDTH - 1),
		13329 => to_unsigned(31372, LUT_AMPL_WIDTH - 1),
		13330 => to_unsigned(31372, LUT_AMPL_WIDTH - 1),
		13331 => to_unsigned(31373, LUT_AMPL_WIDTH - 1),
		13332 => to_unsigned(31374, LUT_AMPL_WIDTH - 1),
		13333 => to_unsigned(31375, LUT_AMPL_WIDTH - 1),
		13334 => to_unsigned(31376, LUT_AMPL_WIDTH - 1),
		13335 => to_unsigned(31377, LUT_AMPL_WIDTH - 1),
		13336 => to_unsigned(31378, LUT_AMPL_WIDTH - 1),
		13337 => to_unsigned(31379, LUT_AMPL_WIDTH - 1),
		13338 => to_unsigned(31380, LUT_AMPL_WIDTH - 1),
		13339 => to_unsigned(31381, LUT_AMPL_WIDTH - 1),
		13340 => to_unsigned(31381, LUT_AMPL_WIDTH - 1),
		13341 => to_unsigned(31382, LUT_AMPL_WIDTH - 1),
		13342 => to_unsigned(31383, LUT_AMPL_WIDTH - 1),
		13343 => to_unsigned(31384, LUT_AMPL_WIDTH - 1),
		13344 => to_unsigned(31385, LUT_AMPL_WIDTH - 1),
		13345 => to_unsigned(31386, LUT_AMPL_WIDTH - 1),
		13346 => to_unsigned(31387, LUT_AMPL_WIDTH - 1),
		13347 => to_unsigned(31388, LUT_AMPL_WIDTH - 1),
		13348 => to_unsigned(31389, LUT_AMPL_WIDTH - 1),
		13349 => to_unsigned(31390, LUT_AMPL_WIDTH - 1),
		13350 => to_unsigned(31391, LUT_AMPL_WIDTH - 1),
		13351 => to_unsigned(31391, LUT_AMPL_WIDTH - 1),
		13352 => to_unsigned(31392, LUT_AMPL_WIDTH - 1),
		13353 => to_unsigned(31393, LUT_AMPL_WIDTH - 1),
		13354 => to_unsigned(31394, LUT_AMPL_WIDTH - 1),
		13355 => to_unsigned(31395, LUT_AMPL_WIDTH - 1),
		13356 => to_unsigned(31396, LUT_AMPL_WIDTH - 1),
		13357 => to_unsigned(31397, LUT_AMPL_WIDTH - 1),
		13358 => to_unsigned(31398, LUT_AMPL_WIDTH - 1),
		13359 => to_unsigned(31399, LUT_AMPL_WIDTH - 1),
		13360 => to_unsigned(31400, LUT_AMPL_WIDTH - 1),
		13361 => to_unsigned(31400, LUT_AMPL_WIDTH - 1),
		13362 => to_unsigned(31401, LUT_AMPL_WIDTH - 1),
		13363 => to_unsigned(31402, LUT_AMPL_WIDTH - 1),
		13364 => to_unsigned(31403, LUT_AMPL_WIDTH - 1),
		13365 => to_unsigned(31404, LUT_AMPL_WIDTH - 1),
		13366 => to_unsigned(31405, LUT_AMPL_WIDTH - 1),
		13367 => to_unsigned(31406, LUT_AMPL_WIDTH - 1),
		13368 => to_unsigned(31407, LUT_AMPL_WIDTH - 1),
		13369 => to_unsigned(31408, LUT_AMPL_WIDTH - 1),
		13370 => to_unsigned(31408, LUT_AMPL_WIDTH - 1),
		13371 => to_unsigned(31409, LUT_AMPL_WIDTH - 1),
		13372 => to_unsigned(31410, LUT_AMPL_WIDTH - 1),
		13373 => to_unsigned(31411, LUT_AMPL_WIDTH - 1),
		13374 => to_unsigned(31412, LUT_AMPL_WIDTH - 1),
		13375 => to_unsigned(31413, LUT_AMPL_WIDTH - 1),
		13376 => to_unsigned(31414, LUT_AMPL_WIDTH - 1),
		13377 => to_unsigned(31415, LUT_AMPL_WIDTH - 1),
		13378 => to_unsigned(31416, LUT_AMPL_WIDTH - 1),
		13379 => to_unsigned(31417, LUT_AMPL_WIDTH - 1),
		13380 => to_unsigned(31417, LUT_AMPL_WIDTH - 1),
		13381 => to_unsigned(31418, LUT_AMPL_WIDTH - 1),
		13382 => to_unsigned(31419, LUT_AMPL_WIDTH - 1),
		13383 => to_unsigned(31420, LUT_AMPL_WIDTH - 1),
		13384 => to_unsigned(31421, LUT_AMPL_WIDTH - 1),
		13385 => to_unsigned(31422, LUT_AMPL_WIDTH - 1),
		13386 => to_unsigned(31423, LUT_AMPL_WIDTH - 1),
		13387 => to_unsigned(31424, LUT_AMPL_WIDTH - 1),
		13388 => to_unsigned(31425, LUT_AMPL_WIDTH - 1),
		13389 => to_unsigned(31425, LUT_AMPL_WIDTH - 1),
		13390 => to_unsigned(31426, LUT_AMPL_WIDTH - 1),
		13391 => to_unsigned(31427, LUT_AMPL_WIDTH - 1),
		13392 => to_unsigned(31428, LUT_AMPL_WIDTH - 1),
		13393 => to_unsigned(31429, LUT_AMPL_WIDTH - 1),
		13394 => to_unsigned(31430, LUT_AMPL_WIDTH - 1),
		13395 => to_unsigned(31431, LUT_AMPL_WIDTH - 1),
		13396 => to_unsigned(31432, LUT_AMPL_WIDTH - 1),
		13397 => to_unsigned(31433, LUT_AMPL_WIDTH - 1),
		13398 => to_unsigned(31433, LUT_AMPL_WIDTH - 1),
		13399 => to_unsigned(31434, LUT_AMPL_WIDTH - 1),
		13400 => to_unsigned(31435, LUT_AMPL_WIDTH - 1),
		13401 => to_unsigned(31436, LUT_AMPL_WIDTH - 1),
		13402 => to_unsigned(31437, LUT_AMPL_WIDTH - 1),
		13403 => to_unsigned(31438, LUT_AMPL_WIDTH - 1),
		13404 => to_unsigned(31439, LUT_AMPL_WIDTH - 1),
		13405 => to_unsigned(31440, LUT_AMPL_WIDTH - 1),
		13406 => to_unsigned(31441, LUT_AMPL_WIDTH - 1),
		13407 => to_unsigned(31441, LUT_AMPL_WIDTH - 1),
		13408 => to_unsigned(31442, LUT_AMPL_WIDTH - 1),
		13409 => to_unsigned(31443, LUT_AMPL_WIDTH - 1),
		13410 => to_unsigned(31444, LUT_AMPL_WIDTH - 1),
		13411 => to_unsigned(31445, LUT_AMPL_WIDTH - 1),
		13412 => to_unsigned(31446, LUT_AMPL_WIDTH - 1),
		13413 => to_unsigned(31447, LUT_AMPL_WIDTH - 1),
		13414 => to_unsigned(31448, LUT_AMPL_WIDTH - 1),
		13415 => to_unsigned(31448, LUT_AMPL_WIDTH - 1),
		13416 => to_unsigned(31449, LUT_AMPL_WIDTH - 1),
		13417 => to_unsigned(31450, LUT_AMPL_WIDTH - 1),
		13418 => to_unsigned(31451, LUT_AMPL_WIDTH - 1),
		13419 => to_unsigned(31452, LUT_AMPL_WIDTH - 1),
		13420 => to_unsigned(31453, LUT_AMPL_WIDTH - 1),
		13421 => to_unsigned(31454, LUT_AMPL_WIDTH - 1),
		13422 => to_unsigned(31455, LUT_AMPL_WIDTH - 1),
		13423 => to_unsigned(31456, LUT_AMPL_WIDTH - 1),
		13424 => to_unsigned(31456, LUT_AMPL_WIDTH - 1),
		13425 => to_unsigned(31457, LUT_AMPL_WIDTH - 1),
		13426 => to_unsigned(31458, LUT_AMPL_WIDTH - 1),
		13427 => to_unsigned(31459, LUT_AMPL_WIDTH - 1),
		13428 => to_unsigned(31460, LUT_AMPL_WIDTH - 1),
		13429 => to_unsigned(31461, LUT_AMPL_WIDTH - 1),
		13430 => to_unsigned(31462, LUT_AMPL_WIDTH - 1),
		13431 => to_unsigned(31463, LUT_AMPL_WIDTH - 1),
		13432 => to_unsigned(31463, LUT_AMPL_WIDTH - 1),
		13433 => to_unsigned(31464, LUT_AMPL_WIDTH - 1),
		13434 => to_unsigned(31465, LUT_AMPL_WIDTH - 1),
		13435 => to_unsigned(31466, LUT_AMPL_WIDTH - 1),
		13436 => to_unsigned(31467, LUT_AMPL_WIDTH - 1),
		13437 => to_unsigned(31468, LUT_AMPL_WIDTH - 1),
		13438 => to_unsigned(31469, LUT_AMPL_WIDTH - 1),
		13439 => to_unsigned(31470, LUT_AMPL_WIDTH - 1),
		13440 => to_unsigned(31470, LUT_AMPL_WIDTH - 1),
		13441 => to_unsigned(31471, LUT_AMPL_WIDTH - 1),
		13442 => to_unsigned(31472, LUT_AMPL_WIDTH - 1),
		13443 => to_unsigned(31473, LUT_AMPL_WIDTH - 1),
		13444 => to_unsigned(31474, LUT_AMPL_WIDTH - 1),
		13445 => to_unsigned(31475, LUT_AMPL_WIDTH - 1),
		13446 => to_unsigned(31476, LUT_AMPL_WIDTH - 1),
		13447 => to_unsigned(31477, LUT_AMPL_WIDTH - 1),
		13448 => to_unsigned(31477, LUT_AMPL_WIDTH - 1),
		13449 => to_unsigned(31478, LUT_AMPL_WIDTH - 1),
		13450 => to_unsigned(31479, LUT_AMPL_WIDTH - 1),
		13451 => to_unsigned(31480, LUT_AMPL_WIDTH - 1),
		13452 => to_unsigned(31481, LUT_AMPL_WIDTH - 1),
		13453 => to_unsigned(31482, LUT_AMPL_WIDTH - 1),
		13454 => to_unsigned(31483, LUT_AMPL_WIDTH - 1),
		13455 => to_unsigned(31484, LUT_AMPL_WIDTH - 1),
		13456 => to_unsigned(31484, LUT_AMPL_WIDTH - 1),
		13457 => to_unsigned(31485, LUT_AMPL_WIDTH - 1),
		13458 => to_unsigned(31486, LUT_AMPL_WIDTH - 1),
		13459 => to_unsigned(31487, LUT_AMPL_WIDTH - 1),
		13460 => to_unsigned(31488, LUT_AMPL_WIDTH - 1),
		13461 => to_unsigned(31489, LUT_AMPL_WIDTH - 1),
		13462 => to_unsigned(31490, LUT_AMPL_WIDTH - 1),
		13463 => to_unsigned(31490, LUT_AMPL_WIDTH - 1),
		13464 => to_unsigned(31491, LUT_AMPL_WIDTH - 1),
		13465 => to_unsigned(31492, LUT_AMPL_WIDTH - 1),
		13466 => to_unsigned(31493, LUT_AMPL_WIDTH - 1),
		13467 => to_unsigned(31494, LUT_AMPL_WIDTH - 1),
		13468 => to_unsigned(31495, LUT_AMPL_WIDTH - 1),
		13469 => to_unsigned(31496, LUT_AMPL_WIDTH - 1),
		13470 => to_unsigned(31497, LUT_AMPL_WIDTH - 1),
		13471 => to_unsigned(31497, LUT_AMPL_WIDTH - 1),
		13472 => to_unsigned(31498, LUT_AMPL_WIDTH - 1),
		13473 => to_unsigned(31499, LUT_AMPL_WIDTH - 1),
		13474 => to_unsigned(31500, LUT_AMPL_WIDTH - 1),
		13475 => to_unsigned(31501, LUT_AMPL_WIDTH - 1),
		13476 => to_unsigned(31502, LUT_AMPL_WIDTH - 1),
		13477 => to_unsigned(31503, LUT_AMPL_WIDTH - 1),
		13478 => to_unsigned(31503, LUT_AMPL_WIDTH - 1),
		13479 => to_unsigned(31504, LUT_AMPL_WIDTH - 1),
		13480 => to_unsigned(31505, LUT_AMPL_WIDTH - 1),
		13481 => to_unsigned(31506, LUT_AMPL_WIDTH - 1),
		13482 => to_unsigned(31507, LUT_AMPL_WIDTH - 1),
		13483 => to_unsigned(31508, LUT_AMPL_WIDTH - 1),
		13484 => to_unsigned(31509, LUT_AMPL_WIDTH - 1),
		13485 => to_unsigned(31510, LUT_AMPL_WIDTH - 1),
		13486 => to_unsigned(31510, LUT_AMPL_WIDTH - 1),
		13487 => to_unsigned(31511, LUT_AMPL_WIDTH - 1),
		13488 => to_unsigned(31512, LUT_AMPL_WIDTH - 1),
		13489 => to_unsigned(31513, LUT_AMPL_WIDTH - 1),
		13490 => to_unsigned(31514, LUT_AMPL_WIDTH - 1),
		13491 => to_unsigned(31515, LUT_AMPL_WIDTH - 1),
		13492 => to_unsigned(31516, LUT_AMPL_WIDTH - 1),
		13493 => to_unsigned(31516, LUT_AMPL_WIDTH - 1),
		13494 => to_unsigned(31517, LUT_AMPL_WIDTH - 1),
		13495 => to_unsigned(31518, LUT_AMPL_WIDTH - 1),
		13496 => to_unsigned(31519, LUT_AMPL_WIDTH - 1),
		13497 => to_unsigned(31520, LUT_AMPL_WIDTH - 1),
		13498 => to_unsigned(31521, LUT_AMPL_WIDTH - 1),
		13499 => to_unsigned(31522, LUT_AMPL_WIDTH - 1),
		13500 => to_unsigned(31522, LUT_AMPL_WIDTH - 1),
		13501 => to_unsigned(31523, LUT_AMPL_WIDTH - 1),
		13502 => to_unsigned(31524, LUT_AMPL_WIDTH - 1),
		13503 => to_unsigned(31525, LUT_AMPL_WIDTH - 1),
		13504 => to_unsigned(31526, LUT_AMPL_WIDTH - 1),
		13505 => to_unsigned(31527, LUT_AMPL_WIDTH - 1),
		13506 => to_unsigned(31528, LUT_AMPL_WIDTH - 1),
		13507 => to_unsigned(31528, LUT_AMPL_WIDTH - 1),
		13508 => to_unsigned(31529, LUT_AMPL_WIDTH - 1),
		13509 => to_unsigned(31530, LUT_AMPL_WIDTH - 1),
		13510 => to_unsigned(31531, LUT_AMPL_WIDTH - 1),
		13511 => to_unsigned(31532, LUT_AMPL_WIDTH - 1),
		13512 => to_unsigned(31533, LUT_AMPL_WIDTH - 1),
		13513 => to_unsigned(31534, LUT_AMPL_WIDTH - 1),
		13514 => to_unsigned(31534, LUT_AMPL_WIDTH - 1),
		13515 => to_unsigned(31535, LUT_AMPL_WIDTH - 1),
		13516 => to_unsigned(31536, LUT_AMPL_WIDTH - 1),
		13517 => to_unsigned(31537, LUT_AMPL_WIDTH - 1),
		13518 => to_unsigned(31538, LUT_AMPL_WIDTH - 1),
		13519 => to_unsigned(31539, LUT_AMPL_WIDTH - 1),
		13520 => to_unsigned(31539, LUT_AMPL_WIDTH - 1),
		13521 => to_unsigned(31540, LUT_AMPL_WIDTH - 1),
		13522 => to_unsigned(31541, LUT_AMPL_WIDTH - 1),
		13523 => to_unsigned(31542, LUT_AMPL_WIDTH - 1),
		13524 => to_unsigned(31543, LUT_AMPL_WIDTH - 1),
		13525 => to_unsigned(31544, LUT_AMPL_WIDTH - 1),
		13526 => to_unsigned(31545, LUT_AMPL_WIDTH - 1),
		13527 => to_unsigned(31545, LUT_AMPL_WIDTH - 1),
		13528 => to_unsigned(31546, LUT_AMPL_WIDTH - 1),
		13529 => to_unsigned(31547, LUT_AMPL_WIDTH - 1),
		13530 => to_unsigned(31548, LUT_AMPL_WIDTH - 1),
		13531 => to_unsigned(31549, LUT_AMPL_WIDTH - 1),
		13532 => to_unsigned(31550, LUT_AMPL_WIDTH - 1),
		13533 => to_unsigned(31551, LUT_AMPL_WIDTH - 1),
		13534 => to_unsigned(31551, LUT_AMPL_WIDTH - 1),
		13535 => to_unsigned(31552, LUT_AMPL_WIDTH - 1),
		13536 => to_unsigned(31553, LUT_AMPL_WIDTH - 1),
		13537 => to_unsigned(31554, LUT_AMPL_WIDTH - 1),
		13538 => to_unsigned(31555, LUT_AMPL_WIDTH - 1),
		13539 => to_unsigned(31556, LUT_AMPL_WIDTH - 1),
		13540 => to_unsigned(31556, LUT_AMPL_WIDTH - 1),
		13541 => to_unsigned(31557, LUT_AMPL_WIDTH - 1),
		13542 => to_unsigned(31558, LUT_AMPL_WIDTH - 1),
		13543 => to_unsigned(31559, LUT_AMPL_WIDTH - 1),
		13544 => to_unsigned(31560, LUT_AMPL_WIDTH - 1),
		13545 => to_unsigned(31561, LUT_AMPL_WIDTH - 1),
		13546 => to_unsigned(31562, LUT_AMPL_WIDTH - 1),
		13547 => to_unsigned(31562, LUT_AMPL_WIDTH - 1),
		13548 => to_unsigned(31563, LUT_AMPL_WIDTH - 1),
		13549 => to_unsigned(31564, LUT_AMPL_WIDTH - 1),
		13550 => to_unsigned(31565, LUT_AMPL_WIDTH - 1),
		13551 => to_unsigned(31566, LUT_AMPL_WIDTH - 1),
		13552 => to_unsigned(31567, LUT_AMPL_WIDTH - 1),
		13553 => to_unsigned(31567, LUT_AMPL_WIDTH - 1),
		13554 => to_unsigned(31568, LUT_AMPL_WIDTH - 1),
		13555 => to_unsigned(31569, LUT_AMPL_WIDTH - 1),
		13556 => to_unsigned(31570, LUT_AMPL_WIDTH - 1),
		13557 => to_unsigned(31571, LUT_AMPL_WIDTH - 1),
		13558 => to_unsigned(31572, LUT_AMPL_WIDTH - 1),
		13559 => to_unsigned(31572, LUT_AMPL_WIDTH - 1),
		13560 => to_unsigned(31573, LUT_AMPL_WIDTH - 1),
		13561 => to_unsigned(31574, LUT_AMPL_WIDTH - 1),
		13562 => to_unsigned(31575, LUT_AMPL_WIDTH - 1),
		13563 => to_unsigned(31576, LUT_AMPL_WIDTH - 1),
		13564 => to_unsigned(31577, LUT_AMPL_WIDTH - 1),
		13565 => to_unsigned(31578, LUT_AMPL_WIDTH - 1),
		13566 => to_unsigned(31578, LUT_AMPL_WIDTH - 1),
		13567 => to_unsigned(31579, LUT_AMPL_WIDTH - 1),
		13568 => to_unsigned(31580, LUT_AMPL_WIDTH - 1),
		13569 => to_unsigned(31581, LUT_AMPL_WIDTH - 1),
		13570 => to_unsigned(31582, LUT_AMPL_WIDTH - 1),
		13571 => to_unsigned(31583, LUT_AMPL_WIDTH - 1),
		13572 => to_unsigned(31583, LUT_AMPL_WIDTH - 1),
		13573 => to_unsigned(31584, LUT_AMPL_WIDTH - 1),
		13574 => to_unsigned(31585, LUT_AMPL_WIDTH - 1),
		13575 => to_unsigned(31586, LUT_AMPL_WIDTH - 1),
		13576 => to_unsigned(31587, LUT_AMPL_WIDTH - 1),
		13577 => to_unsigned(31588, LUT_AMPL_WIDTH - 1),
		13578 => to_unsigned(31588, LUT_AMPL_WIDTH - 1),
		13579 => to_unsigned(31589, LUT_AMPL_WIDTH - 1),
		13580 => to_unsigned(31590, LUT_AMPL_WIDTH - 1),
		13581 => to_unsigned(31591, LUT_AMPL_WIDTH - 1),
		13582 => to_unsigned(31592, LUT_AMPL_WIDTH - 1),
		13583 => to_unsigned(31593, LUT_AMPL_WIDTH - 1),
		13584 => to_unsigned(31593, LUT_AMPL_WIDTH - 1),
		13585 => to_unsigned(31594, LUT_AMPL_WIDTH - 1),
		13586 => to_unsigned(31595, LUT_AMPL_WIDTH - 1),
		13587 => to_unsigned(31596, LUT_AMPL_WIDTH - 1),
		13588 => to_unsigned(31597, LUT_AMPL_WIDTH - 1),
		13589 => to_unsigned(31598, LUT_AMPL_WIDTH - 1),
		13590 => to_unsigned(31598, LUT_AMPL_WIDTH - 1),
		13591 => to_unsigned(31599, LUT_AMPL_WIDTH - 1),
		13592 => to_unsigned(31600, LUT_AMPL_WIDTH - 1),
		13593 => to_unsigned(31601, LUT_AMPL_WIDTH - 1),
		13594 => to_unsigned(31602, LUT_AMPL_WIDTH - 1),
		13595 => to_unsigned(31603, LUT_AMPL_WIDTH - 1),
		13596 => to_unsigned(31603, LUT_AMPL_WIDTH - 1),
		13597 => to_unsigned(31604, LUT_AMPL_WIDTH - 1),
		13598 => to_unsigned(31605, LUT_AMPL_WIDTH - 1),
		13599 => to_unsigned(31606, LUT_AMPL_WIDTH - 1),
		13600 => to_unsigned(31607, LUT_AMPL_WIDTH - 1),
		13601 => to_unsigned(31608, LUT_AMPL_WIDTH - 1),
		13602 => to_unsigned(31608, LUT_AMPL_WIDTH - 1),
		13603 => to_unsigned(31609, LUT_AMPL_WIDTH - 1),
		13604 => to_unsigned(31610, LUT_AMPL_WIDTH - 1),
		13605 => to_unsigned(31611, LUT_AMPL_WIDTH - 1),
		13606 => to_unsigned(31612, LUT_AMPL_WIDTH - 1),
		13607 => to_unsigned(31613, LUT_AMPL_WIDTH - 1),
		13608 => to_unsigned(31613, LUT_AMPL_WIDTH - 1),
		13609 => to_unsigned(31614, LUT_AMPL_WIDTH - 1),
		13610 => to_unsigned(31615, LUT_AMPL_WIDTH - 1),
		13611 => to_unsigned(31616, LUT_AMPL_WIDTH - 1),
		13612 => to_unsigned(31617, LUT_AMPL_WIDTH - 1),
		13613 => to_unsigned(31617, LUT_AMPL_WIDTH - 1),
		13614 => to_unsigned(31618, LUT_AMPL_WIDTH - 1),
		13615 => to_unsigned(31619, LUT_AMPL_WIDTH - 1),
		13616 => to_unsigned(31620, LUT_AMPL_WIDTH - 1),
		13617 => to_unsigned(31621, LUT_AMPL_WIDTH - 1),
		13618 => to_unsigned(31622, LUT_AMPL_WIDTH - 1),
		13619 => to_unsigned(31622, LUT_AMPL_WIDTH - 1),
		13620 => to_unsigned(31623, LUT_AMPL_WIDTH - 1),
		13621 => to_unsigned(31624, LUT_AMPL_WIDTH - 1),
		13622 => to_unsigned(31625, LUT_AMPL_WIDTH - 1),
		13623 => to_unsigned(31626, LUT_AMPL_WIDTH - 1),
		13624 => to_unsigned(31627, LUT_AMPL_WIDTH - 1),
		13625 => to_unsigned(31627, LUT_AMPL_WIDTH - 1),
		13626 => to_unsigned(31628, LUT_AMPL_WIDTH - 1),
		13627 => to_unsigned(31629, LUT_AMPL_WIDTH - 1),
		13628 => to_unsigned(31630, LUT_AMPL_WIDTH - 1),
		13629 => to_unsigned(31631, LUT_AMPL_WIDTH - 1),
		13630 => to_unsigned(31631, LUT_AMPL_WIDTH - 1),
		13631 => to_unsigned(31632, LUT_AMPL_WIDTH - 1),
		13632 => to_unsigned(31633, LUT_AMPL_WIDTH - 1),
		13633 => to_unsigned(31634, LUT_AMPL_WIDTH - 1),
		13634 => to_unsigned(31635, LUT_AMPL_WIDTH - 1),
		13635 => to_unsigned(31636, LUT_AMPL_WIDTH - 1),
		13636 => to_unsigned(31636, LUT_AMPL_WIDTH - 1),
		13637 => to_unsigned(31637, LUT_AMPL_WIDTH - 1),
		13638 => to_unsigned(31638, LUT_AMPL_WIDTH - 1),
		13639 => to_unsigned(31639, LUT_AMPL_WIDTH - 1),
		13640 => to_unsigned(31640, LUT_AMPL_WIDTH - 1),
		13641 => to_unsigned(31640, LUT_AMPL_WIDTH - 1),
		13642 => to_unsigned(31641, LUT_AMPL_WIDTH - 1),
		13643 => to_unsigned(31642, LUT_AMPL_WIDTH - 1),
		13644 => to_unsigned(31643, LUT_AMPL_WIDTH - 1),
		13645 => to_unsigned(31644, LUT_AMPL_WIDTH - 1),
		13646 => to_unsigned(31645, LUT_AMPL_WIDTH - 1),
		13647 => to_unsigned(31645, LUT_AMPL_WIDTH - 1),
		13648 => to_unsigned(31646, LUT_AMPL_WIDTH - 1),
		13649 => to_unsigned(31647, LUT_AMPL_WIDTH - 1),
		13650 => to_unsigned(31648, LUT_AMPL_WIDTH - 1),
		13651 => to_unsigned(31649, LUT_AMPL_WIDTH - 1),
		13652 => to_unsigned(31649, LUT_AMPL_WIDTH - 1),
		13653 => to_unsigned(31650, LUT_AMPL_WIDTH - 1),
		13654 => to_unsigned(31651, LUT_AMPL_WIDTH - 1),
		13655 => to_unsigned(31652, LUT_AMPL_WIDTH - 1),
		13656 => to_unsigned(31653, LUT_AMPL_WIDTH - 1),
		13657 => to_unsigned(31653, LUT_AMPL_WIDTH - 1),
		13658 => to_unsigned(31654, LUT_AMPL_WIDTH - 1),
		13659 => to_unsigned(31655, LUT_AMPL_WIDTH - 1),
		13660 => to_unsigned(31656, LUT_AMPL_WIDTH - 1),
		13661 => to_unsigned(31657, LUT_AMPL_WIDTH - 1),
		13662 => to_unsigned(31658, LUT_AMPL_WIDTH - 1),
		13663 => to_unsigned(31658, LUT_AMPL_WIDTH - 1),
		13664 => to_unsigned(31659, LUT_AMPL_WIDTH - 1),
		13665 => to_unsigned(31660, LUT_AMPL_WIDTH - 1),
		13666 => to_unsigned(31661, LUT_AMPL_WIDTH - 1),
		13667 => to_unsigned(31662, LUT_AMPL_WIDTH - 1),
		13668 => to_unsigned(31662, LUT_AMPL_WIDTH - 1),
		13669 => to_unsigned(31663, LUT_AMPL_WIDTH - 1),
		13670 => to_unsigned(31664, LUT_AMPL_WIDTH - 1),
		13671 => to_unsigned(31665, LUT_AMPL_WIDTH - 1),
		13672 => to_unsigned(31666, LUT_AMPL_WIDTH - 1),
		13673 => to_unsigned(31666, LUT_AMPL_WIDTH - 1),
		13674 => to_unsigned(31667, LUT_AMPL_WIDTH - 1),
		13675 => to_unsigned(31668, LUT_AMPL_WIDTH - 1),
		13676 => to_unsigned(31669, LUT_AMPL_WIDTH - 1),
		13677 => to_unsigned(31670, LUT_AMPL_WIDTH - 1),
		13678 => to_unsigned(31670, LUT_AMPL_WIDTH - 1),
		13679 => to_unsigned(31671, LUT_AMPL_WIDTH - 1),
		13680 => to_unsigned(31672, LUT_AMPL_WIDTH - 1),
		13681 => to_unsigned(31673, LUT_AMPL_WIDTH - 1),
		13682 => to_unsigned(31674, LUT_AMPL_WIDTH - 1),
		13683 => to_unsigned(31674, LUT_AMPL_WIDTH - 1),
		13684 => to_unsigned(31675, LUT_AMPL_WIDTH - 1),
		13685 => to_unsigned(31676, LUT_AMPL_WIDTH - 1),
		13686 => to_unsigned(31677, LUT_AMPL_WIDTH - 1),
		13687 => to_unsigned(31678, LUT_AMPL_WIDTH - 1),
		13688 => to_unsigned(31679, LUT_AMPL_WIDTH - 1),
		13689 => to_unsigned(31679, LUT_AMPL_WIDTH - 1),
		13690 => to_unsigned(31680, LUT_AMPL_WIDTH - 1),
		13691 => to_unsigned(31681, LUT_AMPL_WIDTH - 1),
		13692 => to_unsigned(31682, LUT_AMPL_WIDTH - 1),
		13693 => to_unsigned(31683, LUT_AMPL_WIDTH - 1),
		13694 => to_unsigned(31683, LUT_AMPL_WIDTH - 1),
		13695 => to_unsigned(31684, LUT_AMPL_WIDTH - 1),
		13696 => to_unsigned(31685, LUT_AMPL_WIDTH - 1),
		13697 => to_unsigned(31686, LUT_AMPL_WIDTH - 1),
		13698 => to_unsigned(31687, LUT_AMPL_WIDTH - 1),
		13699 => to_unsigned(31687, LUT_AMPL_WIDTH - 1),
		13700 => to_unsigned(31688, LUT_AMPL_WIDTH - 1),
		13701 => to_unsigned(31689, LUT_AMPL_WIDTH - 1),
		13702 => to_unsigned(31690, LUT_AMPL_WIDTH - 1),
		13703 => to_unsigned(31691, LUT_AMPL_WIDTH - 1),
		13704 => to_unsigned(31691, LUT_AMPL_WIDTH - 1),
		13705 => to_unsigned(31692, LUT_AMPL_WIDTH - 1),
		13706 => to_unsigned(31693, LUT_AMPL_WIDTH - 1),
		13707 => to_unsigned(31694, LUT_AMPL_WIDTH - 1),
		13708 => to_unsigned(31695, LUT_AMPL_WIDTH - 1),
		13709 => to_unsigned(31695, LUT_AMPL_WIDTH - 1),
		13710 => to_unsigned(31696, LUT_AMPL_WIDTH - 1),
		13711 => to_unsigned(31697, LUT_AMPL_WIDTH - 1),
		13712 => to_unsigned(31698, LUT_AMPL_WIDTH - 1),
		13713 => to_unsigned(31698, LUT_AMPL_WIDTH - 1),
		13714 => to_unsigned(31699, LUT_AMPL_WIDTH - 1),
		13715 => to_unsigned(31700, LUT_AMPL_WIDTH - 1),
		13716 => to_unsigned(31701, LUT_AMPL_WIDTH - 1),
		13717 => to_unsigned(31702, LUT_AMPL_WIDTH - 1),
		13718 => to_unsigned(31702, LUT_AMPL_WIDTH - 1),
		13719 => to_unsigned(31703, LUT_AMPL_WIDTH - 1),
		13720 => to_unsigned(31704, LUT_AMPL_WIDTH - 1),
		13721 => to_unsigned(31705, LUT_AMPL_WIDTH - 1),
		13722 => to_unsigned(31706, LUT_AMPL_WIDTH - 1),
		13723 => to_unsigned(31706, LUT_AMPL_WIDTH - 1),
		13724 => to_unsigned(31707, LUT_AMPL_WIDTH - 1),
		13725 => to_unsigned(31708, LUT_AMPL_WIDTH - 1),
		13726 => to_unsigned(31709, LUT_AMPL_WIDTH - 1),
		13727 => to_unsigned(31710, LUT_AMPL_WIDTH - 1),
		13728 => to_unsigned(31710, LUT_AMPL_WIDTH - 1),
		13729 => to_unsigned(31711, LUT_AMPL_WIDTH - 1),
		13730 => to_unsigned(31712, LUT_AMPL_WIDTH - 1),
		13731 => to_unsigned(31713, LUT_AMPL_WIDTH - 1),
		13732 => to_unsigned(31714, LUT_AMPL_WIDTH - 1),
		13733 => to_unsigned(31714, LUT_AMPL_WIDTH - 1),
		13734 => to_unsigned(31715, LUT_AMPL_WIDTH - 1),
		13735 => to_unsigned(31716, LUT_AMPL_WIDTH - 1),
		13736 => to_unsigned(31717, LUT_AMPL_WIDTH - 1),
		13737 => to_unsigned(31718, LUT_AMPL_WIDTH - 1),
		13738 => to_unsigned(31718, LUT_AMPL_WIDTH - 1),
		13739 => to_unsigned(31719, LUT_AMPL_WIDTH - 1),
		13740 => to_unsigned(31720, LUT_AMPL_WIDTH - 1),
		13741 => to_unsigned(31721, LUT_AMPL_WIDTH - 1),
		13742 => to_unsigned(31721, LUT_AMPL_WIDTH - 1),
		13743 => to_unsigned(31722, LUT_AMPL_WIDTH - 1),
		13744 => to_unsigned(31723, LUT_AMPL_WIDTH - 1),
		13745 => to_unsigned(31724, LUT_AMPL_WIDTH - 1),
		13746 => to_unsigned(31725, LUT_AMPL_WIDTH - 1),
		13747 => to_unsigned(31725, LUT_AMPL_WIDTH - 1),
		13748 => to_unsigned(31726, LUT_AMPL_WIDTH - 1),
		13749 => to_unsigned(31727, LUT_AMPL_WIDTH - 1),
		13750 => to_unsigned(31728, LUT_AMPL_WIDTH - 1),
		13751 => to_unsigned(31729, LUT_AMPL_WIDTH - 1),
		13752 => to_unsigned(31729, LUT_AMPL_WIDTH - 1),
		13753 => to_unsigned(31730, LUT_AMPL_WIDTH - 1),
		13754 => to_unsigned(31731, LUT_AMPL_WIDTH - 1),
		13755 => to_unsigned(31732, LUT_AMPL_WIDTH - 1),
		13756 => to_unsigned(31732, LUT_AMPL_WIDTH - 1),
		13757 => to_unsigned(31733, LUT_AMPL_WIDTH - 1),
		13758 => to_unsigned(31734, LUT_AMPL_WIDTH - 1),
		13759 => to_unsigned(31735, LUT_AMPL_WIDTH - 1),
		13760 => to_unsigned(31736, LUT_AMPL_WIDTH - 1),
		13761 => to_unsigned(31736, LUT_AMPL_WIDTH - 1),
		13762 => to_unsigned(31737, LUT_AMPL_WIDTH - 1),
		13763 => to_unsigned(31738, LUT_AMPL_WIDTH - 1),
		13764 => to_unsigned(31739, LUT_AMPL_WIDTH - 1),
		13765 => to_unsigned(31739, LUT_AMPL_WIDTH - 1),
		13766 => to_unsigned(31740, LUT_AMPL_WIDTH - 1),
		13767 => to_unsigned(31741, LUT_AMPL_WIDTH - 1),
		13768 => to_unsigned(31742, LUT_AMPL_WIDTH - 1),
		13769 => to_unsigned(31743, LUT_AMPL_WIDTH - 1),
		13770 => to_unsigned(31743, LUT_AMPL_WIDTH - 1),
		13771 => to_unsigned(31744, LUT_AMPL_WIDTH - 1),
		13772 => to_unsigned(31745, LUT_AMPL_WIDTH - 1),
		13773 => to_unsigned(31746, LUT_AMPL_WIDTH - 1),
		13774 => to_unsigned(31746, LUT_AMPL_WIDTH - 1),
		13775 => to_unsigned(31747, LUT_AMPL_WIDTH - 1),
		13776 => to_unsigned(31748, LUT_AMPL_WIDTH - 1),
		13777 => to_unsigned(31749, LUT_AMPL_WIDTH - 1),
		13778 => to_unsigned(31750, LUT_AMPL_WIDTH - 1),
		13779 => to_unsigned(31750, LUT_AMPL_WIDTH - 1),
		13780 => to_unsigned(31751, LUT_AMPL_WIDTH - 1),
		13781 => to_unsigned(31752, LUT_AMPL_WIDTH - 1),
		13782 => to_unsigned(31753, LUT_AMPL_WIDTH - 1),
		13783 => to_unsigned(31753, LUT_AMPL_WIDTH - 1),
		13784 => to_unsigned(31754, LUT_AMPL_WIDTH - 1),
		13785 => to_unsigned(31755, LUT_AMPL_WIDTH - 1),
		13786 => to_unsigned(31756, LUT_AMPL_WIDTH - 1),
		13787 => to_unsigned(31757, LUT_AMPL_WIDTH - 1),
		13788 => to_unsigned(31757, LUT_AMPL_WIDTH - 1),
		13789 => to_unsigned(31758, LUT_AMPL_WIDTH - 1),
		13790 => to_unsigned(31759, LUT_AMPL_WIDTH - 1),
		13791 => to_unsigned(31760, LUT_AMPL_WIDTH - 1),
		13792 => to_unsigned(31760, LUT_AMPL_WIDTH - 1),
		13793 => to_unsigned(31761, LUT_AMPL_WIDTH - 1),
		13794 => to_unsigned(31762, LUT_AMPL_WIDTH - 1),
		13795 => to_unsigned(31763, LUT_AMPL_WIDTH - 1),
		13796 => to_unsigned(31764, LUT_AMPL_WIDTH - 1),
		13797 => to_unsigned(31764, LUT_AMPL_WIDTH - 1),
		13798 => to_unsigned(31765, LUT_AMPL_WIDTH - 1),
		13799 => to_unsigned(31766, LUT_AMPL_WIDTH - 1),
		13800 => to_unsigned(31767, LUT_AMPL_WIDTH - 1),
		13801 => to_unsigned(31767, LUT_AMPL_WIDTH - 1),
		13802 => to_unsigned(31768, LUT_AMPL_WIDTH - 1),
		13803 => to_unsigned(31769, LUT_AMPL_WIDTH - 1),
		13804 => to_unsigned(31770, LUT_AMPL_WIDTH - 1),
		13805 => to_unsigned(31770, LUT_AMPL_WIDTH - 1),
		13806 => to_unsigned(31771, LUT_AMPL_WIDTH - 1),
		13807 => to_unsigned(31772, LUT_AMPL_WIDTH - 1),
		13808 => to_unsigned(31773, LUT_AMPL_WIDTH - 1),
		13809 => to_unsigned(31774, LUT_AMPL_WIDTH - 1),
		13810 => to_unsigned(31774, LUT_AMPL_WIDTH - 1),
		13811 => to_unsigned(31775, LUT_AMPL_WIDTH - 1),
		13812 => to_unsigned(31776, LUT_AMPL_WIDTH - 1),
		13813 => to_unsigned(31777, LUT_AMPL_WIDTH - 1),
		13814 => to_unsigned(31777, LUT_AMPL_WIDTH - 1),
		13815 => to_unsigned(31778, LUT_AMPL_WIDTH - 1),
		13816 => to_unsigned(31779, LUT_AMPL_WIDTH - 1),
		13817 => to_unsigned(31780, LUT_AMPL_WIDTH - 1),
		13818 => to_unsigned(31780, LUT_AMPL_WIDTH - 1),
		13819 => to_unsigned(31781, LUT_AMPL_WIDTH - 1),
		13820 => to_unsigned(31782, LUT_AMPL_WIDTH - 1),
		13821 => to_unsigned(31783, LUT_AMPL_WIDTH - 1),
		13822 => to_unsigned(31783, LUT_AMPL_WIDTH - 1),
		13823 => to_unsigned(31784, LUT_AMPL_WIDTH - 1),
		13824 => to_unsigned(31785, LUT_AMPL_WIDTH - 1),
		13825 => to_unsigned(31786, LUT_AMPL_WIDTH - 1),
		13826 => to_unsigned(31787, LUT_AMPL_WIDTH - 1),
		13827 => to_unsigned(31787, LUT_AMPL_WIDTH - 1),
		13828 => to_unsigned(31788, LUT_AMPL_WIDTH - 1),
		13829 => to_unsigned(31789, LUT_AMPL_WIDTH - 1),
		13830 => to_unsigned(31790, LUT_AMPL_WIDTH - 1),
		13831 => to_unsigned(31790, LUT_AMPL_WIDTH - 1),
		13832 => to_unsigned(31791, LUT_AMPL_WIDTH - 1),
		13833 => to_unsigned(31792, LUT_AMPL_WIDTH - 1),
		13834 => to_unsigned(31793, LUT_AMPL_WIDTH - 1),
		13835 => to_unsigned(31793, LUT_AMPL_WIDTH - 1),
		13836 => to_unsigned(31794, LUT_AMPL_WIDTH - 1),
		13837 => to_unsigned(31795, LUT_AMPL_WIDTH - 1),
		13838 => to_unsigned(31796, LUT_AMPL_WIDTH - 1),
		13839 => to_unsigned(31796, LUT_AMPL_WIDTH - 1),
		13840 => to_unsigned(31797, LUT_AMPL_WIDTH - 1),
		13841 => to_unsigned(31798, LUT_AMPL_WIDTH - 1),
		13842 => to_unsigned(31799, LUT_AMPL_WIDTH - 1),
		13843 => to_unsigned(31799, LUT_AMPL_WIDTH - 1),
		13844 => to_unsigned(31800, LUT_AMPL_WIDTH - 1),
		13845 => to_unsigned(31801, LUT_AMPL_WIDTH - 1),
		13846 => to_unsigned(31802, LUT_AMPL_WIDTH - 1),
		13847 => to_unsigned(31802, LUT_AMPL_WIDTH - 1),
		13848 => to_unsigned(31803, LUT_AMPL_WIDTH - 1),
		13849 => to_unsigned(31804, LUT_AMPL_WIDTH - 1),
		13850 => to_unsigned(31805, LUT_AMPL_WIDTH - 1),
		13851 => to_unsigned(31806, LUT_AMPL_WIDTH - 1),
		13852 => to_unsigned(31806, LUT_AMPL_WIDTH - 1),
		13853 => to_unsigned(31807, LUT_AMPL_WIDTH - 1),
		13854 => to_unsigned(31808, LUT_AMPL_WIDTH - 1),
		13855 => to_unsigned(31809, LUT_AMPL_WIDTH - 1),
		13856 => to_unsigned(31809, LUT_AMPL_WIDTH - 1),
		13857 => to_unsigned(31810, LUT_AMPL_WIDTH - 1),
		13858 => to_unsigned(31811, LUT_AMPL_WIDTH - 1),
		13859 => to_unsigned(31812, LUT_AMPL_WIDTH - 1),
		13860 => to_unsigned(31812, LUT_AMPL_WIDTH - 1),
		13861 => to_unsigned(31813, LUT_AMPL_WIDTH - 1),
		13862 => to_unsigned(31814, LUT_AMPL_WIDTH - 1),
		13863 => to_unsigned(31815, LUT_AMPL_WIDTH - 1),
		13864 => to_unsigned(31815, LUT_AMPL_WIDTH - 1),
		13865 => to_unsigned(31816, LUT_AMPL_WIDTH - 1),
		13866 => to_unsigned(31817, LUT_AMPL_WIDTH - 1),
		13867 => to_unsigned(31818, LUT_AMPL_WIDTH - 1),
		13868 => to_unsigned(31818, LUT_AMPL_WIDTH - 1),
		13869 => to_unsigned(31819, LUT_AMPL_WIDTH - 1),
		13870 => to_unsigned(31820, LUT_AMPL_WIDTH - 1),
		13871 => to_unsigned(31821, LUT_AMPL_WIDTH - 1),
		13872 => to_unsigned(31821, LUT_AMPL_WIDTH - 1),
		13873 => to_unsigned(31822, LUT_AMPL_WIDTH - 1),
		13874 => to_unsigned(31823, LUT_AMPL_WIDTH - 1),
		13875 => to_unsigned(31824, LUT_AMPL_WIDTH - 1),
		13876 => to_unsigned(31824, LUT_AMPL_WIDTH - 1),
		13877 => to_unsigned(31825, LUT_AMPL_WIDTH - 1),
		13878 => to_unsigned(31826, LUT_AMPL_WIDTH - 1),
		13879 => to_unsigned(31827, LUT_AMPL_WIDTH - 1),
		13880 => to_unsigned(31827, LUT_AMPL_WIDTH - 1),
		13881 => to_unsigned(31828, LUT_AMPL_WIDTH - 1),
		13882 => to_unsigned(31829, LUT_AMPL_WIDTH - 1),
		13883 => to_unsigned(31830, LUT_AMPL_WIDTH - 1),
		13884 => to_unsigned(31830, LUT_AMPL_WIDTH - 1),
		13885 => to_unsigned(31831, LUT_AMPL_WIDTH - 1),
		13886 => to_unsigned(31832, LUT_AMPL_WIDTH - 1),
		13887 => to_unsigned(31833, LUT_AMPL_WIDTH - 1),
		13888 => to_unsigned(31833, LUT_AMPL_WIDTH - 1),
		13889 => to_unsigned(31834, LUT_AMPL_WIDTH - 1),
		13890 => to_unsigned(31835, LUT_AMPL_WIDTH - 1),
		13891 => to_unsigned(31836, LUT_AMPL_WIDTH - 1),
		13892 => to_unsigned(31836, LUT_AMPL_WIDTH - 1),
		13893 => to_unsigned(31837, LUT_AMPL_WIDTH - 1),
		13894 => to_unsigned(31838, LUT_AMPL_WIDTH - 1),
		13895 => to_unsigned(31838, LUT_AMPL_WIDTH - 1),
		13896 => to_unsigned(31839, LUT_AMPL_WIDTH - 1),
		13897 => to_unsigned(31840, LUT_AMPL_WIDTH - 1),
		13898 => to_unsigned(31841, LUT_AMPL_WIDTH - 1),
		13899 => to_unsigned(31841, LUT_AMPL_WIDTH - 1),
		13900 => to_unsigned(31842, LUT_AMPL_WIDTH - 1),
		13901 => to_unsigned(31843, LUT_AMPL_WIDTH - 1),
		13902 => to_unsigned(31844, LUT_AMPL_WIDTH - 1),
		13903 => to_unsigned(31844, LUT_AMPL_WIDTH - 1),
		13904 => to_unsigned(31845, LUT_AMPL_WIDTH - 1),
		13905 => to_unsigned(31846, LUT_AMPL_WIDTH - 1),
		13906 => to_unsigned(31847, LUT_AMPL_WIDTH - 1),
		13907 => to_unsigned(31847, LUT_AMPL_WIDTH - 1),
		13908 => to_unsigned(31848, LUT_AMPL_WIDTH - 1),
		13909 => to_unsigned(31849, LUT_AMPL_WIDTH - 1),
		13910 => to_unsigned(31850, LUT_AMPL_WIDTH - 1),
		13911 => to_unsigned(31850, LUT_AMPL_WIDTH - 1),
		13912 => to_unsigned(31851, LUT_AMPL_WIDTH - 1),
		13913 => to_unsigned(31852, LUT_AMPL_WIDTH - 1),
		13914 => to_unsigned(31853, LUT_AMPL_WIDTH - 1),
		13915 => to_unsigned(31853, LUT_AMPL_WIDTH - 1),
		13916 => to_unsigned(31854, LUT_AMPL_WIDTH - 1),
		13917 => to_unsigned(31855, LUT_AMPL_WIDTH - 1),
		13918 => to_unsigned(31855, LUT_AMPL_WIDTH - 1),
		13919 => to_unsigned(31856, LUT_AMPL_WIDTH - 1),
		13920 => to_unsigned(31857, LUT_AMPL_WIDTH - 1),
		13921 => to_unsigned(31858, LUT_AMPL_WIDTH - 1),
		13922 => to_unsigned(31858, LUT_AMPL_WIDTH - 1),
		13923 => to_unsigned(31859, LUT_AMPL_WIDTH - 1),
		13924 => to_unsigned(31860, LUT_AMPL_WIDTH - 1),
		13925 => to_unsigned(31861, LUT_AMPL_WIDTH - 1),
		13926 => to_unsigned(31861, LUT_AMPL_WIDTH - 1),
		13927 => to_unsigned(31862, LUT_AMPL_WIDTH - 1),
		13928 => to_unsigned(31863, LUT_AMPL_WIDTH - 1),
		13929 => to_unsigned(31864, LUT_AMPL_WIDTH - 1),
		13930 => to_unsigned(31864, LUT_AMPL_WIDTH - 1),
		13931 => to_unsigned(31865, LUT_AMPL_WIDTH - 1),
		13932 => to_unsigned(31866, LUT_AMPL_WIDTH - 1),
		13933 => to_unsigned(31866, LUT_AMPL_WIDTH - 1),
		13934 => to_unsigned(31867, LUT_AMPL_WIDTH - 1),
		13935 => to_unsigned(31868, LUT_AMPL_WIDTH - 1),
		13936 => to_unsigned(31869, LUT_AMPL_WIDTH - 1),
		13937 => to_unsigned(31869, LUT_AMPL_WIDTH - 1),
		13938 => to_unsigned(31870, LUT_AMPL_WIDTH - 1),
		13939 => to_unsigned(31871, LUT_AMPL_WIDTH - 1),
		13940 => to_unsigned(31872, LUT_AMPL_WIDTH - 1),
		13941 => to_unsigned(31872, LUT_AMPL_WIDTH - 1),
		13942 => to_unsigned(31873, LUT_AMPL_WIDTH - 1),
		13943 => to_unsigned(31874, LUT_AMPL_WIDTH - 1),
		13944 => to_unsigned(31875, LUT_AMPL_WIDTH - 1),
		13945 => to_unsigned(31875, LUT_AMPL_WIDTH - 1),
		13946 => to_unsigned(31876, LUT_AMPL_WIDTH - 1),
		13947 => to_unsigned(31877, LUT_AMPL_WIDTH - 1),
		13948 => to_unsigned(31877, LUT_AMPL_WIDTH - 1),
		13949 => to_unsigned(31878, LUT_AMPL_WIDTH - 1),
		13950 => to_unsigned(31879, LUT_AMPL_WIDTH - 1),
		13951 => to_unsigned(31880, LUT_AMPL_WIDTH - 1),
		13952 => to_unsigned(31880, LUT_AMPL_WIDTH - 1),
		13953 => to_unsigned(31881, LUT_AMPL_WIDTH - 1),
		13954 => to_unsigned(31882, LUT_AMPL_WIDTH - 1),
		13955 => to_unsigned(31882, LUT_AMPL_WIDTH - 1),
		13956 => to_unsigned(31883, LUT_AMPL_WIDTH - 1),
		13957 => to_unsigned(31884, LUT_AMPL_WIDTH - 1),
		13958 => to_unsigned(31885, LUT_AMPL_WIDTH - 1),
		13959 => to_unsigned(31885, LUT_AMPL_WIDTH - 1),
		13960 => to_unsigned(31886, LUT_AMPL_WIDTH - 1),
		13961 => to_unsigned(31887, LUT_AMPL_WIDTH - 1),
		13962 => to_unsigned(31888, LUT_AMPL_WIDTH - 1),
		13963 => to_unsigned(31888, LUT_AMPL_WIDTH - 1),
		13964 => to_unsigned(31889, LUT_AMPL_WIDTH - 1),
		13965 => to_unsigned(31890, LUT_AMPL_WIDTH - 1),
		13966 => to_unsigned(31890, LUT_AMPL_WIDTH - 1),
		13967 => to_unsigned(31891, LUT_AMPL_WIDTH - 1),
		13968 => to_unsigned(31892, LUT_AMPL_WIDTH - 1),
		13969 => to_unsigned(31893, LUT_AMPL_WIDTH - 1),
		13970 => to_unsigned(31893, LUT_AMPL_WIDTH - 1),
		13971 => to_unsigned(31894, LUT_AMPL_WIDTH - 1),
		13972 => to_unsigned(31895, LUT_AMPL_WIDTH - 1),
		13973 => to_unsigned(31896, LUT_AMPL_WIDTH - 1),
		13974 => to_unsigned(31896, LUT_AMPL_WIDTH - 1),
		13975 => to_unsigned(31897, LUT_AMPL_WIDTH - 1),
		13976 => to_unsigned(31898, LUT_AMPL_WIDTH - 1),
		13977 => to_unsigned(31898, LUT_AMPL_WIDTH - 1),
		13978 => to_unsigned(31899, LUT_AMPL_WIDTH - 1),
		13979 => to_unsigned(31900, LUT_AMPL_WIDTH - 1),
		13980 => to_unsigned(31901, LUT_AMPL_WIDTH - 1),
		13981 => to_unsigned(31901, LUT_AMPL_WIDTH - 1),
		13982 => to_unsigned(31902, LUT_AMPL_WIDTH - 1),
		13983 => to_unsigned(31903, LUT_AMPL_WIDTH - 1),
		13984 => to_unsigned(31903, LUT_AMPL_WIDTH - 1),
		13985 => to_unsigned(31904, LUT_AMPL_WIDTH - 1),
		13986 => to_unsigned(31905, LUT_AMPL_WIDTH - 1),
		13987 => to_unsigned(31906, LUT_AMPL_WIDTH - 1),
		13988 => to_unsigned(31906, LUT_AMPL_WIDTH - 1),
		13989 => to_unsigned(31907, LUT_AMPL_WIDTH - 1),
		13990 => to_unsigned(31908, LUT_AMPL_WIDTH - 1),
		13991 => to_unsigned(31908, LUT_AMPL_WIDTH - 1),
		13992 => to_unsigned(31909, LUT_AMPL_WIDTH - 1),
		13993 => to_unsigned(31910, LUT_AMPL_WIDTH - 1),
		13994 => to_unsigned(31911, LUT_AMPL_WIDTH - 1),
		13995 => to_unsigned(31911, LUT_AMPL_WIDTH - 1),
		13996 => to_unsigned(31912, LUT_AMPL_WIDTH - 1),
		13997 => to_unsigned(31913, LUT_AMPL_WIDTH - 1),
		13998 => to_unsigned(31913, LUT_AMPL_WIDTH - 1),
		13999 => to_unsigned(31914, LUT_AMPL_WIDTH - 1),
		14000 => to_unsigned(31915, LUT_AMPL_WIDTH - 1),
		14001 => to_unsigned(31916, LUT_AMPL_WIDTH - 1),
		14002 => to_unsigned(31916, LUT_AMPL_WIDTH - 1),
		14003 => to_unsigned(31917, LUT_AMPL_WIDTH - 1),
		14004 => to_unsigned(31918, LUT_AMPL_WIDTH - 1),
		14005 => to_unsigned(31918, LUT_AMPL_WIDTH - 1),
		14006 => to_unsigned(31919, LUT_AMPL_WIDTH - 1),
		14007 => to_unsigned(31920, LUT_AMPL_WIDTH - 1),
		14008 => to_unsigned(31921, LUT_AMPL_WIDTH - 1),
		14009 => to_unsigned(31921, LUT_AMPL_WIDTH - 1),
		14010 => to_unsigned(31922, LUT_AMPL_WIDTH - 1),
		14011 => to_unsigned(31923, LUT_AMPL_WIDTH - 1),
		14012 => to_unsigned(31923, LUT_AMPL_WIDTH - 1),
		14013 => to_unsigned(31924, LUT_AMPL_WIDTH - 1),
		14014 => to_unsigned(31925, LUT_AMPL_WIDTH - 1),
		14015 => to_unsigned(31925, LUT_AMPL_WIDTH - 1),
		14016 => to_unsigned(31926, LUT_AMPL_WIDTH - 1),
		14017 => to_unsigned(31927, LUT_AMPL_WIDTH - 1),
		14018 => to_unsigned(31928, LUT_AMPL_WIDTH - 1),
		14019 => to_unsigned(31928, LUT_AMPL_WIDTH - 1),
		14020 => to_unsigned(31929, LUT_AMPL_WIDTH - 1),
		14021 => to_unsigned(31930, LUT_AMPL_WIDTH - 1),
		14022 => to_unsigned(31930, LUT_AMPL_WIDTH - 1),
		14023 => to_unsigned(31931, LUT_AMPL_WIDTH - 1),
		14024 => to_unsigned(31932, LUT_AMPL_WIDTH - 1),
		14025 => to_unsigned(31933, LUT_AMPL_WIDTH - 1),
		14026 => to_unsigned(31933, LUT_AMPL_WIDTH - 1),
		14027 => to_unsigned(31934, LUT_AMPL_WIDTH - 1),
		14028 => to_unsigned(31935, LUT_AMPL_WIDTH - 1),
		14029 => to_unsigned(31935, LUT_AMPL_WIDTH - 1),
		14030 => to_unsigned(31936, LUT_AMPL_WIDTH - 1),
		14031 => to_unsigned(31937, LUT_AMPL_WIDTH - 1),
		14032 => to_unsigned(31937, LUT_AMPL_WIDTH - 1),
		14033 => to_unsigned(31938, LUT_AMPL_WIDTH - 1),
		14034 => to_unsigned(31939, LUT_AMPL_WIDTH - 1),
		14035 => to_unsigned(31940, LUT_AMPL_WIDTH - 1),
		14036 => to_unsigned(31940, LUT_AMPL_WIDTH - 1),
		14037 => to_unsigned(31941, LUT_AMPL_WIDTH - 1),
		14038 => to_unsigned(31942, LUT_AMPL_WIDTH - 1),
		14039 => to_unsigned(31942, LUT_AMPL_WIDTH - 1),
		14040 => to_unsigned(31943, LUT_AMPL_WIDTH - 1),
		14041 => to_unsigned(31944, LUT_AMPL_WIDTH - 1),
		14042 => to_unsigned(31944, LUT_AMPL_WIDTH - 1),
		14043 => to_unsigned(31945, LUT_AMPL_WIDTH - 1),
		14044 => to_unsigned(31946, LUT_AMPL_WIDTH - 1),
		14045 => to_unsigned(31947, LUT_AMPL_WIDTH - 1),
		14046 => to_unsigned(31947, LUT_AMPL_WIDTH - 1),
		14047 => to_unsigned(31948, LUT_AMPL_WIDTH - 1),
		14048 => to_unsigned(31949, LUT_AMPL_WIDTH - 1),
		14049 => to_unsigned(31949, LUT_AMPL_WIDTH - 1),
		14050 => to_unsigned(31950, LUT_AMPL_WIDTH - 1),
		14051 => to_unsigned(31951, LUT_AMPL_WIDTH - 1),
		14052 => to_unsigned(31951, LUT_AMPL_WIDTH - 1),
		14053 => to_unsigned(31952, LUT_AMPL_WIDTH - 1),
		14054 => to_unsigned(31953, LUT_AMPL_WIDTH - 1),
		14055 => to_unsigned(31954, LUT_AMPL_WIDTH - 1),
		14056 => to_unsigned(31954, LUT_AMPL_WIDTH - 1),
		14057 => to_unsigned(31955, LUT_AMPL_WIDTH - 1),
		14058 => to_unsigned(31956, LUT_AMPL_WIDTH - 1),
		14059 => to_unsigned(31956, LUT_AMPL_WIDTH - 1),
		14060 => to_unsigned(31957, LUT_AMPL_WIDTH - 1),
		14061 => to_unsigned(31958, LUT_AMPL_WIDTH - 1),
		14062 => to_unsigned(31958, LUT_AMPL_WIDTH - 1),
		14063 => to_unsigned(31959, LUT_AMPL_WIDTH - 1),
		14064 => to_unsigned(31960, LUT_AMPL_WIDTH - 1),
		14065 => to_unsigned(31960, LUT_AMPL_WIDTH - 1),
		14066 => to_unsigned(31961, LUT_AMPL_WIDTH - 1),
		14067 => to_unsigned(31962, LUT_AMPL_WIDTH - 1),
		14068 => to_unsigned(31963, LUT_AMPL_WIDTH - 1),
		14069 => to_unsigned(31963, LUT_AMPL_WIDTH - 1),
		14070 => to_unsigned(31964, LUT_AMPL_WIDTH - 1),
		14071 => to_unsigned(31965, LUT_AMPL_WIDTH - 1),
		14072 => to_unsigned(31965, LUT_AMPL_WIDTH - 1),
		14073 => to_unsigned(31966, LUT_AMPL_WIDTH - 1),
		14074 => to_unsigned(31967, LUT_AMPL_WIDTH - 1),
		14075 => to_unsigned(31967, LUT_AMPL_WIDTH - 1),
		14076 => to_unsigned(31968, LUT_AMPL_WIDTH - 1),
		14077 => to_unsigned(31969, LUT_AMPL_WIDTH - 1),
		14078 => to_unsigned(31969, LUT_AMPL_WIDTH - 1),
		14079 => to_unsigned(31970, LUT_AMPL_WIDTH - 1),
		14080 => to_unsigned(31971, LUT_AMPL_WIDTH - 1),
		14081 => to_unsigned(31972, LUT_AMPL_WIDTH - 1),
		14082 => to_unsigned(31972, LUT_AMPL_WIDTH - 1),
		14083 => to_unsigned(31973, LUT_AMPL_WIDTH - 1),
		14084 => to_unsigned(31974, LUT_AMPL_WIDTH - 1),
		14085 => to_unsigned(31974, LUT_AMPL_WIDTH - 1),
		14086 => to_unsigned(31975, LUT_AMPL_WIDTH - 1),
		14087 => to_unsigned(31976, LUT_AMPL_WIDTH - 1),
		14088 => to_unsigned(31976, LUT_AMPL_WIDTH - 1),
		14089 => to_unsigned(31977, LUT_AMPL_WIDTH - 1),
		14090 => to_unsigned(31978, LUT_AMPL_WIDTH - 1),
		14091 => to_unsigned(31978, LUT_AMPL_WIDTH - 1),
		14092 => to_unsigned(31979, LUT_AMPL_WIDTH - 1),
		14093 => to_unsigned(31980, LUT_AMPL_WIDTH - 1),
		14094 => to_unsigned(31980, LUT_AMPL_WIDTH - 1),
		14095 => to_unsigned(31981, LUT_AMPL_WIDTH - 1),
		14096 => to_unsigned(31982, LUT_AMPL_WIDTH - 1),
		14097 => to_unsigned(31982, LUT_AMPL_WIDTH - 1),
		14098 => to_unsigned(31983, LUT_AMPL_WIDTH - 1),
		14099 => to_unsigned(31984, LUT_AMPL_WIDTH - 1),
		14100 => to_unsigned(31985, LUT_AMPL_WIDTH - 1),
		14101 => to_unsigned(31985, LUT_AMPL_WIDTH - 1),
		14102 => to_unsigned(31986, LUT_AMPL_WIDTH - 1),
		14103 => to_unsigned(31987, LUT_AMPL_WIDTH - 1),
		14104 => to_unsigned(31987, LUT_AMPL_WIDTH - 1),
		14105 => to_unsigned(31988, LUT_AMPL_WIDTH - 1),
		14106 => to_unsigned(31989, LUT_AMPL_WIDTH - 1),
		14107 => to_unsigned(31989, LUT_AMPL_WIDTH - 1),
		14108 => to_unsigned(31990, LUT_AMPL_WIDTH - 1),
		14109 => to_unsigned(31991, LUT_AMPL_WIDTH - 1),
		14110 => to_unsigned(31991, LUT_AMPL_WIDTH - 1),
		14111 => to_unsigned(31992, LUT_AMPL_WIDTH - 1),
		14112 => to_unsigned(31993, LUT_AMPL_WIDTH - 1),
		14113 => to_unsigned(31993, LUT_AMPL_WIDTH - 1),
		14114 => to_unsigned(31994, LUT_AMPL_WIDTH - 1),
		14115 => to_unsigned(31995, LUT_AMPL_WIDTH - 1),
		14116 => to_unsigned(31995, LUT_AMPL_WIDTH - 1),
		14117 => to_unsigned(31996, LUT_AMPL_WIDTH - 1),
		14118 => to_unsigned(31997, LUT_AMPL_WIDTH - 1),
		14119 => to_unsigned(31997, LUT_AMPL_WIDTH - 1),
		14120 => to_unsigned(31998, LUT_AMPL_WIDTH - 1),
		14121 => to_unsigned(31999, LUT_AMPL_WIDTH - 1),
		14122 => to_unsigned(31999, LUT_AMPL_WIDTH - 1),
		14123 => to_unsigned(32000, LUT_AMPL_WIDTH - 1),
		14124 => to_unsigned(32001, LUT_AMPL_WIDTH - 1),
		14125 => to_unsigned(32002, LUT_AMPL_WIDTH - 1),
		14126 => to_unsigned(32002, LUT_AMPL_WIDTH - 1),
		14127 => to_unsigned(32003, LUT_AMPL_WIDTH - 1),
		14128 => to_unsigned(32004, LUT_AMPL_WIDTH - 1),
		14129 => to_unsigned(32004, LUT_AMPL_WIDTH - 1),
		14130 => to_unsigned(32005, LUT_AMPL_WIDTH - 1),
		14131 => to_unsigned(32006, LUT_AMPL_WIDTH - 1),
		14132 => to_unsigned(32006, LUT_AMPL_WIDTH - 1),
		14133 => to_unsigned(32007, LUT_AMPL_WIDTH - 1),
		14134 => to_unsigned(32008, LUT_AMPL_WIDTH - 1),
		14135 => to_unsigned(32008, LUT_AMPL_WIDTH - 1),
		14136 => to_unsigned(32009, LUT_AMPL_WIDTH - 1),
		14137 => to_unsigned(32010, LUT_AMPL_WIDTH - 1),
		14138 => to_unsigned(32010, LUT_AMPL_WIDTH - 1),
		14139 => to_unsigned(32011, LUT_AMPL_WIDTH - 1),
		14140 => to_unsigned(32012, LUT_AMPL_WIDTH - 1),
		14141 => to_unsigned(32012, LUT_AMPL_WIDTH - 1),
		14142 => to_unsigned(32013, LUT_AMPL_WIDTH - 1),
		14143 => to_unsigned(32014, LUT_AMPL_WIDTH - 1),
		14144 => to_unsigned(32014, LUT_AMPL_WIDTH - 1),
		14145 => to_unsigned(32015, LUT_AMPL_WIDTH - 1),
		14146 => to_unsigned(32016, LUT_AMPL_WIDTH - 1),
		14147 => to_unsigned(32016, LUT_AMPL_WIDTH - 1),
		14148 => to_unsigned(32017, LUT_AMPL_WIDTH - 1),
		14149 => to_unsigned(32018, LUT_AMPL_WIDTH - 1),
		14150 => to_unsigned(32018, LUT_AMPL_WIDTH - 1),
		14151 => to_unsigned(32019, LUT_AMPL_WIDTH - 1),
		14152 => to_unsigned(32020, LUT_AMPL_WIDTH - 1),
		14153 => to_unsigned(32020, LUT_AMPL_WIDTH - 1),
		14154 => to_unsigned(32021, LUT_AMPL_WIDTH - 1),
		14155 => to_unsigned(32022, LUT_AMPL_WIDTH - 1),
		14156 => to_unsigned(32022, LUT_AMPL_WIDTH - 1),
		14157 => to_unsigned(32023, LUT_AMPL_WIDTH - 1),
		14158 => to_unsigned(32024, LUT_AMPL_WIDTH - 1),
		14159 => to_unsigned(32024, LUT_AMPL_WIDTH - 1),
		14160 => to_unsigned(32025, LUT_AMPL_WIDTH - 1),
		14161 => to_unsigned(32026, LUT_AMPL_WIDTH - 1),
		14162 => to_unsigned(32026, LUT_AMPL_WIDTH - 1),
		14163 => to_unsigned(32027, LUT_AMPL_WIDTH - 1),
		14164 => to_unsigned(32028, LUT_AMPL_WIDTH - 1),
		14165 => to_unsigned(32028, LUT_AMPL_WIDTH - 1),
		14166 => to_unsigned(32029, LUT_AMPL_WIDTH - 1),
		14167 => to_unsigned(32030, LUT_AMPL_WIDTH - 1),
		14168 => to_unsigned(32030, LUT_AMPL_WIDTH - 1),
		14169 => to_unsigned(32031, LUT_AMPL_WIDTH - 1),
		14170 => to_unsigned(32032, LUT_AMPL_WIDTH - 1),
		14171 => to_unsigned(32032, LUT_AMPL_WIDTH - 1),
		14172 => to_unsigned(32033, LUT_AMPL_WIDTH - 1),
		14173 => to_unsigned(32034, LUT_AMPL_WIDTH - 1),
		14174 => to_unsigned(32034, LUT_AMPL_WIDTH - 1),
		14175 => to_unsigned(32035, LUT_AMPL_WIDTH - 1),
		14176 => to_unsigned(32036, LUT_AMPL_WIDTH - 1),
		14177 => to_unsigned(32036, LUT_AMPL_WIDTH - 1),
		14178 => to_unsigned(32037, LUT_AMPL_WIDTH - 1),
		14179 => to_unsigned(32038, LUT_AMPL_WIDTH - 1),
		14180 => to_unsigned(32038, LUT_AMPL_WIDTH - 1),
		14181 => to_unsigned(32039, LUT_AMPL_WIDTH - 1),
		14182 => to_unsigned(32040, LUT_AMPL_WIDTH - 1),
		14183 => to_unsigned(32040, LUT_AMPL_WIDTH - 1),
		14184 => to_unsigned(32041, LUT_AMPL_WIDTH - 1),
		14185 => to_unsigned(32041, LUT_AMPL_WIDTH - 1),
		14186 => to_unsigned(32042, LUT_AMPL_WIDTH - 1),
		14187 => to_unsigned(32043, LUT_AMPL_WIDTH - 1),
		14188 => to_unsigned(32043, LUT_AMPL_WIDTH - 1),
		14189 => to_unsigned(32044, LUT_AMPL_WIDTH - 1),
		14190 => to_unsigned(32045, LUT_AMPL_WIDTH - 1),
		14191 => to_unsigned(32045, LUT_AMPL_WIDTH - 1),
		14192 => to_unsigned(32046, LUT_AMPL_WIDTH - 1),
		14193 => to_unsigned(32047, LUT_AMPL_WIDTH - 1),
		14194 => to_unsigned(32047, LUT_AMPL_WIDTH - 1),
		14195 => to_unsigned(32048, LUT_AMPL_WIDTH - 1),
		14196 => to_unsigned(32049, LUT_AMPL_WIDTH - 1),
		14197 => to_unsigned(32049, LUT_AMPL_WIDTH - 1),
		14198 => to_unsigned(32050, LUT_AMPL_WIDTH - 1),
		14199 => to_unsigned(32051, LUT_AMPL_WIDTH - 1),
		14200 => to_unsigned(32051, LUT_AMPL_WIDTH - 1),
		14201 => to_unsigned(32052, LUT_AMPL_WIDTH - 1),
		14202 => to_unsigned(32053, LUT_AMPL_WIDTH - 1),
		14203 => to_unsigned(32053, LUT_AMPL_WIDTH - 1),
		14204 => to_unsigned(32054, LUT_AMPL_WIDTH - 1),
		14205 => to_unsigned(32055, LUT_AMPL_WIDTH - 1),
		14206 => to_unsigned(32055, LUT_AMPL_WIDTH - 1),
		14207 => to_unsigned(32056, LUT_AMPL_WIDTH - 1),
		14208 => to_unsigned(32057, LUT_AMPL_WIDTH - 1),
		14209 => to_unsigned(32057, LUT_AMPL_WIDTH - 1),
		14210 => to_unsigned(32058, LUT_AMPL_WIDTH - 1),
		14211 => to_unsigned(32058, LUT_AMPL_WIDTH - 1),
		14212 => to_unsigned(32059, LUT_AMPL_WIDTH - 1),
		14213 => to_unsigned(32060, LUT_AMPL_WIDTH - 1),
		14214 => to_unsigned(32060, LUT_AMPL_WIDTH - 1),
		14215 => to_unsigned(32061, LUT_AMPL_WIDTH - 1),
		14216 => to_unsigned(32062, LUT_AMPL_WIDTH - 1),
		14217 => to_unsigned(32062, LUT_AMPL_WIDTH - 1),
		14218 => to_unsigned(32063, LUT_AMPL_WIDTH - 1),
		14219 => to_unsigned(32064, LUT_AMPL_WIDTH - 1),
		14220 => to_unsigned(32064, LUT_AMPL_WIDTH - 1),
		14221 => to_unsigned(32065, LUT_AMPL_WIDTH - 1),
		14222 => to_unsigned(32066, LUT_AMPL_WIDTH - 1),
		14223 => to_unsigned(32066, LUT_AMPL_WIDTH - 1),
		14224 => to_unsigned(32067, LUT_AMPL_WIDTH - 1),
		14225 => to_unsigned(32068, LUT_AMPL_WIDTH - 1),
		14226 => to_unsigned(32068, LUT_AMPL_WIDTH - 1),
		14227 => to_unsigned(32069, LUT_AMPL_WIDTH - 1),
		14228 => to_unsigned(32069, LUT_AMPL_WIDTH - 1),
		14229 => to_unsigned(32070, LUT_AMPL_WIDTH - 1),
		14230 => to_unsigned(32071, LUT_AMPL_WIDTH - 1),
		14231 => to_unsigned(32071, LUT_AMPL_WIDTH - 1),
		14232 => to_unsigned(32072, LUT_AMPL_WIDTH - 1),
		14233 => to_unsigned(32073, LUT_AMPL_WIDTH - 1),
		14234 => to_unsigned(32073, LUT_AMPL_WIDTH - 1),
		14235 => to_unsigned(32074, LUT_AMPL_WIDTH - 1),
		14236 => to_unsigned(32075, LUT_AMPL_WIDTH - 1),
		14237 => to_unsigned(32075, LUT_AMPL_WIDTH - 1),
		14238 => to_unsigned(32076, LUT_AMPL_WIDTH - 1),
		14239 => to_unsigned(32077, LUT_AMPL_WIDTH - 1),
		14240 => to_unsigned(32077, LUT_AMPL_WIDTH - 1),
		14241 => to_unsigned(32078, LUT_AMPL_WIDTH - 1),
		14242 => to_unsigned(32078, LUT_AMPL_WIDTH - 1),
		14243 => to_unsigned(32079, LUT_AMPL_WIDTH - 1),
		14244 => to_unsigned(32080, LUT_AMPL_WIDTH - 1),
		14245 => to_unsigned(32080, LUT_AMPL_WIDTH - 1),
		14246 => to_unsigned(32081, LUT_AMPL_WIDTH - 1),
		14247 => to_unsigned(32082, LUT_AMPL_WIDTH - 1),
		14248 => to_unsigned(32082, LUT_AMPL_WIDTH - 1),
		14249 => to_unsigned(32083, LUT_AMPL_WIDTH - 1),
		14250 => to_unsigned(32084, LUT_AMPL_WIDTH - 1),
		14251 => to_unsigned(32084, LUT_AMPL_WIDTH - 1),
		14252 => to_unsigned(32085, LUT_AMPL_WIDTH - 1),
		14253 => to_unsigned(32086, LUT_AMPL_WIDTH - 1),
		14254 => to_unsigned(32086, LUT_AMPL_WIDTH - 1),
		14255 => to_unsigned(32087, LUT_AMPL_WIDTH - 1),
		14256 => to_unsigned(32087, LUT_AMPL_WIDTH - 1),
		14257 => to_unsigned(32088, LUT_AMPL_WIDTH - 1),
		14258 => to_unsigned(32089, LUT_AMPL_WIDTH - 1),
		14259 => to_unsigned(32089, LUT_AMPL_WIDTH - 1),
		14260 => to_unsigned(32090, LUT_AMPL_WIDTH - 1),
		14261 => to_unsigned(32091, LUT_AMPL_WIDTH - 1),
		14262 => to_unsigned(32091, LUT_AMPL_WIDTH - 1),
		14263 => to_unsigned(32092, LUT_AMPL_WIDTH - 1),
		14264 => to_unsigned(32092, LUT_AMPL_WIDTH - 1),
		14265 => to_unsigned(32093, LUT_AMPL_WIDTH - 1),
		14266 => to_unsigned(32094, LUT_AMPL_WIDTH - 1),
		14267 => to_unsigned(32094, LUT_AMPL_WIDTH - 1),
		14268 => to_unsigned(32095, LUT_AMPL_WIDTH - 1),
		14269 => to_unsigned(32096, LUT_AMPL_WIDTH - 1),
		14270 => to_unsigned(32096, LUT_AMPL_WIDTH - 1),
		14271 => to_unsigned(32097, LUT_AMPL_WIDTH - 1),
		14272 => to_unsigned(32098, LUT_AMPL_WIDTH - 1),
		14273 => to_unsigned(32098, LUT_AMPL_WIDTH - 1),
		14274 => to_unsigned(32099, LUT_AMPL_WIDTH - 1),
		14275 => to_unsigned(32099, LUT_AMPL_WIDTH - 1),
		14276 => to_unsigned(32100, LUT_AMPL_WIDTH - 1),
		14277 => to_unsigned(32101, LUT_AMPL_WIDTH - 1),
		14278 => to_unsigned(32101, LUT_AMPL_WIDTH - 1),
		14279 => to_unsigned(32102, LUT_AMPL_WIDTH - 1),
		14280 => to_unsigned(32103, LUT_AMPL_WIDTH - 1),
		14281 => to_unsigned(32103, LUT_AMPL_WIDTH - 1),
		14282 => to_unsigned(32104, LUT_AMPL_WIDTH - 1),
		14283 => to_unsigned(32104, LUT_AMPL_WIDTH - 1),
		14284 => to_unsigned(32105, LUT_AMPL_WIDTH - 1),
		14285 => to_unsigned(32106, LUT_AMPL_WIDTH - 1),
		14286 => to_unsigned(32106, LUT_AMPL_WIDTH - 1),
		14287 => to_unsigned(32107, LUT_AMPL_WIDTH - 1),
		14288 => to_unsigned(32108, LUT_AMPL_WIDTH - 1),
		14289 => to_unsigned(32108, LUT_AMPL_WIDTH - 1),
		14290 => to_unsigned(32109, LUT_AMPL_WIDTH - 1),
		14291 => to_unsigned(32110, LUT_AMPL_WIDTH - 1),
		14292 => to_unsigned(32110, LUT_AMPL_WIDTH - 1),
		14293 => to_unsigned(32111, LUT_AMPL_WIDTH - 1),
		14294 => to_unsigned(32111, LUT_AMPL_WIDTH - 1),
		14295 => to_unsigned(32112, LUT_AMPL_WIDTH - 1),
		14296 => to_unsigned(32113, LUT_AMPL_WIDTH - 1),
		14297 => to_unsigned(32113, LUT_AMPL_WIDTH - 1),
		14298 => to_unsigned(32114, LUT_AMPL_WIDTH - 1),
		14299 => to_unsigned(32115, LUT_AMPL_WIDTH - 1),
		14300 => to_unsigned(32115, LUT_AMPL_WIDTH - 1),
		14301 => to_unsigned(32116, LUT_AMPL_WIDTH - 1),
		14302 => to_unsigned(32116, LUT_AMPL_WIDTH - 1),
		14303 => to_unsigned(32117, LUT_AMPL_WIDTH - 1),
		14304 => to_unsigned(32118, LUT_AMPL_WIDTH - 1),
		14305 => to_unsigned(32118, LUT_AMPL_WIDTH - 1),
		14306 => to_unsigned(32119, LUT_AMPL_WIDTH - 1),
		14307 => to_unsigned(32119, LUT_AMPL_WIDTH - 1),
		14308 => to_unsigned(32120, LUT_AMPL_WIDTH - 1),
		14309 => to_unsigned(32121, LUT_AMPL_WIDTH - 1),
		14310 => to_unsigned(32121, LUT_AMPL_WIDTH - 1),
		14311 => to_unsigned(32122, LUT_AMPL_WIDTH - 1),
		14312 => to_unsigned(32123, LUT_AMPL_WIDTH - 1),
		14313 => to_unsigned(32123, LUT_AMPL_WIDTH - 1),
		14314 => to_unsigned(32124, LUT_AMPL_WIDTH - 1),
		14315 => to_unsigned(32124, LUT_AMPL_WIDTH - 1),
		14316 => to_unsigned(32125, LUT_AMPL_WIDTH - 1),
		14317 => to_unsigned(32126, LUT_AMPL_WIDTH - 1),
		14318 => to_unsigned(32126, LUT_AMPL_WIDTH - 1),
		14319 => to_unsigned(32127, LUT_AMPL_WIDTH - 1),
		14320 => to_unsigned(32128, LUT_AMPL_WIDTH - 1),
		14321 => to_unsigned(32128, LUT_AMPL_WIDTH - 1),
		14322 => to_unsigned(32129, LUT_AMPL_WIDTH - 1),
		14323 => to_unsigned(32129, LUT_AMPL_WIDTH - 1),
		14324 => to_unsigned(32130, LUT_AMPL_WIDTH - 1),
		14325 => to_unsigned(32131, LUT_AMPL_WIDTH - 1),
		14326 => to_unsigned(32131, LUT_AMPL_WIDTH - 1),
		14327 => to_unsigned(32132, LUT_AMPL_WIDTH - 1),
		14328 => to_unsigned(32132, LUT_AMPL_WIDTH - 1),
		14329 => to_unsigned(32133, LUT_AMPL_WIDTH - 1),
		14330 => to_unsigned(32134, LUT_AMPL_WIDTH - 1),
		14331 => to_unsigned(32134, LUT_AMPL_WIDTH - 1),
		14332 => to_unsigned(32135, LUT_AMPL_WIDTH - 1),
		14333 => to_unsigned(32136, LUT_AMPL_WIDTH - 1),
		14334 => to_unsigned(32136, LUT_AMPL_WIDTH - 1),
		14335 => to_unsigned(32137, LUT_AMPL_WIDTH - 1),
		14336 => to_unsigned(32137, LUT_AMPL_WIDTH - 1),
		14337 => to_unsigned(32138, LUT_AMPL_WIDTH - 1),
		14338 => to_unsigned(32139, LUT_AMPL_WIDTH - 1),
		14339 => to_unsigned(32139, LUT_AMPL_WIDTH - 1),
		14340 => to_unsigned(32140, LUT_AMPL_WIDTH - 1),
		14341 => to_unsigned(32140, LUT_AMPL_WIDTH - 1),
		14342 => to_unsigned(32141, LUT_AMPL_WIDTH - 1),
		14343 => to_unsigned(32142, LUT_AMPL_WIDTH - 1),
		14344 => to_unsigned(32142, LUT_AMPL_WIDTH - 1),
		14345 => to_unsigned(32143, LUT_AMPL_WIDTH - 1),
		14346 => to_unsigned(32144, LUT_AMPL_WIDTH - 1),
		14347 => to_unsigned(32144, LUT_AMPL_WIDTH - 1),
		14348 => to_unsigned(32145, LUT_AMPL_WIDTH - 1),
		14349 => to_unsigned(32145, LUT_AMPL_WIDTH - 1),
		14350 => to_unsigned(32146, LUT_AMPL_WIDTH - 1),
		14351 => to_unsigned(32147, LUT_AMPL_WIDTH - 1),
		14352 => to_unsigned(32147, LUT_AMPL_WIDTH - 1),
		14353 => to_unsigned(32148, LUT_AMPL_WIDTH - 1),
		14354 => to_unsigned(32148, LUT_AMPL_WIDTH - 1),
		14355 => to_unsigned(32149, LUT_AMPL_WIDTH - 1),
		14356 => to_unsigned(32150, LUT_AMPL_WIDTH - 1),
		14357 => to_unsigned(32150, LUT_AMPL_WIDTH - 1),
		14358 => to_unsigned(32151, LUT_AMPL_WIDTH - 1),
		14359 => to_unsigned(32151, LUT_AMPL_WIDTH - 1),
		14360 => to_unsigned(32152, LUT_AMPL_WIDTH - 1),
		14361 => to_unsigned(32153, LUT_AMPL_WIDTH - 1),
		14362 => to_unsigned(32153, LUT_AMPL_WIDTH - 1),
		14363 => to_unsigned(32154, LUT_AMPL_WIDTH - 1),
		14364 => to_unsigned(32154, LUT_AMPL_WIDTH - 1),
		14365 => to_unsigned(32155, LUT_AMPL_WIDTH - 1),
		14366 => to_unsigned(32156, LUT_AMPL_WIDTH - 1),
		14367 => to_unsigned(32156, LUT_AMPL_WIDTH - 1),
		14368 => to_unsigned(32157, LUT_AMPL_WIDTH - 1),
		14369 => to_unsigned(32157, LUT_AMPL_WIDTH - 1),
		14370 => to_unsigned(32158, LUT_AMPL_WIDTH - 1),
		14371 => to_unsigned(32159, LUT_AMPL_WIDTH - 1),
		14372 => to_unsigned(32159, LUT_AMPL_WIDTH - 1),
		14373 => to_unsigned(32160, LUT_AMPL_WIDTH - 1),
		14374 => to_unsigned(32160, LUT_AMPL_WIDTH - 1),
		14375 => to_unsigned(32161, LUT_AMPL_WIDTH - 1),
		14376 => to_unsigned(32162, LUT_AMPL_WIDTH - 1),
		14377 => to_unsigned(32162, LUT_AMPL_WIDTH - 1),
		14378 => to_unsigned(32163, LUT_AMPL_WIDTH - 1),
		14379 => to_unsigned(32163, LUT_AMPL_WIDTH - 1),
		14380 => to_unsigned(32164, LUT_AMPL_WIDTH - 1),
		14381 => to_unsigned(32165, LUT_AMPL_WIDTH - 1),
		14382 => to_unsigned(32165, LUT_AMPL_WIDTH - 1),
		14383 => to_unsigned(32166, LUT_AMPL_WIDTH - 1),
		14384 => to_unsigned(32166, LUT_AMPL_WIDTH - 1),
		14385 => to_unsigned(32167, LUT_AMPL_WIDTH - 1),
		14386 => to_unsigned(32168, LUT_AMPL_WIDTH - 1),
		14387 => to_unsigned(32168, LUT_AMPL_WIDTH - 1),
		14388 => to_unsigned(32169, LUT_AMPL_WIDTH - 1),
		14389 => to_unsigned(32169, LUT_AMPL_WIDTH - 1),
		14390 => to_unsigned(32170, LUT_AMPL_WIDTH - 1),
		14391 => to_unsigned(32171, LUT_AMPL_WIDTH - 1),
		14392 => to_unsigned(32171, LUT_AMPL_WIDTH - 1),
		14393 => to_unsigned(32172, LUT_AMPL_WIDTH - 1),
		14394 => to_unsigned(32172, LUT_AMPL_WIDTH - 1),
		14395 => to_unsigned(32173, LUT_AMPL_WIDTH - 1),
		14396 => to_unsigned(32174, LUT_AMPL_WIDTH - 1),
		14397 => to_unsigned(32174, LUT_AMPL_WIDTH - 1),
		14398 => to_unsigned(32175, LUT_AMPL_WIDTH - 1),
		14399 => to_unsigned(32175, LUT_AMPL_WIDTH - 1),
		14400 => to_unsigned(32176, LUT_AMPL_WIDTH - 1),
		14401 => to_unsigned(32177, LUT_AMPL_WIDTH - 1),
		14402 => to_unsigned(32177, LUT_AMPL_WIDTH - 1),
		14403 => to_unsigned(32178, LUT_AMPL_WIDTH - 1),
		14404 => to_unsigned(32178, LUT_AMPL_WIDTH - 1),
		14405 => to_unsigned(32179, LUT_AMPL_WIDTH - 1),
		14406 => to_unsigned(32180, LUT_AMPL_WIDTH - 1),
		14407 => to_unsigned(32180, LUT_AMPL_WIDTH - 1),
		14408 => to_unsigned(32181, LUT_AMPL_WIDTH - 1),
		14409 => to_unsigned(32181, LUT_AMPL_WIDTH - 1),
		14410 => to_unsigned(32182, LUT_AMPL_WIDTH - 1),
		14411 => to_unsigned(32183, LUT_AMPL_WIDTH - 1),
		14412 => to_unsigned(32183, LUT_AMPL_WIDTH - 1),
		14413 => to_unsigned(32184, LUT_AMPL_WIDTH - 1),
		14414 => to_unsigned(32184, LUT_AMPL_WIDTH - 1),
		14415 => to_unsigned(32185, LUT_AMPL_WIDTH - 1),
		14416 => to_unsigned(32185, LUT_AMPL_WIDTH - 1),
		14417 => to_unsigned(32186, LUT_AMPL_WIDTH - 1),
		14418 => to_unsigned(32187, LUT_AMPL_WIDTH - 1),
		14419 => to_unsigned(32187, LUT_AMPL_WIDTH - 1),
		14420 => to_unsigned(32188, LUT_AMPL_WIDTH - 1),
		14421 => to_unsigned(32188, LUT_AMPL_WIDTH - 1),
		14422 => to_unsigned(32189, LUT_AMPL_WIDTH - 1),
		14423 => to_unsigned(32190, LUT_AMPL_WIDTH - 1),
		14424 => to_unsigned(32190, LUT_AMPL_WIDTH - 1),
		14425 => to_unsigned(32191, LUT_AMPL_WIDTH - 1),
		14426 => to_unsigned(32191, LUT_AMPL_WIDTH - 1),
		14427 => to_unsigned(32192, LUT_AMPL_WIDTH - 1),
		14428 => to_unsigned(32193, LUT_AMPL_WIDTH - 1),
		14429 => to_unsigned(32193, LUT_AMPL_WIDTH - 1),
		14430 => to_unsigned(32194, LUT_AMPL_WIDTH - 1),
		14431 => to_unsigned(32194, LUT_AMPL_WIDTH - 1),
		14432 => to_unsigned(32195, LUT_AMPL_WIDTH - 1),
		14433 => to_unsigned(32195, LUT_AMPL_WIDTH - 1),
		14434 => to_unsigned(32196, LUT_AMPL_WIDTH - 1),
		14435 => to_unsigned(32197, LUT_AMPL_WIDTH - 1),
		14436 => to_unsigned(32197, LUT_AMPL_WIDTH - 1),
		14437 => to_unsigned(32198, LUT_AMPL_WIDTH - 1),
		14438 => to_unsigned(32198, LUT_AMPL_WIDTH - 1),
		14439 => to_unsigned(32199, LUT_AMPL_WIDTH - 1),
		14440 => to_unsigned(32200, LUT_AMPL_WIDTH - 1),
		14441 => to_unsigned(32200, LUT_AMPL_WIDTH - 1),
		14442 => to_unsigned(32201, LUT_AMPL_WIDTH - 1),
		14443 => to_unsigned(32201, LUT_AMPL_WIDTH - 1),
		14444 => to_unsigned(32202, LUT_AMPL_WIDTH - 1),
		14445 => to_unsigned(32202, LUT_AMPL_WIDTH - 1),
		14446 => to_unsigned(32203, LUT_AMPL_WIDTH - 1),
		14447 => to_unsigned(32204, LUT_AMPL_WIDTH - 1),
		14448 => to_unsigned(32204, LUT_AMPL_WIDTH - 1),
		14449 => to_unsigned(32205, LUT_AMPL_WIDTH - 1),
		14450 => to_unsigned(32205, LUT_AMPL_WIDTH - 1),
		14451 => to_unsigned(32206, LUT_AMPL_WIDTH - 1),
		14452 => to_unsigned(32206, LUT_AMPL_WIDTH - 1),
		14453 => to_unsigned(32207, LUT_AMPL_WIDTH - 1),
		14454 => to_unsigned(32208, LUT_AMPL_WIDTH - 1),
		14455 => to_unsigned(32208, LUT_AMPL_WIDTH - 1),
		14456 => to_unsigned(32209, LUT_AMPL_WIDTH - 1),
		14457 => to_unsigned(32209, LUT_AMPL_WIDTH - 1),
		14458 => to_unsigned(32210, LUT_AMPL_WIDTH - 1),
		14459 => to_unsigned(32211, LUT_AMPL_WIDTH - 1),
		14460 => to_unsigned(32211, LUT_AMPL_WIDTH - 1),
		14461 => to_unsigned(32212, LUT_AMPL_WIDTH - 1),
		14462 => to_unsigned(32212, LUT_AMPL_WIDTH - 1),
		14463 => to_unsigned(32213, LUT_AMPL_WIDTH - 1),
		14464 => to_unsigned(32213, LUT_AMPL_WIDTH - 1),
		14465 => to_unsigned(32214, LUT_AMPL_WIDTH - 1),
		14466 => to_unsigned(32215, LUT_AMPL_WIDTH - 1),
		14467 => to_unsigned(32215, LUT_AMPL_WIDTH - 1),
		14468 => to_unsigned(32216, LUT_AMPL_WIDTH - 1),
		14469 => to_unsigned(32216, LUT_AMPL_WIDTH - 1),
		14470 => to_unsigned(32217, LUT_AMPL_WIDTH - 1),
		14471 => to_unsigned(32217, LUT_AMPL_WIDTH - 1),
		14472 => to_unsigned(32218, LUT_AMPL_WIDTH - 1),
		14473 => to_unsigned(32219, LUT_AMPL_WIDTH - 1),
		14474 => to_unsigned(32219, LUT_AMPL_WIDTH - 1),
		14475 => to_unsigned(32220, LUT_AMPL_WIDTH - 1),
		14476 => to_unsigned(32220, LUT_AMPL_WIDTH - 1),
		14477 => to_unsigned(32221, LUT_AMPL_WIDTH - 1),
		14478 => to_unsigned(32221, LUT_AMPL_WIDTH - 1),
		14479 => to_unsigned(32222, LUT_AMPL_WIDTH - 1),
		14480 => to_unsigned(32223, LUT_AMPL_WIDTH - 1),
		14481 => to_unsigned(32223, LUT_AMPL_WIDTH - 1),
		14482 => to_unsigned(32224, LUT_AMPL_WIDTH - 1),
		14483 => to_unsigned(32224, LUT_AMPL_WIDTH - 1),
		14484 => to_unsigned(32225, LUT_AMPL_WIDTH - 1),
		14485 => to_unsigned(32225, LUT_AMPL_WIDTH - 1),
		14486 => to_unsigned(32226, LUT_AMPL_WIDTH - 1),
		14487 => to_unsigned(32227, LUT_AMPL_WIDTH - 1),
		14488 => to_unsigned(32227, LUT_AMPL_WIDTH - 1),
		14489 => to_unsigned(32228, LUT_AMPL_WIDTH - 1),
		14490 => to_unsigned(32228, LUT_AMPL_WIDTH - 1),
		14491 => to_unsigned(32229, LUT_AMPL_WIDTH - 1),
		14492 => to_unsigned(32229, LUT_AMPL_WIDTH - 1),
		14493 => to_unsigned(32230, LUT_AMPL_WIDTH - 1),
		14494 => to_unsigned(32231, LUT_AMPL_WIDTH - 1),
		14495 => to_unsigned(32231, LUT_AMPL_WIDTH - 1),
		14496 => to_unsigned(32232, LUT_AMPL_WIDTH - 1),
		14497 => to_unsigned(32232, LUT_AMPL_WIDTH - 1),
		14498 => to_unsigned(32233, LUT_AMPL_WIDTH - 1),
		14499 => to_unsigned(32233, LUT_AMPL_WIDTH - 1),
		14500 => to_unsigned(32234, LUT_AMPL_WIDTH - 1),
		14501 => to_unsigned(32234, LUT_AMPL_WIDTH - 1),
		14502 => to_unsigned(32235, LUT_AMPL_WIDTH - 1),
		14503 => to_unsigned(32236, LUT_AMPL_WIDTH - 1),
		14504 => to_unsigned(32236, LUT_AMPL_WIDTH - 1),
		14505 => to_unsigned(32237, LUT_AMPL_WIDTH - 1),
		14506 => to_unsigned(32237, LUT_AMPL_WIDTH - 1),
		14507 => to_unsigned(32238, LUT_AMPL_WIDTH - 1),
		14508 => to_unsigned(32238, LUT_AMPL_WIDTH - 1),
		14509 => to_unsigned(32239, LUT_AMPL_WIDTH - 1),
		14510 => to_unsigned(32240, LUT_AMPL_WIDTH - 1),
		14511 => to_unsigned(32240, LUT_AMPL_WIDTH - 1),
		14512 => to_unsigned(32241, LUT_AMPL_WIDTH - 1),
		14513 => to_unsigned(32241, LUT_AMPL_WIDTH - 1),
		14514 => to_unsigned(32242, LUT_AMPL_WIDTH - 1),
		14515 => to_unsigned(32242, LUT_AMPL_WIDTH - 1),
		14516 => to_unsigned(32243, LUT_AMPL_WIDTH - 1),
		14517 => to_unsigned(32243, LUT_AMPL_WIDTH - 1),
		14518 => to_unsigned(32244, LUT_AMPL_WIDTH - 1),
		14519 => to_unsigned(32245, LUT_AMPL_WIDTH - 1),
		14520 => to_unsigned(32245, LUT_AMPL_WIDTH - 1),
		14521 => to_unsigned(32246, LUT_AMPL_WIDTH - 1),
		14522 => to_unsigned(32246, LUT_AMPL_WIDTH - 1),
		14523 => to_unsigned(32247, LUT_AMPL_WIDTH - 1),
		14524 => to_unsigned(32247, LUT_AMPL_WIDTH - 1),
		14525 => to_unsigned(32248, LUT_AMPL_WIDTH - 1),
		14526 => to_unsigned(32248, LUT_AMPL_WIDTH - 1),
		14527 => to_unsigned(32249, LUT_AMPL_WIDTH - 1),
		14528 => to_unsigned(32250, LUT_AMPL_WIDTH - 1),
		14529 => to_unsigned(32250, LUT_AMPL_WIDTH - 1),
		14530 => to_unsigned(32251, LUT_AMPL_WIDTH - 1),
		14531 => to_unsigned(32251, LUT_AMPL_WIDTH - 1),
		14532 => to_unsigned(32252, LUT_AMPL_WIDTH - 1),
		14533 => to_unsigned(32252, LUT_AMPL_WIDTH - 1),
		14534 => to_unsigned(32253, LUT_AMPL_WIDTH - 1),
		14535 => to_unsigned(32253, LUT_AMPL_WIDTH - 1),
		14536 => to_unsigned(32254, LUT_AMPL_WIDTH - 1),
		14537 => to_unsigned(32255, LUT_AMPL_WIDTH - 1),
		14538 => to_unsigned(32255, LUT_AMPL_WIDTH - 1),
		14539 => to_unsigned(32256, LUT_AMPL_WIDTH - 1),
		14540 => to_unsigned(32256, LUT_AMPL_WIDTH - 1),
		14541 => to_unsigned(32257, LUT_AMPL_WIDTH - 1),
		14542 => to_unsigned(32257, LUT_AMPL_WIDTH - 1),
		14543 => to_unsigned(32258, LUT_AMPL_WIDTH - 1),
		14544 => to_unsigned(32258, LUT_AMPL_WIDTH - 1),
		14545 => to_unsigned(32259, LUT_AMPL_WIDTH - 1),
		14546 => to_unsigned(32260, LUT_AMPL_WIDTH - 1),
		14547 => to_unsigned(32260, LUT_AMPL_WIDTH - 1),
		14548 => to_unsigned(32261, LUT_AMPL_WIDTH - 1),
		14549 => to_unsigned(32261, LUT_AMPL_WIDTH - 1),
		14550 => to_unsigned(32262, LUT_AMPL_WIDTH - 1),
		14551 => to_unsigned(32262, LUT_AMPL_WIDTH - 1),
		14552 => to_unsigned(32263, LUT_AMPL_WIDTH - 1),
		14553 => to_unsigned(32263, LUT_AMPL_WIDTH - 1),
		14554 => to_unsigned(32264, LUT_AMPL_WIDTH - 1),
		14555 => to_unsigned(32265, LUT_AMPL_WIDTH - 1),
		14556 => to_unsigned(32265, LUT_AMPL_WIDTH - 1),
		14557 => to_unsigned(32266, LUT_AMPL_WIDTH - 1),
		14558 => to_unsigned(32266, LUT_AMPL_WIDTH - 1),
		14559 => to_unsigned(32267, LUT_AMPL_WIDTH - 1),
		14560 => to_unsigned(32267, LUT_AMPL_WIDTH - 1),
		14561 => to_unsigned(32268, LUT_AMPL_WIDTH - 1),
		14562 => to_unsigned(32268, LUT_AMPL_WIDTH - 1),
		14563 => to_unsigned(32269, LUT_AMPL_WIDTH - 1),
		14564 => to_unsigned(32269, LUT_AMPL_WIDTH - 1),
		14565 => to_unsigned(32270, LUT_AMPL_WIDTH - 1),
		14566 => to_unsigned(32271, LUT_AMPL_WIDTH - 1),
		14567 => to_unsigned(32271, LUT_AMPL_WIDTH - 1),
		14568 => to_unsigned(32272, LUT_AMPL_WIDTH - 1),
		14569 => to_unsigned(32272, LUT_AMPL_WIDTH - 1),
		14570 => to_unsigned(32273, LUT_AMPL_WIDTH - 1),
		14571 => to_unsigned(32273, LUT_AMPL_WIDTH - 1),
		14572 => to_unsigned(32274, LUT_AMPL_WIDTH - 1),
		14573 => to_unsigned(32274, LUT_AMPL_WIDTH - 1),
		14574 => to_unsigned(32275, LUT_AMPL_WIDTH - 1),
		14575 => to_unsigned(32275, LUT_AMPL_WIDTH - 1),
		14576 => to_unsigned(32276, LUT_AMPL_WIDTH - 1),
		14577 => to_unsigned(32277, LUT_AMPL_WIDTH - 1),
		14578 => to_unsigned(32277, LUT_AMPL_WIDTH - 1),
		14579 => to_unsigned(32278, LUT_AMPL_WIDTH - 1),
		14580 => to_unsigned(32278, LUT_AMPL_WIDTH - 1),
		14581 => to_unsigned(32279, LUT_AMPL_WIDTH - 1),
		14582 => to_unsigned(32279, LUT_AMPL_WIDTH - 1),
		14583 => to_unsigned(32280, LUT_AMPL_WIDTH - 1),
		14584 => to_unsigned(32280, LUT_AMPL_WIDTH - 1),
		14585 => to_unsigned(32281, LUT_AMPL_WIDTH - 1),
		14586 => to_unsigned(32281, LUT_AMPL_WIDTH - 1),
		14587 => to_unsigned(32282, LUT_AMPL_WIDTH - 1),
		14588 => to_unsigned(32282, LUT_AMPL_WIDTH - 1),
		14589 => to_unsigned(32283, LUT_AMPL_WIDTH - 1),
		14590 => to_unsigned(32284, LUT_AMPL_WIDTH - 1),
		14591 => to_unsigned(32284, LUT_AMPL_WIDTH - 1),
		14592 => to_unsigned(32285, LUT_AMPL_WIDTH - 1),
		14593 => to_unsigned(32285, LUT_AMPL_WIDTH - 1),
		14594 => to_unsigned(32286, LUT_AMPL_WIDTH - 1),
		14595 => to_unsigned(32286, LUT_AMPL_WIDTH - 1),
		14596 => to_unsigned(32287, LUT_AMPL_WIDTH - 1),
		14597 => to_unsigned(32287, LUT_AMPL_WIDTH - 1),
		14598 => to_unsigned(32288, LUT_AMPL_WIDTH - 1),
		14599 => to_unsigned(32288, LUT_AMPL_WIDTH - 1),
		14600 => to_unsigned(32289, LUT_AMPL_WIDTH - 1),
		14601 => to_unsigned(32289, LUT_AMPL_WIDTH - 1),
		14602 => to_unsigned(32290, LUT_AMPL_WIDTH - 1),
		14603 => to_unsigned(32290, LUT_AMPL_WIDTH - 1),
		14604 => to_unsigned(32291, LUT_AMPL_WIDTH - 1),
		14605 => to_unsigned(32292, LUT_AMPL_WIDTH - 1),
		14606 => to_unsigned(32292, LUT_AMPL_WIDTH - 1),
		14607 => to_unsigned(32293, LUT_AMPL_WIDTH - 1),
		14608 => to_unsigned(32293, LUT_AMPL_WIDTH - 1),
		14609 => to_unsigned(32294, LUT_AMPL_WIDTH - 1),
		14610 => to_unsigned(32294, LUT_AMPL_WIDTH - 1),
		14611 => to_unsigned(32295, LUT_AMPL_WIDTH - 1),
		14612 => to_unsigned(32295, LUT_AMPL_WIDTH - 1),
		14613 => to_unsigned(32296, LUT_AMPL_WIDTH - 1),
		14614 => to_unsigned(32296, LUT_AMPL_WIDTH - 1),
		14615 => to_unsigned(32297, LUT_AMPL_WIDTH - 1),
		14616 => to_unsigned(32297, LUT_AMPL_WIDTH - 1),
		14617 => to_unsigned(32298, LUT_AMPL_WIDTH - 1),
		14618 => to_unsigned(32298, LUT_AMPL_WIDTH - 1),
		14619 => to_unsigned(32299, LUT_AMPL_WIDTH - 1),
		14620 => to_unsigned(32300, LUT_AMPL_WIDTH - 1),
		14621 => to_unsigned(32300, LUT_AMPL_WIDTH - 1),
		14622 => to_unsigned(32301, LUT_AMPL_WIDTH - 1),
		14623 => to_unsigned(32301, LUT_AMPL_WIDTH - 1),
		14624 => to_unsigned(32302, LUT_AMPL_WIDTH - 1),
		14625 => to_unsigned(32302, LUT_AMPL_WIDTH - 1),
		14626 => to_unsigned(32303, LUT_AMPL_WIDTH - 1),
		14627 => to_unsigned(32303, LUT_AMPL_WIDTH - 1),
		14628 => to_unsigned(32304, LUT_AMPL_WIDTH - 1),
		14629 => to_unsigned(32304, LUT_AMPL_WIDTH - 1),
		14630 => to_unsigned(32305, LUT_AMPL_WIDTH - 1),
		14631 => to_unsigned(32305, LUT_AMPL_WIDTH - 1),
		14632 => to_unsigned(32306, LUT_AMPL_WIDTH - 1),
		14633 => to_unsigned(32306, LUT_AMPL_WIDTH - 1),
		14634 => to_unsigned(32307, LUT_AMPL_WIDTH - 1),
		14635 => to_unsigned(32307, LUT_AMPL_WIDTH - 1),
		14636 => to_unsigned(32308, LUT_AMPL_WIDTH - 1),
		14637 => to_unsigned(32308, LUT_AMPL_WIDTH - 1),
		14638 => to_unsigned(32309, LUT_AMPL_WIDTH - 1),
		14639 => to_unsigned(32310, LUT_AMPL_WIDTH - 1),
		14640 => to_unsigned(32310, LUT_AMPL_WIDTH - 1),
		14641 => to_unsigned(32311, LUT_AMPL_WIDTH - 1),
		14642 => to_unsigned(32311, LUT_AMPL_WIDTH - 1),
		14643 => to_unsigned(32312, LUT_AMPL_WIDTH - 1),
		14644 => to_unsigned(32312, LUT_AMPL_WIDTH - 1),
		14645 => to_unsigned(32313, LUT_AMPL_WIDTH - 1),
		14646 => to_unsigned(32313, LUT_AMPL_WIDTH - 1),
		14647 => to_unsigned(32314, LUT_AMPL_WIDTH - 1),
		14648 => to_unsigned(32314, LUT_AMPL_WIDTH - 1),
		14649 => to_unsigned(32315, LUT_AMPL_WIDTH - 1),
		14650 => to_unsigned(32315, LUT_AMPL_WIDTH - 1),
		14651 => to_unsigned(32316, LUT_AMPL_WIDTH - 1),
		14652 => to_unsigned(32316, LUT_AMPL_WIDTH - 1),
		14653 => to_unsigned(32317, LUT_AMPL_WIDTH - 1),
		14654 => to_unsigned(32317, LUT_AMPL_WIDTH - 1),
		14655 => to_unsigned(32318, LUT_AMPL_WIDTH - 1),
		14656 => to_unsigned(32318, LUT_AMPL_WIDTH - 1),
		14657 => to_unsigned(32319, LUT_AMPL_WIDTH - 1),
		14658 => to_unsigned(32319, LUT_AMPL_WIDTH - 1),
		14659 => to_unsigned(32320, LUT_AMPL_WIDTH - 1),
		14660 => to_unsigned(32320, LUT_AMPL_WIDTH - 1),
		14661 => to_unsigned(32321, LUT_AMPL_WIDTH - 1),
		14662 => to_unsigned(32321, LUT_AMPL_WIDTH - 1),
		14663 => to_unsigned(32322, LUT_AMPL_WIDTH - 1),
		14664 => to_unsigned(32322, LUT_AMPL_WIDTH - 1),
		14665 => to_unsigned(32323, LUT_AMPL_WIDTH - 1),
		14666 => to_unsigned(32324, LUT_AMPL_WIDTH - 1),
		14667 => to_unsigned(32324, LUT_AMPL_WIDTH - 1),
		14668 => to_unsigned(32325, LUT_AMPL_WIDTH - 1),
		14669 => to_unsigned(32325, LUT_AMPL_WIDTH - 1),
		14670 => to_unsigned(32326, LUT_AMPL_WIDTH - 1),
		14671 => to_unsigned(32326, LUT_AMPL_WIDTH - 1),
		14672 => to_unsigned(32327, LUT_AMPL_WIDTH - 1),
		14673 => to_unsigned(32327, LUT_AMPL_WIDTH - 1),
		14674 => to_unsigned(32328, LUT_AMPL_WIDTH - 1),
		14675 => to_unsigned(32328, LUT_AMPL_WIDTH - 1),
		14676 => to_unsigned(32329, LUT_AMPL_WIDTH - 1),
		14677 => to_unsigned(32329, LUT_AMPL_WIDTH - 1),
		14678 => to_unsigned(32330, LUT_AMPL_WIDTH - 1),
		14679 => to_unsigned(32330, LUT_AMPL_WIDTH - 1),
		14680 => to_unsigned(32331, LUT_AMPL_WIDTH - 1),
		14681 => to_unsigned(32331, LUT_AMPL_WIDTH - 1),
		14682 => to_unsigned(32332, LUT_AMPL_WIDTH - 1),
		14683 => to_unsigned(32332, LUT_AMPL_WIDTH - 1),
		14684 => to_unsigned(32333, LUT_AMPL_WIDTH - 1),
		14685 => to_unsigned(32333, LUT_AMPL_WIDTH - 1),
		14686 => to_unsigned(32334, LUT_AMPL_WIDTH - 1),
		14687 => to_unsigned(32334, LUT_AMPL_WIDTH - 1),
		14688 => to_unsigned(32335, LUT_AMPL_WIDTH - 1),
		14689 => to_unsigned(32335, LUT_AMPL_WIDTH - 1),
		14690 => to_unsigned(32336, LUT_AMPL_WIDTH - 1),
		14691 => to_unsigned(32336, LUT_AMPL_WIDTH - 1),
		14692 => to_unsigned(32337, LUT_AMPL_WIDTH - 1),
		14693 => to_unsigned(32337, LUT_AMPL_WIDTH - 1),
		14694 => to_unsigned(32338, LUT_AMPL_WIDTH - 1),
		14695 => to_unsigned(32338, LUT_AMPL_WIDTH - 1),
		14696 => to_unsigned(32339, LUT_AMPL_WIDTH - 1),
		14697 => to_unsigned(32339, LUT_AMPL_WIDTH - 1),
		14698 => to_unsigned(32340, LUT_AMPL_WIDTH - 1),
		14699 => to_unsigned(32340, LUT_AMPL_WIDTH - 1),
		14700 => to_unsigned(32341, LUT_AMPL_WIDTH - 1),
		14701 => to_unsigned(32341, LUT_AMPL_WIDTH - 1),
		14702 => to_unsigned(32342, LUT_AMPL_WIDTH - 1),
		14703 => to_unsigned(32342, LUT_AMPL_WIDTH - 1),
		14704 => to_unsigned(32343, LUT_AMPL_WIDTH - 1),
		14705 => to_unsigned(32343, LUT_AMPL_WIDTH - 1),
		14706 => to_unsigned(32344, LUT_AMPL_WIDTH - 1),
		14707 => to_unsigned(32344, LUT_AMPL_WIDTH - 1),
		14708 => to_unsigned(32345, LUT_AMPL_WIDTH - 1),
		14709 => to_unsigned(32345, LUT_AMPL_WIDTH - 1),
		14710 => to_unsigned(32346, LUT_AMPL_WIDTH - 1),
		14711 => to_unsigned(32346, LUT_AMPL_WIDTH - 1),
		14712 => to_unsigned(32347, LUT_AMPL_WIDTH - 1),
		14713 => to_unsigned(32347, LUT_AMPL_WIDTH - 1),
		14714 => to_unsigned(32348, LUT_AMPL_WIDTH - 1),
		14715 => to_unsigned(32348, LUT_AMPL_WIDTH - 1),
		14716 => to_unsigned(32349, LUT_AMPL_WIDTH - 1),
		14717 => to_unsigned(32349, LUT_AMPL_WIDTH - 1),
		14718 => to_unsigned(32350, LUT_AMPL_WIDTH - 1),
		14719 => to_unsigned(32350, LUT_AMPL_WIDTH - 1),
		14720 => to_unsigned(32351, LUT_AMPL_WIDTH - 1),
		14721 => to_unsigned(32351, LUT_AMPL_WIDTH - 1),
		14722 => to_unsigned(32352, LUT_AMPL_WIDTH - 1),
		14723 => to_unsigned(32352, LUT_AMPL_WIDTH - 1),
		14724 => to_unsigned(32353, LUT_AMPL_WIDTH - 1),
		14725 => to_unsigned(32353, LUT_AMPL_WIDTH - 1),
		14726 => to_unsigned(32354, LUT_AMPL_WIDTH - 1),
		14727 => to_unsigned(32354, LUT_AMPL_WIDTH - 1),
		14728 => to_unsigned(32355, LUT_AMPL_WIDTH - 1),
		14729 => to_unsigned(32355, LUT_AMPL_WIDTH - 1),
		14730 => to_unsigned(32356, LUT_AMPL_WIDTH - 1),
		14731 => to_unsigned(32356, LUT_AMPL_WIDTH - 1),
		14732 => to_unsigned(32357, LUT_AMPL_WIDTH - 1),
		14733 => to_unsigned(32357, LUT_AMPL_WIDTH - 1),
		14734 => to_unsigned(32358, LUT_AMPL_WIDTH - 1),
		14735 => to_unsigned(32358, LUT_AMPL_WIDTH - 1),
		14736 => to_unsigned(32359, LUT_AMPL_WIDTH - 1),
		14737 => to_unsigned(32359, LUT_AMPL_WIDTH - 1),
		14738 => to_unsigned(32360, LUT_AMPL_WIDTH - 1),
		14739 => to_unsigned(32360, LUT_AMPL_WIDTH - 1),
		14740 => to_unsigned(32361, LUT_AMPL_WIDTH - 1),
		14741 => to_unsigned(32361, LUT_AMPL_WIDTH - 1),
		14742 => to_unsigned(32362, LUT_AMPL_WIDTH - 1),
		14743 => to_unsigned(32362, LUT_AMPL_WIDTH - 1),
		14744 => to_unsigned(32363, LUT_AMPL_WIDTH - 1),
		14745 => to_unsigned(32363, LUT_AMPL_WIDTH - 1),
		14746 => to_unsigned(32364, LUT_AMPL_WIDTH - 1),
		14747 => to_unsigned(32364, LUT_AMPL_WIDTH - 1),
		14748 => to_unsigned(32365, LUT_AMPL_WIDTH - 1),
		14749 => to_unsigned(32365, LUT_AMPL_WIDTH - 1),
		14750 => to_unsigned(32366, LUT_AMPL_WIDTH - 1),
		14751 => to_unsigned(32366, LUT_AMPL_WIDTH - 1),
		14752 => to_unsigned(32367, LUT_AMPL_WIDTH - 1),
		14753 => to_unsigned(32367, LUT_AMPL_WIDTH - 1),
		14754 => to_unsigned(32368, LUT_AMPL_WIDTH - 1),
		14755 => to_unsigned(32368, LUT_AMPL_WIDTH - 1),
		14756 => to_unsigned(32369, LUT_AMPL_WIDTH - 1),
		14757 => to_unsigned(32369, LUT_AMPL_WIDTH - 1),
		14758 => to_unsigned(32370, LUT_AMPL_WIDTH - 1),
		14759 => to_unsigned(32370, LUT_AMPL_WIDTH - 1),
		14760 => to_unsigned(32371, LUT_AMPL_WIDTH - 1),
		14761 => to_unsigned(32371, LUT_AMPL_WIDTH - 1),
		14762 => to_unsigned(32372, LUT_AMPL_WIDTH - 1),
		14763 => to_unsigned(32372, LUT_AMPL_WIDTH - 1),
		14764 => to_unsigned(32373, LUT_AMPL_WIDTH - 1),
		14765 => to_unsigned(32373, LUT_AMPL_WIDTH - 1),
		14766 => to_unsigned(32374, LUT_AMPL_WIDTH - 1),
		14767 => to_unsigned(32374, LUT_AMPL_WIDTH - 1),
		14768 => to_unsigned(32375, LUT_AMPL_WIDTH - 1),
		14769 => to_unsigned(32375, LUT_AMPL_WIDTH - 1),
		14770 => to_unsigned(32375, LUT_AMPL_WIDTH - 1),
		14771 => to_unsigned(32376, LUT_AMPL_WIDTH - 1),
		14772 => to_unsigned(32376, LUT_AMPL_WIDTH - 1),
		14773 => to_unsigned(32377, LUT_AMPL_WIDTH - 1),
		14774 => to_unsigned(32377, LUT_AMPL_WIDTH - 1),
		14775 => to_unsigned(32378, LUT_AMPL_WIDTH - 1),
		14776 => to_unsigned(32378, LUT_AMPL_WIDTH - 1),
		14777 => to_unsigned(32379, LUT_AMPL_WIDTH - 1),
		14778 => to_unsigned(32379, LUT_AMPL_WIDTH - 1),
		14779 => to_unsigned(32380, LUT_AMPL_WIDTH - 1),
		14780 => to_unsigned(32380, LUT_AMPL_WIDTH - 1),
		14781 => to_unsigned(32381, LUT_AMPL_WIDTH - 1),
		14782 => to_unsigned(32381, LUT_AMPL_WIDTH - 1),
		14783 => to_unsigned(32382, LUT_AMPL_WIDTH - 1),
		14784 => to_unsigned(32382, LUT_AMPL_WIDTH - 1),
		14785 => to_unsigned(32383, LUT_AMPL_WIDTH - 1),
		14786 => to_unsigned(32383, LUT_AMPL_WIDTH - 1),
		14787 => to_unsigned(32384, LUT_AMPL_WIDTH - 1),
		14788 => to_unsigned(32384, LUT_AMPL_WIDTH - 1),
		14789 => to_unsigned(32385, LUT_AMPL_WIDTH - 1),
		14790 => to_unsigned(32385, LUT_AMPL_WIDTH - 1),
		14791 => to_unsigned(32386, LUT_AMPL_WIDTH - 1),
		14792 => to_unsigned(32386, LUT_AMPL_WIDTH - 1),
		14793 => to_unsigned(32387, LUT_AMPL_WIDTH - 1),
		14794 => to_unsigned(32387, LUT_AMPL_WIDTH - 1),
		14795 => to_unsigned(32387, LUT_AMPL_WIDTH - 1),
		14796 => to_unsigned(32388, LUT_AMPL_WIDTH - 1),
		14797 => to_unsigned(32388, LUT_AMPL_WIDTH - 1),
		14798 => to_unsigned(32389, LUT_AMPL_WIDTH - 1),
		14799 => to_unsigned(32389, LUT_AMPL_WIDTH - 1),
		14800 => to_unsigned(32390, LUT_AMPL_WIDTH - 1),
		14801 => to_unsigned(32390, LUT_AMPL_WIDTH - 1),
		14802 => to_unsigned(32391, LUT_AMPL_WIDTH - 1),
		14803 => to_unsigned(32391, LUT_AMPL_WIDTH - 1),
		14804 => to_unsigned(32392, LUT_AMPL_WIDTH - 1),
		14805 => to_unsigned(32392, LUT_AMPL_WIDTH - 1),
		14806 => to_unsigned(32393, LUT_AMPL_WIDTH - 1),
		14807 => to_unsigned(32393, LUT_AMPL_WIDTH - 1),
		14808 => to_unsigned(32394, LUT_AMPL_WIDTH - 1),
		14809 => to_unsigned(32394, LUT_AMPL_WIDTH - 1),
		14810 => to_unsigned(32395, LUT_AMPL_WIDTH - 1),
		14811 => to_unsigned(32395, LUT_AMPL_WIDTH - 1),
		14812 => to_unsigned(32396, LUT_AMPL_WIDTH - 1),
		14813 => to_unsigned(32396, LUT_AMPL_WIDTH - 1),
		14814 => to_unsigned(32397, LUT_AMPL_WIDTH - 1),
		14815 => to_unsigned(32397, LUT_AMPL_WIDTH - 1),
		14816 => to_unsigned(32397, LUT_AMPL_WIDTH - 1),
		14817 => to_unsigned(32398, LUT_AMPL_WIDTH - 1),
		14818 => to_unsigned(32398, LUT_AMPL_WIDTH - 1),
		14819 => to_unsigned(32399, LUT_AMPL_WIDTH - 1),
		14820 => to_unsigned(32399, LUT_AMPL_WIDTH - 1),
		14821 => to_unsigned(32400, LUT_AMPL_WIDTH - 1),
		14822 => to_unsigned(32400, LUT_AMPL_WIDTH - 1),
		14823 => to_unsigned(32401, LUT_AMPL_WIDTH - 1),
		14824 => to_unsigned(32401, LUT_AMPL_WIDTH - 1),
		14825 => to_unsigned(32402, LUT_AMPL_WIDTH - 1),
		14826 => to_unsigned(32402, LUT_AMPL_WIDTH - 1),
		14827 => to_unsigned(32403, LUT_AMPL_WIDTH - 1),
		14828 => to_unsigned(32403, LUT_AMPL_WIDTH - 1),
		14829 => to_unsigned(32404, LUT_AMPL_WIDTH - 1),
		14830 => to_unsigned(32404, LUT_AMPL_WIDTH - 1),
		14831 => to_unsigned(32404, LUT_AMPL_WIDTH - 1),
		14832 => to_unsigned(32405, LUT_AMPL_WIDTH - 1),
		14833 => to_unsigned(32405, LUT_AMPL_WIDTH - 1),
		14834 => to_unsigned(32406, LUT_AMPL_WIDTH - 1),
		14835 => to_unsigned(32406, LUT_AMPL_WIDTH - 1),
		14836 => to_unsigned(32407, LUT_AMPL_WIDTH - 1),
		14837 => to_unsigned(32407, LUT_AMPL_WIDTH - 1),
		14838 => to_unsigned(32408, LUT_AMPL_WIDTH - 1),
		14839 => to_unsigned(32408, LUT_AMPL_WIDTH - 1),
		14840 => to_unsigned(32409, LUT_AMPL_WIDTH - 1),
		14841 => to_unsigned(32409, LUT_AMPL_WIDTH - 1),
		14842 => to_unsigned(32410, LUT_AMPL_WIDTH - 1),
		14843 => to_unsigned(32410, LUT_AMPL_WIDTH - 1),
		14844 => to_unsigned(32411, LUT_AMPL_WIDTH - 1),
		14845 => to_unsigned(32411, LUT_AMPL_WIDTH - 1),
		14846 => to_unsigned(32411, LUT_AMPL_WIDTH - 1),
		14847 => to_unsigned(32412, LUT_AMPL_WIDTH - 1),
		14848 => to_unsigned(32412, LUT_AMPL_WIDTH - 1),
		14849 => to_unsigned(32413, LUT_AMPL_WIDTH - 1),
		14850 => to_unsigned(32413, LUT_AMPL_WIDTH - 1),
		14851 => to_unsigned(32414, LUT_AMPL_WIDTH - 1),
		14852 => to_unsigned(32414, LUT_AMPL_WIDTH - 1),
		14853 => to_unsigned(32415, LUT_AMPL_WIDTH - 1),
		14854 => to_unsigned(32415, LUT_AMPL_WIDTH - 1),
		14855 => to_unsigned(32416, LUT_AMPL_WIDTH - 1),
		14856 => to_unsigned(32416, LUT_AMPL_WIDTH - 1),
		14857 => to_unsigned(32416, LUT_AMPL_WIDTH - 1),
		14858 => to_unsigned(32417, LUT_AMPL_WIDTH - 1),
		14859 => to_unsigned(32417, LUT_AMPL_WIDTH - 1),
		14860 => to_unsigned(32418, LUT_AMPL_WIDTH - 1),
		14861 => to_unsigned(32418, LUT_AMPL_WIDTH - 1),
		14862 => to_unsigned(32419, LUT_AMPL_WIDTH - 1),
		14863 => to_unsigned(32419, LUT_AMPL_WIDTH - 1),
		14864 => to_unsigned(32420, LUT_AMPL_WIDTH - 1),
		14865 => to_unsigned(32420, LUT_AMPL_WIDTH - 1),
		14866 => to_unsigned(32421, LUT_AMPL_WIDTH - 1),
		14867 => to_unsigned(32421, LUT_AMPL_WIDTH - 1),
		14868 => to_unsigned(32422, LUT_AMPL_WIDTH - 1),
		14869 => to_unsigned(32422, LUT_AMPL_WIDTH - 1),
		14870 => to_unsigned(32422, LUT_AMPL_WIDTH - 1),
		14871 => to_unsigned(32423, LUT_AMPL_WIDTH - 1),
		14872 => to_unsigned(32423, LUT_AMPL_WIDTH - 1),
		14873 => to_unsigned(32424, LUT_AMPL_WIDTH - 1),
		14874 => to_unsigned(32424, LUT_AMPL_WIDTH - 1),
		14875 => to_unsigned(32425, LUT_AMPL_WIDTH - 1),
		14876 => to_unsigned(32425, LUT_AMPL_WIDTH - 1),
		14877 => to_unsigned(32426, LUT_AMPL_WIDTH - 1),
		14878 => to_unsigned(32426, LUT_AMPL_WIDTH - 1),
		14879 => to_unsigned(32426, LUT_AMPL_WIDTH - 1),
		14880 => to_unsigned(32427, LUT_AMPL_WIDTH - 1),
		14881 => to_unsigned(32427, LUT_AMPL_WIDTH - 1),
		14882 => to_unsigned(32428, LUT_AMPL_WIDTH - 1),
		14883 => to_unsigned(32428, LUT_AMPL_WIDTH - 1),
		14884 => to_unsigned(32429, LUT_AMPL_WIDTH - 1),
		14885 => to_unsigned(32429, LUT_AMPL_WIDTH - 1),
		14886 => to_unsigned(32430, LUT_AMPL_WIDTH - 1),
		14887 => to_unsigned(32430, LUT_AMPL_WIDTH - 1),
		14888 => to_unsigned(32431, LUT_AMPL_WIDTH - 1),
		14889 => to_unsigned(32431, LUT_AMPL_WIDTH - 1),
		14890 => to_unsigned(32431, LUT_AMPL_WIDTH - 1),
		14891 => to_unsigned(32432, LUT_AMPL_WIDTH - 1),
		14892 => to_unsigned(32432, LUT_AMPL_WIDTH - 1),
		14893 => to_unsigned(32433, LUT_AMPL_WIDTH - 1),
		14894 => to_unsigned(32433, LUT_AMPL_WIDTH - 1),
		14895 => to_unsigned(32434, LUT_AMPL_WIDTH - 1),
		14896 => to_unsigned(32434, LUT_AMPL_WIDTH - 1),
		14897 => to_unsigned(32435, LUT_AMPL_WIDTH - 1),
		14898 => to_unsigned(32435, LUT_AMPL_WIDTH - 1),
		14899 => to_unsigned(32435, LUT_AMPL_WIDTH - 1),
		14900 => to_unsigned(32436, LUT_AMPL_WIDTH - 1),
		14901 => to_unsigned(32436, LUT_AMPL_WIDTH - 1),
		14902 => to_unsigned(32437, LUT_AMPL_WIDTH - 1),
		14903 => to_unsigned(32437, LUT_AMPL_WIDTH - 1),
		14904 => to_unsigned(32438, LUT_AMPL_WIDTH - 1),
		14905 => to_unsigned(32438, LUT_AMPL_WIDTH - 1),
		14906 => to_unsigned(32439, LUT_AMPL_WIDTH - 1),
		14907 => to_unsigned(32439, LUT_AMPL_WIDTH - 1),
		14908 => to_unsigned(32439, LUT_AMPL_WIDTH - 1),
		14909 => to_unsigned(32440, LUT_AMPL_WIDTH - 1),
		14910 => to_unsigned(32440, LUT_AMPL_WIDTH - 1),
		14911 => to_unsigned(32441, LUT_AMPL_WIDTH - 1),
		14912 => to_unsigned(32441, LUT_AMPL_WIDTH - 1),
		14913 => to_unsigned(32442, LUT_AMPL_WIDTH - 1),
		14914 => to_unsigned(32442, LUT_AMPL_WIDTH - 1),
		14915 => to_unsigned(32443, LUT_AMPL_WIDTH - 1),
		14916 => to_unsigned(32443, LUT_AMPL_WIDTH - 1),
		14917 => to_unsigned(32443, LUT_AMPL_WIDTH - 1),
		14918 => to_unsigned(32444, LUT_AMPL_WIDTH - 1),
		14919 => to_unsigned(32444, LUT_AMPL_WIDTH - 1),
		14920 => to_unsigned(32445, LUT_AMPL_WIDTH - 1),
		14921 => to_unsigned(32445, LUT_AMPL_WIDTH - 1),
		14922 => to_unsigned(32446, LUT_AMPL_WIDTH - 1),
		14923 => to_unsigned(32446, LUT_AMPL_WIDTH - 1),
		14924 => to_unsigned(32447, LUT_AMPL_WIDTH - 1),
		14925 => to_unsigned(32447, LUT_AMPL_WIDTH - 1),
		14926 => to_unsigned(32447, LUT_AMPL_WIDTH - 1),
		14927 => to_unsigned(32448, LUT_AMPL_WIDTH - 1),
		14928 => to_unsigned(32448, LUT_AMPL_WIDTH - 1),
		14929 => to_unsigned(32449, LUT_AMPL_WIDTH - 1),
		14930 => to_unsigned(32449, LUT_AMPL_WIDTH - 1),
		14931 => to_unsigned(32450, LUT_AMPL_WIDTH - 1),
		14932 => to_unsigned(32450, LUT_AMPL_WIDTH - 1),
		14933 => to_unsigned(32450, LUT_AMPL_WIDTH - 1),
		14934 => to_unsigned(32451, LUT_AMPL_WIDTH - 1),
		14935 => to_unsigned(32451, LUT_AMPL_WIDTH - 1),
		14936 => to_unsigned(32452, LUT_AMPL_WIDTH - 1),
		14937 => to_unsigned(32452, LUT_AMPL_WIDTH - 1),
		14938 => to_unsigned(32453, LUT_AMPL_WIDTH - 1),
		14939 => to_unsigned(32453, LUT_AMPL_WIDTH - 1),
		14940 => to_unsigned(32453, LUT_AMPL_WIDTH - 1),
		14941 => to_unsigned(32454, LUT_AMPL_WIDTH - 1),
		14942 => to_unsigned(32454, LUT_AMPL_WIDTH - 1),
		14943 => to_unsigned(32455, LUT_AMPL_WIDTH - 1),
		14944 => to_unsigned(32455, LUT_AMPL_WIDTH - 1),
		14945 => to_unsigned(32456, LUT_AMPL_WIDTH - 1),
		14946 => to_unsigned(32456, LUT_AMPL_WIDTH - 1),
		14947 => to_unsigned(32457, LUT_AMPL_WIDTH - 1),
		14948 => to_unsigned(32457, LUT_AMPL_WIDTH - 1),
		14949 => to_unsigned(32457, LUT_AMPL_WIDTH - 1),
		14950 => to_unsigned(32458, LUT_AMPL_WIDTH - 1),
		14951 => to_unsigned(32458, LUT_AMPL_WIDTH - 1),
		14952 => to_unsigned(32459, LUT_AMPL_WIDTH - 1),
		14953 => to_unsigned(32459, LUT_AMPL_WIDTH - 1),
		14954 => to_unsigned(32460, LUT_AMPL_WIDTH - 1),
		14955 => to_unsigned(32460, LUT_AMPL_WIDTH - 1),
		14956 => to_unsigned(32460, LUT_AMPL_WIDTH - 1),
		14957 => to_unsigned(32461, LUT_AMPL_WIDTH - 1),
		14958 => to_unsigned(32461, LUT_AMPL_WIDTH - 1),
		14959 => to_unsigned(32462, LUT_AMPL_WIDTH - 1),
		14960 => to_unsigned(32462, LUT_AMPL_WIDTH - 1),
		14961 => to_unsigned(32463, LUT_AMPL_WIDTH - 1),
		14962 => to_unsigned(32463, LUT_AMPL_WIDTH - 1),
		14963 => to_unsigned(32463, LUT_AMPL_WIDTH - 1),
		14964 => to_unsigned(32464, LUT_AMPL_WIDTH - 1),
		14965 => to_unsigned(32464, LUT_AMPL_WIDTH - 1),
		14966 => to_unsigned(32465, LUT_AMPL_WIDTH - 1),
		14967 => to_unsigned(32465, LUT_AMPL_WIDTH - 1),
		14968 => to_unsigned(32466, LUT_AMPL_WIDTH - 1),
		14969 => to_unsigned(32466, LUT_AMPL_WIDTH - 1),
		14970 => to_unsigned(32466, LUT_AMPL_WIDTH - 1),
		14971 => to_unsigned(32467, LUT_AMPL_WIDTH - 1),
		14972 => to_unsigned(32467, LUT_AMPL_WIDTH - 1),
		14973 => to_unsigned(32468, LUT_AMPL_WIDTH - 1),
		14974 => to_unsigned(32468, LUT_AMPL_WIDTH - 1),
		14975 => to_unsigned(32468, LUT_AMPL_WIDTH - 1),
		14976 => to_unsigned(32469, LUT_AMPL_WIDTH - 1),
		14977 => to_unsigned(32469, LUT_AMPL_WIDTH - 1),
		14978 => to_unsigned(32470, LUT_AMPL_WIDTH - 1),
		14979 => to_unsigned(32470, LUT_AMPL_WIDTH - 1),
		14980 => to_unsigned(32471, LUT_AMPL_WIDTH - 1),
		14981 => to_unsigned(32471, LUT_AMPL_WIDTH - 1),
		14982 => to_unsigned(32471, LUT_AMPL_WIDTH - 1),
		14983 => to_unsigned(32472, LUT_AMPL_WIDTH - 1),
		14984 => to_unsigned(32472, LUT_AMPL_WIDTH - 1),
		14985 => to_unsigned(32473, LUT_AMPL_WIDTH - 1),
		14986 => to_unsigned(32473, LUT_AMPL_WIDTH - 1),
		14987 => to_unsigned(32474, LUT_AMPL_WIDTH - 1),
		14988 => to_unsigned(32474, LUT_AMPL_WIDTH - 1),
		14989 => to_unsigned(32474, LUT_AMPL_WIDTH - 1),
		14990 => to_unsigned(32475, LUT_AMPL_WIDTH - 1),
		14991 => to_unsigned(32475, LUT_AMPL_WIDTH - 1),
		14992 => to_unsigned(32476, LUT_AMPL_WIDTH - 1),
		14993 => to_unsigned(32476, LUT_AMPL_WIDTH - 1),
		14994 => to_unsigned(32476, LUT_AMPL_WIDTH - 1),
		14995 => to_unsigned(32477, LUT_AMPL_WIDTH - 1),
		14996 => to_unsigned(32477, LUT_AMPL_WIDTH - 1),
		14997 => to_unsigned(32478, LUT_AMPL_WIDTH - 1),
		14998 => to_unsigned(32478, LUT_AMPL_WIDTH - 1),
		14999 => to_unsigned(32479, LUT_AMPL_WIDTH - 1),
		15000 => to_unsigned(32479, LUT_AMPL_WIDTH - 1),
		15001 => to_unsigned(32479, LUT_AMPL_WIDTH - 1),
		15002 => to_unsigned(32480, LUT_AMPL_WIDTH - 1),
		15003 => to_unsigned(32480, LUT_AMPL_WIDTH - 1),
		15004 => to_unsigned(32481, LUT_AMPL_WIDTH - 1),
		15005 => to_unsigned(32481, LUT_AMPL_WIDTH - 1),
		15006 => to_unsigned(32481, LUT_AMPL_WIDTH - 1),
		15007 => to_unsigned(32482, LUT_AMPL_WIDTH - 1),
		15008 => to_unsigned(32482, LUT_AMPL_WIDTH - 1),
		15009 => to_unsigned(32483, LUT_AMPL_WIDTH - 1),
		15010 => to_unsigned(32483, LUT_AMPL_WIDTH - 1),
		15011 => to_unsigned(32484, LUT_AMPL_WIDTH - 1),
		15012 => to_unsigned(32484, LUT_AMPL_WIDTH - 1),
		15013 => to_unsigned(32484, LUT_AMPL_WIDTH - 1),
		15014 => to_unsigned(32485, LUT_AMPL_WIDTH - 1),
		15015 => to_unsigned(32485, LUT_AMPL_WIDTH - 1),
		15016 => to_unsigned(32486, LUT_AMPL_WIDTH - 1),
		15017 => to_unsigned(32486, LUT_AMPL_WIDTH - 1),
		15018 => to_unsigned(32486, LUT_AMPL_WIDTH - 1),
		15019 => to_unsigned(32487, LUT_AMPL_WIDTH - 1),
		15020 => to_unsigned(32487, LUT_AMPL_WIDTH - 1),
		15021 => to_unsigned(32488, LUT_AMPL_WIDTH - 1),
		15022 => to_unsigned(32488, LUT_AMPL_WIDTH - 1),
		15023 => to_unsigned(32488, LUT_AMPL_WIDTH - 1),
		15024 => to_unsigned(32489, LUT_AMPL_WIDTH - 1),
		15025 => to_unsigned(32489, LUT_AMPL_WIDTH - 1),
		15026 => to_unsigned(32490, LUT_AMPL_WIDTH - 1),
		15027 => to_unsigned(32490, LUT_AMPL_WIDTH - 1),
		15028 => to_unsigned(32490, LUT_AMPL_WIDTH - 1),
		15029 => to_unsigned(32491, LUT_AMPL_WIDTH - 1),
		15030 => to_unsigned(32491, LUT_AMPL_WIDTH - 1),
		15031 => to_unsigned(32492, LUT_AMPL_WIDTH - 1),
		15032 => to_unsigned(32492, LUT_AMPL_WIDTH - 1),
		15033 => to_unsigned(32493, LUT_AMPL_WIDTH - 1),
		15034 => to_unsigned(32493, LUT_AMPL_WIDTH - 1),
		15035 => to_unsigned(32493, LUT_AMPL_WIDTH - 1),
		15036 => to_unsigned(32494, LUT_AMPL_WIDTH - 1),
		15037 => to_unsigned(32494, LUT_AMPL_WIDTH - 1),
		15038 => to_unsigned(32495, LUT_AMPL_WIDTH - 1),
		15039 => to_unsigned(32495, LUT_AMPL_WIDTH - 1),
		15040 => to_unsigned(32495, LUT_AMPL_WIDTH - 1),
		15041 => to_unsigned(32496, LUT_AMPL_WIDTH - 1),
		15042 => to_unsigned(32496, LUT_AMPL_WIDTH - 1),
		15043 => to_unsigned(32497, LUT_AMPL_WIDTH - 1),
		15044 => to_unsigned(32497, LUT_AMPL_WIDTH - 1),
		15045 => to_unsigned(32497, LUT_AMPL_WIDTH - 1),
		15046 => to_unsigned(32498, LUT_AMPL_WIDTH - 1),
		15047 => to_unsigned(32498, LUT_AMPL_WIDTH - 1),
		15048 => to_unsigned(32499, LUT_AMPL_WIDTH - 1),
		15049 => to_unsigned(32499, LUT_AMPL_WIDTH - 1),
		15050 => to_unsigned(32499, LUT_AMPL_WIDTH - 1),
		15051 => to_unsigned(32500, LUT_AMPL_WIDTH - 1),
		15052 => to_unsigned(32500, LUT_AMPL_WIDTH - 1),
		15053 => to_unsigned(32501, LUT_AMPL_WIDTH - 1),
		15054 => to_unsigned(32501, LUT_AMPL_WIDTH - 1),
		15055 => to_unsigned(32501, LUT_AMPL_WIDTH - 1),
		15056 => to_unsigned(32502, LUT_AMPL_WIDTH - 1),
		15057 => to_unsigned(32502, LUT_AMPL_WIDTH - 1),
		15058 => to_unsigned(32503, LUT_AMPL_WIDTH - 1),
		15059 => to_unsigned(32503, LUT_AMPL_WIDTH - 1),
		15060 => to_unsigned(32503, LUT_AMPL_WIDTH - 1),
		15061 => to_unsigned(32504, LUT_AMPL_WIDTH - 1),
		15062 => to_unsigned(32504, LUT_AMPL_WIDTH - 1),
		15063 => to_unsigned(32505, LUT_AMPL_WIDTH - 1),
		15064 => to_unsigned(32505, LUT_AMPL_WIDTH - 1),
		15065 => to_unsigned(32505, LUT_AMPL_WIDTH - 1),
		15066 => to_unsigned(32506, LUT_AMPL_WIDTH - 1),
		15067 => to_unsigned(32506, LUT_AMPL_WIDTH - 1),
		15068 => to_unsigned(32507, LUT_AMPL_WIDTH - 1),
		15069 => to_unsigned(32507, LUT_AMPL_WIDTH - 1),
		15070 => to_unsigned(32507, LUT_AMPL_WIDTH - 1),
		15071 => to_unsigned(32508, LUT_AMPL_WIDTH - 1),
		15072 => to_unsigned(32508, LUT_AMPL_WIDTH - 1),
		15073 => to_unsigned(32509, LUT_AMPL_WIDTH - 1),
		15074 => to_unsigned(32509, LUT_AMPL_WIDTH - 1),
		15075 => to_unsigned(32509, LUT_AMPL_WIDTH - 1),
		15076 => to_unsigned(32510, LUT_AMPL_WIDTH - 1),
		15077 => to_unsigned(32510, LUT_AMPL_WIDTH - 1),
		15078 => to_unsigned(32510, LUT_AMPL_WIDTH - 1),
		15079 => to_unsigned(32511, LUT_AMPL_WIDTH - 1),
		15080 => to_unsigned(32511, LUT_AMPL_WIDTH - 1),
		15081 => to_unsigned(32512, LUT_AMPL_WIDTH - 1),
		15082 => to_unsigned(32512, LUT_AMPL_WIDTH - 1),
		15083 => to_unsigned(32512, LUT_AMPL_WIDTH - 1),
		15084 => to_unsigned(32513, LUT_AMPL_WIDTH - 1),
		15085 => to_unsigned(32513, LUT_AMPL_WIDTH - 1),
		15086 => to_unsigned(32514, LUT_AMPL_WIDTH - 1),
		15087 => to_unsigned(32514, LUT_AMPL_WIDTH - 1),
		15088 => to_unsigned(32514, LUT_AMPL_WIDTH - 1),
		15089 => to_unsigned(32515, LUT_AMPL_WIDTH - 1),
		15090 => to_unsigned(32515, LUT_AMPL_WIDTH - 1),
		15091 => to_unsigned(32516, LUT_AMPL_WIDTH - 1),
		15092 => to_unsigned(32516, LUT_AMPL_WIDTH - 1),
		15093 => to_unsigned(32516, LUT_AMPL_WIDTH - 1),
		15094 => to_unsigned(32517, LUT_AMPL_WIDTH - 1),
		15095 => to_unsigned(32517, LUT_AMPL_WIDTH - 1),
		15096 => to_unsigned(32517, LUT_AMPL_WIDTH - 1),
		15097 => to_unsigned(32518, LUT_AMPL_WIDTH - 1),
		15098 => to_unsigned(32518, LUT_AMPL_WIDTH - 1),
		15099 => to_unsigned(32519, LUT_AMPL_WIDTH - 1),
		15100 => to_unsigned(32519, LUT_AMPL_WIDTH - 1),
		15101 => to_unsigned(32519, LUT_AMPL_WIDTH - 1),
		15102 => to_unsigned(32520, LUT_AMPL_WIDTH - 1),
		15103 => to_unsigned(32520, LUT_AMPL_WIDTH - 1),
		15104 => to_unsigned(32521, LUT_AMPL_WIDTH - 1),
		15105 => to_unsigned(32521, LUT_AMPL_WIDTH - 1),
		15106 => to_unsigned(32521, LUT_AMPL_WIDTH - 1),
		15107 => to_unsigned(32522, LUT_AMPL_WIDTH - 1),
		15108 => to_unsigned(32522, LUT_AMPL_WIDTH - 1),
		15109 => to_unsigned(32522, LUT_AMPL_WIDTH - 1),
		15110 => to_unsigned(32523, LUT_AMPL_WIDTH - 1),
		15111 => to_unsigned(32523, LUT_AMPL_WIDTH - 1),
		15112 => to_unsigned(32524, LUT_AMPL_WIDTH - 1),
		15113 => to_unsigned(32524, LUT_AMPL_WIDTH - 1),
		15114 => to_unsigned(32524, LUT_AMPL_WIDTH - 1),
		15115 => to_unsigned(32525, LUT_AMPL_WIDTH - 1),
		15116 => to_unsigned(32525, LUT_AMPL_WIDTH - 1),
		15117 => to_unsigned(32526, LUT_AMPL_WIDTH - 1),
		15118 => to_unsigned(32526, LUT_AMPL_WIDTH - 1),
		15119 => to_unsigned(32526, LUT_AMPL_WIDTH - 1),
		15120 => to_unsigned(32527, LUT_AMPL_WIDTH - 1),
		15121 => to_unsigned(32527, LUT_AMPL_WIDTH - 1),
		15122 => to_unsigned(32527, LUT_AMPL_WIDTH - 1),
		15123 => to_unsigned(32528, LUT_AMPL_WIDTH - 1),
		15124 => to_unsigned(32528, LUT_AMPL_WIDTH - 1),
		15125 => to_unsigned(32529, LUT_AMPL_WIDTH - 1),
		15126 => to_unsigned(32529, LUT_AMPL_WIDTH - 1),
		15127 => to_unsigned(32529, LUT_AMPL_WIDTH - 1),
		15128 => to_unsigned(32530, LUT_AMPL_WIDTH - 1),
		15129 => to_unsigned(32530, LUT_AMPL_WIDTH - 1),
		15130 => to_unsigned(32530, LUT_AMPL_WIDTH - 1),
		15131 => to_unsigned(32531, LUT_AMPL_WIDTH - 1),
		15132 => to_unsigned(32531, LUT_AMPL_WIDTH - 1),
		15133 => to_unsigned(32532, LUT_AMPL_WIDTH - 1),
		15134 => to_unsigned(32532, LUT_AMPL_WIDTH - 1),
		15135 => to_unsigned(32532, LUT_AMPL_WIDTH - 1),
		15136 => to_unsigned(32533, LUT_AMPL_WIDTH - 1),
		15137 => to_unsigned(32533, LUT_AMPL_WIDTH - 1),
		15138 => to_unsigned(32533, LUT_AMPL_WIDTH - 1),
		15139 => to_unsigned(32534, LUT_AMPL_WIDTH - 1),
		15140 => to_unsigned(32534, LUT_AMPL_WIDTH - 1),
		15141 => to_unsigned(32535, LUT_AMPL_WIDTH - 1),
		15142 => to_unsigned(32535, LUT_AMPL_WIDTH - 1),
		15143 => to_unsigned(32535, LUT_AMPL_WIDTH - 1),
		15144 => to_unsigned(32536, LUT_AMPL_WIDTH - 1),
		15145 => to_unsigned(32536, LUT_AMPL_WIDTH - 1),
		15146 => to_unsigned(32536, LUT_AMPL_WIDTH - 1),
		15147 => to_unsigned(32537, LUT_AMPL_WIDTH - 1),
		15148 => to_unsigned(32537, LUT_AMPL_WIDTH - 1),
		15149 => to_unsigned(32538, LUT_AMPL_WIDTH - 1),
		15150 => to_unsigned(32538, LUT_AMPL_WIDTH - 1),
		15151 => to_unsigned(32538, LUT_AMPL_WIDTH - 1),
		15152 => to_unsigned(32539, LUT_AMPL_WIDTH - 1),
		15153 => to_unsigned(32539, LUT_AMPL_WIDTH - 1),
		15154 => to_unsigned(32539, LUT_AMPL_WIDTH - 1),
		15155 => to_unsigned(32540, LUT_AMPL_WIDTH - 1),
		15156 => to_unsigned(32540, LUT_AMPL_WIDTH - 1),
		15157 => to_unsigned(32541, LUT_AMPL_WIDTH - 1),
		15158 => to_unsigned(32541, LUT_AMPL_WIDTH - 1),
		15159 => to_unsigned(32541, LUT_AMPL_WIDTH - 1),
		15160 => to_unsigned(32542, LUT_AMPL_WIDTH - 1),
		15161 => to_unsigned(32542, LUT_AMPL_WIDTH - 1),
		15162 => to_unsigned(32542, LUT_AMPL_WIDTH - 1),
		15163 => to_unsigned(32543, LUT_AMPL_WIDTH - 1),
		15164 => to_unsigned(32543, LUT_AMPL_WIDTH - 1),
		15165 => to_unsigned(32543, LUT_AMPL_WIDTH - 1),
		15166 => to_unsigned(32544, LUT_AMPL_WIDTH - 1),
		15167 => to_unsigned(32544, LUT_AMPL_WIDTH - 1),
		15168 => to_unsigned(32545, LUT_AMPL_WIDTH - 1),
		15169 => to_unsigned(32545, LUT_AMPL_WIDTH - 1),
		15170 => to_unsigned(32545, LUT_AMPL_WIDTH - 1),
		15171 => to_unsigned(32546, LUT_AMPL_WIDTH - 1),
		15172 => to_unsigned(32546, LUT_AMPL_WIDTH - 1),
		15173 => to_unsigned(32546, LUT_AMPL_WIDTH - 1),
		15174 => to_unsigned(32547, LUT_AMPL_WIDTH - 1),
		15175 => to_unsigned(32547, LUT_AMPL_WIDTH - 1),
		15176 => to_unsigned(32547, LUT_AMPL_WIDTH - 1),
		15177 => to_unsigned(32548, LUT_AMPL_WIDTH - 1),
		15178 => to_unsigned(32548, LUT_AMPL_WIDTH - 1),
		15179 => to_unsigned(32549, LUT_AMPL_WIDTH - 1),
		15180 => to_unsigned(32549, LUT_AMPL_WIDTH - 1),
		15181 => to_unsigned(32549, LUT_AMPL_WIDTH - 1),
		15182 => to_unsigned(32550, LUT_AMPL_WIDTH - 1),
		15183 => to_unsigned(32550, LUT_AMPL_WIDTH - 1),
		15184 => to_unsigned(32550, LUT_AMPL_WIDTH - 1),
		15185 => to_unsigned(32551, LUT_AMPL_WIDTH - 1),
		15186 => to_unsigned(32551, LUT_AMPL_WIDTH - 1),
		15187 => to_unsigned(32551, LUT_AMPL_WIDTH - 1),
		15188 => to_unsigned(32552, LUT_AMPL_WIDTH - 1),
		15189 => to_unsigned(32552, LUT_AMPL_WIDTH - 1),
		15190 => to_unsigned(32553, LUT_AMPL_WIDTH - 1),
		15191 => to_unsigned(32553, LUT_AMPL_WIDTH - 1),
		15192 => to_unsigned(32553, LUT_AMPL_WIDTH - 1),
		15193 => to_unsigned(32554, LUT_AMPL_WIDTH - 1),
		15194 => to_unsigned(32554, LUT_AMPL_WIDTH - 1),
		15195 => to_unsigned(32554, LUT_AMPL_WIDTH - 1),
		15196 => to_unsigned(32555, LUT_AMPL_WIDTH - 1),
		15197 => to_unsigned(32555, LUT_AMPL_WIDTH - 1),
		15198 => to_unsigned(32555, LUT_AMPL_WIDTH - 1),
		15199 => to_unsigned(32556, LUT_AMPL_WIDTH - 1),
		15200 => to_unsigned(32556, LUT_AMPL_WIDTH - 1),
		15201 => to_unsigned(32556, LUT_AMPL_WIDTH - 1),
		15202 => to_unsigned(32557, LUT_AMPL_WIDTH - 1),
		15203 => to_unsigned(32557, LUT_AMPL_WIDTH - 1),
		15204 => to_unsigned(32558, LUT_AMPL_WIDTH - 1),
		15205 => to_unsigned(32558, LUT_AMPL_WIDTH - 1),
		15206 => to_unsigned(32558, LUT_AMPL_WIDTH - 1),
		15207 => to_unsigned(32559, LUT_AMPL_WIDTH - 1),
		15208 => to_unsigned(32559, LUT_AMPL_WIDTH - 1),
		15209 => to_unsigned(32559, LUT_AMPL_WIDTH - 1),
		15210 => to_unsigned(32560, LUT_AMPL_WIDTH - 1),
		15211 => to_unsigned(32560, LUT_AMPL_WIDTH - 1),
		15212 => to_unsigned(32560, LUT_AMPL_WIDTH - 1),
		15213 => to_unsigned(32561, LUT_AMPL_WIDTH - 1),
		15214 => to_unsigned(32561, LUT_AMPL_WIDTH - 1),
		15215 => to_unsigned(32561, LUT_AMPL_WIDTH - 1),
		15216 => to_unsigned(32562, LUT_AMPL_WIDTH - 1),
		15217 => to_unsigned(32562, LUT_AMPL_WIDTH - 1),
		15218 => to_unsigned(32562, LUT_AMPL_WIDTH - 1),
		15219 => to_unsigned(32563, LUT_AMPL_WIDTH - 1),
		15220 => to_unsigned(32563, LUT_AMPL_WIDTH - 1),
		15221 => to_unsigned(32564, LUT_AMPL_WIDTH - 1),
		15222 => to_unsigned(32564, LUT_AMPL_WIDTH - 1),
		15223 => to_unsigned(32564, LUT_AMPL_WIDTH - 1),
		15224 => to_unsigned(32565, LUT_AMPL_WIDTH - 1),
		15225 => to_unsigned(32565, LUT_AMPL_WIDTH - 1),
		15226 => to_unsigned(32565, LUT_AMPL_WIDTH - 1),
		15227 => to_unsigned(32566, LUT_AMPL_WIDTH - 1),
		15228 => to_unsigned(32566, LUT_AMPL_WIDTH - 1),
		15229 => to_unsigned(32566, LUT_AMPL_WIDTH - 1),
		15230 => to_unsigned(32567, LUT_AMPL_WIDTH - 1),
		15231 => to_unsigned(32567, LUT_AMPL_WIDTH - 1),
		15232 => to_unsigned(32567, LUT_AMPL_WIDTH - 1),
		15233 => to_unsigned(32568, LUT_AMPL_WIDTH - 1),
		15234 => to_unsigned(32568, LUT_AMPL_WIDTH - 1),
		15235 => to_unsigned(32568, LUT_AMPL_WIDTH - 1),
		15236 => to_unsigned(32569, LUT_AMPL_WIDTH - 1),
		15237 => to_unsigned(32569, LUT_AMPL_WIDTH - 1),
		15238 => to_unsigned(32569, LUT_AMPL_WIDTH - 1),
		15239 => to_unsigned(32570, LUT_AMPL_WIDTH - 1),
		15240 => to_unsigned(32570, LUT_AMPL_WIDTH - 1),
		15241 => to_unsigned(32570, LUT_AMPL_WIDTH - 1),
		15242 => to_unsigned(32571, LUT_AMPL_WIDTH - 1),
		15243 => to_unsigned(32571, LUT_AMPL_WIDTH - 1),
		15244 => to_unsigned(32571, LUT_AMPL_WIDTH - 1),
		15245 => to_unsigned(32572, LUT_AMPL_WIDTH - 1),
		15246 => to_unsigned(32572, LUT_AMPL_WIDTH - 1),
		15247 => to_unsigned(32573, LUT_AMPL_WIDTH - 1),
		15248 => to_unsigned(32573, LUT_AMPL_WIDTH - 1),
		15249 => to_unsigned(32573, LUT_AMPL_WIDTH - 1),
		15250 => to_unsigned(32574, LUT_AMPL_WIDTH - 1),
		15251 => to_unsigned(32574, LUT_AMPL_WIDTH - 1),
		15252 => to_unsigned(32574, LUT_AMPL_WIDTH - 1),
		15253 => to_unsigned(32575, LUT_AMPL_WIDTH - 1),
		15254 => to_unsigned(32575, LUT_AMPL_WIDTH - 1),
		15255 => to_unsigned(32575, LUT_AMPL_WIDTH - 1),
		15256 => to_unsigned(32576, LUT_AMPL_WIDTH - 1),
		15257 => to_unsigned(32576, LUT_AMPL_WIDTH - 1),
		15258 => to_unsigned(32576, LUT_AMPL_WIDTH - 1),
		15259 => to_unsigned(32577, LUT_AMPL_WIDTH - 1),
		15260 => to_unsigned(32577, LUT_AMPL_WIDTH - 1),
		15261 => to_unsigned(32577, LUT_AMPL_WIDTH - 1),
		15262 => to_unsigned(32578, LUT_AMPL_WIDTH - 1),
		15263 => to_unsigned(32578, LUT_AMPL_WIDTH - 1),
		15264 => to_unsigned(32578, LUT_AMPL_WIDTH - 1),
		15265 => to_unsigned(32579, LUT_AMPL_WIDTH - 1),
		15266 => to_unsigned(32579, LUT_AMPL_WIDTH - 1),
		15267 => to_unsigned(32579, LUT_AMPL_WIDTH - 1),
		15268 => to_unsigned(32580, LUT_AMPL_WIDTH - 1),
		15269 => to_unsigned(32580, LUT_AMPL_WIDTH - 1),
		15270 => to_unsigned(32580, LUT_AMPL_WIDTH - 1),
		15271 => to_unsigned(32581, LUT_AMPL_WIDTH - 1),
		15272 => to_unsigned(32581, LUT_AMPL_WIDTH - 1),
		15273 => to_unsigned(32581, LUT_AMPL_WIDTH - 1),
		15274 => to_unsigned(32582, LUT_AMPL_WIDTH - 1),
		15275 => to_unsigned(32582, LUT_AMPL_WIDTH - 1),
		15276 => to_unsigned(32582, LUT_AMPL_WIDTH - 1),
		15277 => to_unsigned(32583, LUT_AMPL_WIDTH - 1),
		15278 => to_unsigned(32583, LUT_AMPL_WIDTH - 1),
		15279 => to_unsigned(32583, LUT_AMPL_WIDTH - 1),
		15280 => to_unsigned(32584, LUT_AMPL_WIDTH - 1),
		15281 => to_unsigned(32584, LUT_AMPL_WIDTH - 1),
		15282 => to_unsigned(32584, LUT_AMPL_WIDTH - 1),
		15283 => to_unsigned(32585, LUT_AMPL_WIDTH - 1),
		15284 => to_unsigned(32585, LUT_AMPL_WIDTH - 1),
		15285 => to_unsigned(32585, LUT_AMPL_WIDTH - 1),
		15286 => to_unsigned(32586, LUT_AMPL_WIDTH - 1),
		15287 => to_unsigned(32586, LUT_AMPL_WIDTH - 1),
		15288 => to_unsigned(32586, LUT_AMPL_WIDTH - 1),
		15289 => to_unsigned(32587, LUT_AMPL_WIDTH - 1),
		15290 => to_unsigned(32587, LUT_AMPL_WIDTH - 1),
		15291 => to_unsigned(32587, LUT_AMPL_WIDTH - 1),
		15292 => to_unsigned(32588, LUT_AMPL_WIDTH - 1),
		15293 => to_unsigned(32588, LUT_AMPL_WIDTH - 1),
		15294 => to_unsigned(32588, LUT_AMPL_WIDTH - 1),
		15295 => to_unsigned(32589, LUT_AMPL_WIDTH - 1),
		15296 => to_unsigned(32589, LUT_AMPL_WIDTH - 1),
		15297 => to_unsigned(32589, LUT_AMPL_WIDTH - 1),
		15298 => to_unsigned(32590, LUT_AMPL_WIDTH - 1),
		15299 => to_unsigned(32590, LUT_AMPL_WIDTH - 1),
		15300 => to_unsigned(32590, LUT_AMPL_WIDTH - 1),
		15301 => to_unsigned(32591, LUT_AMPL_WIDTH - 1),
		15302 => to_unsigned(32591, LUT_AMPL_WIDTH - 1),
		15303 => to_unsigned(32591, LUT_AMPL_WIDTH - 1),
		15304 => to_unsigned(32592, LUT_AMPL_WIDTH - 1),
		15305 => to_unsigned(32592, LUT_AMPL_WIDTH - 1),
		15306 => to_unsigned(32592, LUT_AMPL_WIDTH - 1),
		15307 => to_unsigned(32592, LUT_AMPL_WIDTH - 1),
		15308 => to_unsigned(32593, LUT_AMPL_WIDTH - 1),
		15309 => to_unsigned(32593, LUT_AMPL_WIDTH - 1),
		15310 => to_unsigned(32593, LUT_AMPL_WIDTH - 1),
		15311 => to_unsigned(32594, LUT_AMPL_WIDTH - 1),
		15312 => to_unsigned(32594, LUT_AMPL_WIDTH - 1),
		15313 => to_unsigned(32594, LUT_AMPL_WIDTH - 1),
		15314 => to_unsigned(32595, LUT_AMPL_WIDTH - 1),
		15315 => to_unsigned(32595, LUT_AMPL_WIDTH - 1),
		15316 => to_unsigned(32595, LUT_AMPL_WIDTH - 1),
		15317 => to_unsigned(32596, LUT_AMPL_WIDTH - 1),
		15318 => to_unsigned(32596, LUT_AMPL_WIDTH - 1),
		15319 => to_unsigned(32596, LUT_AMPL_WIDTH - 1),
		15320 => to_unsigned(32597, LUT_AMPL_WIDTH - 1),
		15321 => to_unsigned(32597, LUT_AMPL_WIDTH - 1),
		15322 => to_unsigned(32597, LUT_AMPL_WIDTH - 1),
		15323 => to_unsigned(32598, LUT_AMPL_WIDTH - 1),
		15324 => to_unsigned(32598, LUT_AMPL_WIDTH - 1),
		15325 => to_unsigned(32598, LUT_AMPL_WIDTH - 1),
		15326 => to_unsigned(32599, LUT_AMPL_WIDTH - 1),
		15327 => to_unsigned(32599, LUT_AMPL_WIDTH - 1),
		15328 => to_unsigned(32599, LUT_AMPL_WIDTH - 1),
		15329 => to_unsigned(32600, LUT_AMPL_WIDTH - 1),
		15330 => to_unsigned(32600, LUT_AMPL_WIDTH - 1),
		15331 => to_unsigned(32600, LUT_AMPL_WIDTH - 1),
		15332 => to_unsigned(32600, LUT_AMPL_WIDTH - 1),
		15333 => to_unsigned(32601, LUT_AMPL_WIDTH - 1),
		15334 => to_unsigned(32601, LUT_AMPL_WIDTH - 1),
		15335 => to_unsigned(32601, LUT_AMPL_WIDTH - 1),
		15336 => to_unsigned(32602, LUT_AMPL_WIDTH - 1),
		15337 => to_unsigned(32602, LUT_AMPL_WIDTH - 1),
		15338 => to_unsigned(32602, LUT_AMPL_WIDTH - 1),
		15339 => to_unsigned(32603, LUT_AMPL_WIDTH - 1),
		15340 => to_unsigned(32603, LUT_AMPL_WIDTH - 1),
		15341 => to_unsigned(32603, LUT_AMPL_WIDTH - 1),
		15342 => to_unsigned(32604, LUT_AMPL_WIDTH - 1),
		15343 => to_unsigned(32604, LUT_AMPL_WIDTH - 1),
		15344 => to_unsigned(32604, LUT_AMPL_WIDTH - 1),
		15345 => to_unsigned(32605, LUT_AMPL_WIDTH - 1),
		15346 => to_unsigned(32605, LUT_AMPL_WIDTH - 1),
		15347 => to_unsigned(32605, LUT_AMPL_WIDTH - 1),
		15348 => to_unsigned(32606, LUT_AMPL_WIDTH - 1),
		15349 => to_unsigned(32606, LUT_AMPL_WIDTH - 1),
		15350 => to_unsigned(32606, LUT_AMPL_WIDTH - 1),
		15351 => to_unsigned(32606, LUT_AMPL_WIDTH - 1),
		15352 => to_unsigned(32607, LUT_AMPL_WIDTH - 1),
		15353 => to_unsigned(32607, LUT_AMPL_WIDTH - 1),
		15354 => to_unsigned(32607, LUT_AMPL_WIDTH - 1),
		15355 => to_unsigned(32608, LUT_AMPL_WIDTH - 1),
		15356 => to_unsigned(32608, LUT_AMPL_WIDTH - 1),
		15357 => to_unsigned(32608, LUT_AMPL_WIDTH - 1),
		15358 => to_unsigned(32609, LUT_AMPL_WIDTH - 1),
		15359 => to_unsigned(32609, LUT_AMPL_WIDTH - 1),
		15360 => to_unsigned(32609, LUT_AMPL_WIDTH - 1),
		15361 => to_unsigned(32610, LUT_AMPL_WIDTH - 1),
		15362 => to_unsigned(32610, LUT_AMPL_WIDTH - 1),
		15363 => to_unsigned(32610, LUT_AMPL_WIDTH - 1),
		15364 => to_unsigned(32610, LUT_AMPL_WIDTH - 1),
		15365 => to_unsigned(32611, LUT_AMPL_WIDTH - 1),
		15366 => to_unsigned(32611, LUT_AMPL_WIDTH - 1),
		15367 => to_unsigned(32611, LUT_AMPL_WIDTH - 1),
		15368 => to_unsigned(32612, LUT_AMPL_WIDTH - 1),
		15369 => to_unsigned(32612, LUT_AMPL_WIDTH - 1),
		15370 => to_unsigned(32612, LUT_AMPL_WIDTH - 1),
		15371 => to_unsigned(32613, LUT_AMPL_WIDTH - 1),
		15372 => to_unsigned(32613, LUT_AMPL_WIDTH - 1),
		15373 => to_unsigned(32613, LUT_AMPL_WIDTH - 1),
		15374 => to_unsigned(32613, LUT_AMPL_WIDTH - 1),
		15375 => to_unsigned(32614, LUT_AMPL_WIDTH - 1),
		15376 => to_unsigned(32614, LUT_AMPL_WIDTH - 1),
		15377 => to_unsigned(32614, LUT_AMPL_WIDTH - 1),
		15378 => to_unsigned(32615, LUT_AMPL_WIDTH - 1),
		15379 => to_unsigned(32615, LUT_AMPL_WIDTH - 1),
		15380 => to_unsigned(32615, LUT_AMPL_WIDTH - 1),
		15381 => to_unsigned(32616, LUT_AMPL_WIDTH - 1),
		15382 => to_unsigned(32616, LUT_AMPL_WIDTH - 1),
		15383 => to_unsigned(32616, LUT_AMPL_WIDTH - 1),
		15384 => to_unsigned(32617, LUT_AMPL_WIDTH - 1),
		15385 => to_unsigned(32617, LUT_AMPL_WIDTH - 1),
		15386 => to_unsigned(32617, LUT_AMPL_WIDTH - 1),
		15387 => to_unsigned(32617, LUT_AMPL_WIDTH - 1),
		15388 => to_unsigned(32618, LUT_AMPL_WIDTH - 1),
		15389 => to_unsigned(32618, LUT_AMPL_WIDTH - 1),
		15390 => to_unsigned(32618, LUT_AMPL_WIDTH - 1),
		15391 => to_unsigned(32619, LUT_AMPL_WIDTH - 1),
		15392 => to_unsigned(32619, LUT_AMPL_WIDTH - 1),
		15393 => to_unsigned(32619, LUT_AMPL_WIDTH - 1),
		15394 => to_unsigned(32620, LUT_AMPL_WIDTH - 1),
		15395 => to_unsigned(32620, LUT_AMPL_WIDTH - 1),
		15396 => to_unsigned(32620, LUT_AMPL_WIDTH - 1),
		15397 => to_unsigned(32620, LUT_AMPL_WIDTH - 1),
		15398 => to_unsigned(32621, LUT_AMPL_WIDTH - 1),
		15399 => to_unsigned(32621, LUT_AMPL_WIDTH - 1),
		15400 => to_unsigned(32621, LUT_AMPL_WIDTH - 1),
		15401 => to_unsigned(32622, LUT_AMPL_WIDTH - 1),
		15402 => to_unsigned(32622, LUT_AMPL_WIDTH - 1),
		15403 => to_unsigned(32622, LUT_AMPL_WIDTH - 1),
		15404 => to_unsigned(32622, LUT_AMPL_WIDTH - 1),
		15405 => to_unsigned(32623, LUT_AMPL_WIDTH - 1),
		15406 => to_unsigned(32623, LUT_AMPL_WIDTH - 1),
		15407 => to_unsigned(32623, LUT_AMPL_WIDTH - 1),
		15408 => to_unsigned(32624, LUT_AMPL_WIDTH - 1),
		15409 => to_unsigned(32624, LUT_AMPL_WIDTH - 1),
		15410 => to_unsigned(32624, LUT_AMPL_WIDTH - 1),
		15411 => to_unsigned(32625, LUT_AMPL_WIDTH - 1),
		15412 => to_unsigned(32625, LUT_AMPL_WIDTH - 1),
		15413 => to_unsigned(32625, LUT_AMPL_WIDTH - 1),
		15414 => to_unsigned(32625, LUT_AMPL_WIDTH - 1),
		15415 => to_unsigned(32626, LUT_AMPL_WIDTH - 1),
		15416 => to_unsigned(32626, LUT_AMPL_WIDTH - 1),
		15417 => to_unsigned(32626, LUT_AMPL_WIDTH - 1),
		15418 => to_unsigned(32627, LUT_AMPL_WIDTH - 1),
		15419 => to_unsigned(32627, LUT_AMPL_WIDTH - 1),
		15420 => to_unsigned(32627, LUT_AMPL_WIDTH - 1),
		15421 => to_unsigned(32627, LUT_AMPL_WIDTH - 1),
		15422 => to_unsigned(32628, LUT_AMPL_WIDTH - 1),
		15423 => to_unsigned(32628, LUT_AMPL_WIDTH - 1),
		15424 => to_unsigned(32628, LUT_AMPL_WIDTH - 1),
		15425 => to_unsigned(32629, LUT_AMPL_WIDTH - 1),
		15426 => to_unsigned(32629, LUT_AMPL_WIDTH - 1),
		15427 => to_unsigned(32629, LUT_AMPL_WIDTH - 1),
		15428 => to_unsigned(32629, LUT_AMPL_WIDTH - 1),
		15429 => to_unsigned(32630, LUT_AMPL_WIDTH - 1),
		15430 => to_unsigned(32630, LUT_AMPL_WIDTH - 1),
		15431 => to_unsigned(32630, LUT_AMPL_WIDTH - 1),
		15432 => to_unsigned(32631, LUT_AMPL_WIDTH - 1),
		15433 => to_unsigned(32631, LUT_AMPL_WIDTH - 1),
		15434 => to_unsigned(32631, LUT_AMPL_WIDTH - 1),
		15435 => to_unsigned(32631, LUT_AMPL_WIDTH - 1),
		15436 => to_unsigned(32632, LUT_AMPL_WIDTH - 1),
		15437 => to_unsigned(32632, LUT_AMPL_WIDTH - 1),
		15438 => to_unsigned(32632, LUT_AMPL_WIDTH - 1),
		15439 => to_unsigned(32633, LUT_AMPL_WIDTH - 1),
		15440 => to_unsigned(32633, LUT_AMPL_WIDTH - 1),
		15441 => to_unsigned(32633, LUT_AMPL_WIDTH - 1),
		15442 => to_unsigned(32633, LUT_AMPL_WIDTH - 1),
		15443 => to_unsigned(32634, LUT_AMPL_WIDTH - 1),
		15444 => to_unsigned(32634, LUT_AMPL_WIDTH - 1),
		15445 => to_unsigned(32634, LUT_AMPL_WIDTH - 1),
		15446 => to_unsigned(32635, LUT_AMPL_WIDTH - 1),
		15447 => to_unsigned(32635, LUT_AMPL_WIDTH - 1),
		15448 => to_unsigned(32635, LUT_AMPL_WIDTH - 1),
		15449 => to_unsigned(32635, LUT_AMPL_WIDTH - 1),
		15450 => to_unsigned(32636, LUT_AMPL_WIDTH - 1),
		15451 => to_unsigned(32636, LUT_AMPL_WIDTH - 1),
		15452 => to_unsigned(32636, LUT_AMPL_WIDTH - 1),
		15453 => to_unsigned(32637, LUT_AMPL_WIDTH - 1),
		15454 => to_unsigned(32637, LUT_AMPL_WIDTH - 1),
		15455 => to_unsigned(32637, LUT_AMPL_WIDTH - 1),
		15456 => to_unsigned(32637, LUT_AMPL_WIDTH - 1),
		15457 => to_unsigned(32638, LUT_AMPL_WIDTH - 1),
		15458 => to_unsigned(32638, LUT_AMPL_WIDTH - 1),
		15459 => to_unsigned(32638, LUT_AMPL_WIDTH - 1),
		15460 => to_unsigned(32639, LUT_AMPL_WIDTH - 1),
		15461 => to_unsigned(32639, LUT_AMPL_WIDTH - 1),
		15462 => to_unsigned(32639, LUT_AMPL_WIDTH - 1),
		15463 => to_unsigned(32639, LUT_AMPL_WIDTH - 1),
		15464 => to_unsigned(32640, LUT_AMPL_WIDTH - 1),
		15465 => to_unsigned(32640, LUT_AMPL_WIDTH - 1),
		15466 => to_unsigned(32640, LUT_AMPL_WIDTH - 1),
		15467 => to_unsigned(32640, LUT_AMPL_WIDTH - 1),
		15468 => to_unsigned(32641, LUT_AMPL_WIDTH - 1),
		15469 => to_unsigned(32641, LUT_AMPL_WIDTH - 1),
		15470 => to_unsigned(32641, LUT_AMPL_WIDTH - 1),
		15471 => to_unsigned(32642, LUT_AMPL_WIDTH - 1),
		15472 => to_unsigned(32642, LUT_AMPL_WIDTH - 1),
		15473 => to_unsigned(32642, LUT_AMPL_WIDTH - 1),
		15474 => to_unsigned(32642, LUT_AMPL_WIDTH - 1),
		15475 => to_unsigned(32643, LUT_AMPL_WIDTH - 1),
		15476 => to_unsigned(32643, LUT_AMPL_WIDTH - 1),
		15477 => to_unsigned(32643, LUT_AMPL_WIDTH - 1),
		15478 => to_unsigned(32643, LUT_AMPL_WIDTH - 1),
		15479 => to_unsigned(32644, LUT_AMPL_WIDTH - 1),
		15480 => to_unsigned(32644, LUT_AMPL_WIDTH - 1),
		15481 => to_unsigned(32644, LUT_AMPL_WIDTH - 1),
		15482 => to_unsigned(32645, LUT_AMPL_WIDTH - 1),
		15483 => to_unsigned(32645, LUT_AMPL_WIDTH - 1),
		15484 => to_unsigned(32645, LUT_AMPL_WIDTH - 1),
		15485 => to_unsigned(32645, LUT_AMPL_WIDTH - 1),
		15486 => to_unsigned(32646, LUT_AMPL_WIDTH - 1),
		15487 => to_unsigned(32646, LUT_AMPL_WIDTH - 1),
		15488 => to_unsigned(32646, LUT_AMPL_WIDTH - 1),
		15489 => to_unsigned(32646, LUT_AMPL_WIDTH - 1),
		15490 => to_unsigned(32647, LUT_AMPL_WIDTH - 1),
		15491 => to_unsigned(32647, LUT_AMPL_WIDTH - 1),
		15492 => to_unsigned(32647, LUT_AMPL_WIDTH - 1),
		15493 => to_unsigned(32648, LUT_AMPL_WIDTH - 1),
		15494 => to_unsigned(32648, LUT_AMPL_WIDTH - 1),
		15495 => to_unsigned(32648, LUT_AMPL_WIDTH - 1),
		15496 => to_unsigned(32648, LUT_AMPL_WIDTH - 1),
		15497 => to_unsigned(32649, LUT_AMPL_WIDTH - 1),
		15498 => to_unsigned(32649, LUT_AMPL_WIDTH - 1),
		15499 => to_unsigned(32649, LUT_AMPL_WIDTH - 1),
		15500 => to_unsigned(32649, LUT_AMPL_WIDTH - 1),
		15501 => to_unsigned(32650, LUT_AMPL_WIDTH - 1),
		15502 => to_unsigned(32650, LUT_AMPL_WIDTH - 1),
		15503 => to_unsigned(32650, LUT_AMPL_WIDTH - 1),
		15504 => to_unsigned(32650, LUT_AMPL_WIDTH - 1),
		15505 => to_unsigned(32651, LUT_AMPL_WIDTH - 1),
		15506 => to_unsigned(32651, LUT_AMPL_WIDTH - 1),
		15507 => to_unsigned(32651, LUT_AMPL_WIDTH - 1),
		15508 => to_unsigned(32652, LUT_AMPL_WIDTH - 1),
		15509 => to_unsigned(32652, LUT_AMPL_WIDTH - 1),
		15510 => to_unsigned(32652, LUT_AMPL_WIDTH - 1),
		15511 => to_unsigned(32652, LUT_AMPL_WIDTH - 1),
		15512 => to_unsigned(32653, LUT_AMPL_WIDTH - 1),
		15513 => to_unsigned(32653, LUT_AMPL_WIDTH - 1),
		15514 => to_unsigned(32653, LUT_AMPL_WIDTH - 1),
		15515 => to_unsigned(32653, LUT_AMPL_WIDTH - 1),
		15516 => to_unsigned(32654, LUT_AMPL_WIDTH - 1),
		15517 => to_unsigned(32654, LUT_AMPL_WIDTH - 1),
		15518 => to_unsigned(32654, LUT_AMPL_WIDTH - 1),
		15519 => to_unsigned(32654, LUT_AMPL_WIDTH - 1),
		15520 => to_unsigned(32655, LUT_AMPL_WIDTH - 1),
		15521 => to_unsigned(32655, LUT_AMPL_WIDTH - 1),
		15522 => to_unsigned(32655, LUT_AMPL_WIDTH - 1),
		15523 => to_unsigned(32655, LUT_AMPL_WIDTH - 1),
		15524 => to_unsigned(32656, LUT_AMPL_WIDTH - 1),
		15525 => to_unsigned(32656, LUT_AMPL_WIDTH - 1),
		15526 => to_unsigned(32656, LUT_AMPL_WIDTH - 1),
		15527 => to_unsigned(32656, LUT_AMPL_WIDTH - 1),
		15528 => to_unsigned(32657, LUT_AMPL_WIDTH - 1),
		15529 => to_unsigned(32657, LUT_AMPL_WIDTH - 1),
		15530 => to_unsigned(32657, LUT_AMPL_WIDTH - 1),
		15531 => to_unsigned(32657, LUT_AMPL_WIDTH - 1),
		15532 => to_unsigned(32658, LUT_AMPL_WIDTH - 1),
		15533 => to_unsigned(32658, LUT_AMPL_WIDTH - 1),
		15534 => to_unsigned(32658, LUT_AMPL_WIDTH - 1),
		15535 => to_unsigned(32659, LUT_AMPL_WIDTH - 1),
		15536 => to_unsigned(32659, LUT_AMPL_WIDTH - 1),
		15537 => to_unsigned(32659, LUT_AMPL_WIDTH - 1),
		15538 => to_unsigned(32659, LUT_AMPL_WIDTH - 1),
		15539 => to_unsigned(32660, LUT_AMPL_WIDTH - 1),
		15540 => to_unsigned(32660, LUT_AMPL_WIDTH - 1),
		15541 => to_unsigned(32660, LUT_AMPL_WIDTH - 1),
		15542 => to_unsigned(32660, LUT_AMPL_WIDTH - 1),
		15543 => to_unsigned(32661, LUT_AMPL_WIDTH - 1),
		15544 => to_unsigned(32661, LUT_AMPL_WIDTH - 1),
		15545 => to_unsigned(32661, LUT_AMPL_WIDTH - 1),
		15546 => to_unsigned(32661, LUT_AMPL_WIDTH - 1),
		15547 => to_unsigned(32662, LUT_AMPL_WIDTH - 1),
		15548 => to_unsigned(32662, LUT_AMPL_WIDTH - 1),
		15549 => to_unsigned(32662, LUT_AMPL_WIDTH - 1),
		15550 => to_unsigned(32662, LUT_AMPL_WIDTH - 1),
		15551 => to_unsigned(32663, LUT_AMPL_WIDTH - 1),
		15552 => to_unsigned(32663, LUT_AMPL_WIDTH - 1),
		15553 => to_unsigned(32663, LUT_AMPL_WIDTH - 1),
		15554 => to_unsigned(32663, LUT_AMPL_WIDTH - 1),
		15555 => to_unsigned(32664, LUT_AMPL_WIDTH - 1),
		15556 => to_unsigned(32664, LUT_AMPL_WIDTH - 1),
		15557 => to_unsigned(32664, LUT_AMPL_WIDTH - 1),
		15558 => to_unsigned(32664, LUT_AMPL_WIDTH - 1),
		15559 => to_unsigned(32665, LUT_AMPL_WIDTH - 1),
		15560 => to_unsigned(32665, LUT_AMPL_WIDTH - 1),
		15561 => to_unsigned(32665, LUT_AMPL_WIDTH - 1),
		15562 => to_unsigned(32665, LUT_AMPL_WIDTH - 1),
		15563 => to_unsigned(32666, LUT_AMPL_WIDTH - 1),
		15564 => to_unsigned(32666, LUT_AMPL_WIDTH - 1),
		15565 => to_unsigned(32666, LUT_AMPL_WIDTH - 1),
		15566 => to_unsigned(32666, LUT_AMPL_WIDTH - 1),
		15567 => to_unsigned(32667, LUT_AMPL_WIDTH - 1),
		15568 => to_unsigned(32667, LUT_AMPL_WIDTH - 1),
		15569 => to_unsigned(32667, LUT_AMPL_WIDTH - 1),
		15570 => to_unsigned(32667, LUT_AMPL_WIDTH - 1),
		15571 => to_unsigned(32668, LUT_AMPL_WIDTH - 1),
		15572 => to_unsigned(32668, LUT_AMPL_WIDTH - 1),
		15573 => to_unsigned(32668, LUT_AMPL_WIDTH - 1),
		15574 => to_unsigned(32668, LUT_AMPL_WIDTH - 1),
		15575 => to_unsigned(32668, LUT_AMPL_WIDTH - 1),
		15576 => to_unsigned(32669, LUT_AMPL_WIDTH - 1),
		15577 => to_unsigned(32669, LUT_AMPL_WIDTH - 1),
		15578 => to_unsigned(32669, LUT_AMPL_WIDTH - 1),
		15579 => to_unsigned(32669, LUT_AMPL_WIDTH - 1),
		15580 => to_unsigned(32670, LUT_AMPL_WIDTH - 1),
		15581 => to_unsigned(32670, LUT_AMPL_WIDTH - 1),
		15582 => to_unsigned(32670, LUT_AMPL_WIDTH - 1),
		15583 => to_unsigned(32670, LUT_AMPL_WIDTH - 1),
		15584 => to_unsigned(32671, LUT_AMPL_WIDTH - 1),
		15585 => to_unsigned(32671, LUT_AMPL_WIDTH - 1),
		15586 => to_unsigned(32671, LUT_AMPL_WIDTH - 1),
		15587 => to_unsigned(32671, LUT_AMPL_WIDTH - 1),
		15588 => to_unsigned(32672, LUT_AMPL_WIDTH - 1),
		15589 => to_unsigned(32672, LUT_AMPL_WIDTH - 1),
		15590 => to_unsigned(32672, LUT_AMPL_WIDTH - 1),
		15591 => to_unsigned(32672, LUT_AMPL_WIDTH - 1),
		15592 => to_unsigned(32673, LUT_AMPL_WIDTH - 1),
		15593 => to_unsigned(32673, LUT_AMPL_WIDTH - 1),
		15594 => to_unsigned(32673, LUT_AMPL_WIDTH - 1),
		15595 => to_unsigned(32673, LUT_AMPL_WIDTH - 1),
		15596 => to_unsigned(32674, LUT_AMPL_WIDTH - 1),
		15597 => to_unsigned(32674, LUT_AMPL_WIDTH - 1),
		15598 => to_unsigned(32674, LUT_AMPL_WIDTH - 1),
		15599 => to_unsigned(32674, LUT_AMPL_WIDTH - 1),
		15600 => to_unsigned(32674, LUT_AMPL_WIDTH - 1),
		15601 => to_unsigned(32675, LUT_AMPL_WIDTH - 1),
		15602 => to_unsigned(32675, LUT_AMPL_WIDTH - 1),
		15603 => to_unsigned(32675, LUT_AMPL_WIDTH - 1),
		15604 => to_unsigned(32675, LUT_AMPL_WIDTH - 1),
		15605 => to_unsigned(32676, LUT_AMPL_WIDTH - 1),
		15606 => to_unsigned(32676, LUT_AMPL_WIDTH - 1),
		15607 => to_unsigned(32676, LUT_AMPL_WIDTH - 1),
		15608 => to_unsigned(32676, LUT_AMPL_WIDTH - 1),
		15609 => to_unsigned(32677, LUT_AMPL_WIDTH - 1),
		15610 => to_unsigned(32677, LUT_AMPL_WIDTH - 1),
		15611 => to_unsigned(32677, LUT_AMPL_WIDTH - 1),
		15612 => to_unsigned(32677, LUT_AMPL_WIDTH - 1),
		15613 => to_unsigned(32678, LUT_AMPL_WIDTH - 1),
		15614 => to_unsigned(32678, LUT_AMPL_WIDTH - 1),
		15615 => to_unsigned(32678, LUT_AMPL_WIDTH - 1),
		15616 => to_unsigned(32678, LUT_AMPL_WIDTH - 1),
		15617 => to_unsigned(32678, LUT_AMPL_WIDTH - 1),
		15618 => to_unsigned(32679, LUT_AMPL_WIDTH - 1),
		15619 => to_unsigned(32679, LUT_AMPL_WIDTH - 1),
		15620 => to_unsigned(32679, LUT_AMPL_WIDTH - 1),
		15621 => to_unsigned(32679, LUT_AMPL_WIDTH - 1),
		15622 => to_unsigned(32680, LUT_AMPL_WIDTH - 1),
		15623 => to_unsigned(32680, LUT_AMPL_WIDTH - 1),
		15624 => to_unsigned(32680, LUT_AMPL_WIDTH - 1),
		15625 => to_unsigned(32680, LUT_AMPL_WIDTH - 1),
		15626 => to_unsigned(32681, LUT_AMPL_WIDTH - 1),
		15627 => to_unsigned(32681, LUT_AMPL_WIDTH - 1),
		15628 => to_unsigned(32681, LUT_AMPL_WIDTH - 1),
		15629 => to_unsigned(32681, LUT_AMPL_WIDTH - 1),
		15630 => to_unsigned(32681, LUT_AMPL_WIDTH - 1),
		15631 => to_unsigned(32682, LUT_AMPL_WIDTH - 1),
		15632 => to_unsigned(32682, LUT_AMPL_WIDTH - 1),
		15633 => to_unsigned(32682, LUT_AMPL_WIDTH - 1),
		15634 => to_unsigned(32682, LUT_AMPL_WIDTH - 1),
		15635 => to_unsigned(32683, LUT_AMPL_WIDTH - 1),
		15636 => to_unsigned(32683, LUT_AMPL_WIDTH - 1),
		15637 => to_unsigned(32683, LUT_AMPL_WIDTH - 1),
		15638 => to_unsigned(32683, LUT_AMPL_WIDTH - 1),
		15639 => to_unsigned(32683, LUT_AMPL_WIDTH - 1),
		15640 => to_unsigned(32684, LUT_AMPL_WIDTH - 1),
		15641 => to_unsigned(32684, LUT_AMPL_WIDTH - 1),
		15642 => to_unsigned(32684, LUT_AMPL_WIDTH - 1),
		15643 => to_unsigned(32684, LUT_AMPL_WIDTH - 1),
		15644 => to_unsigned(32685, LUT_AMPL_WIDTH - 1),
		15645 => to_unsigned(32685, LUT_AMPL_WIDTH - 1),
		15646 => to_unsigned(32685, LUT_AMPL_WIDTH - 1),
		15647 => to_unsigned(32685, LUT_AMPL_WIDTH - 1),
		15648 => to_unsigned(32685, LUT_AMPL_WIDTH - 1),
		15649 => to_unsigned(32686, LUT_AMPL_WIDTH - 1),
		15650 => to_unsigned(32686, LUT_AMPL_WIDTH - 1),
		15651 => to_unsigned(32686, LUT_AMPL_WIDTH - 1),
		15652 => to_unsigned(32686, LUT_AMPL_WIDTH - 1),
		15653 => to_unsigned(32687, LUT_AMPL_WIDTH - 1),
		15654 => to_unsigned(32687, LUT_AMPL_WIDTH - 1),
		15655 => to_unsigned(32687, LUT_AMPL_WIDTH - 1),
		15656 => to_unsigned(32687, LUT_AMPL_WIDTH - 1),
		15657 => to_unsigned(32687, LUT_AMPL_WIDTH - 1),
		15658 => to_unsigned(32688, LUT_AMPL_WIDTH - 1),
		15659 => to_unsigned(32688, LUT_AMPL_WIDTH - 1),
		15660 => to_unsigned(32688, LUT_AMPL_WIDTH - 1),
		15661 => to_unsigned(32688, LUT_AMPL_WIDTH - 1),
		15662 => to_unsigned(32689, LUT_AMPL_WIDTH - 1),
		15663 => to_unsigned(32689, LUT_AMPL_WIDTH - 1),
		15664 => to_unsigned(32689, LUT_AMPL_WIDTH - 1),
		15665 => to_unsigned(32689, LUT_AMPL_WIDTH - 1),
		15666 => to_unsigned(32689, LUT_AMPL_WIDTH - 1),
		15667 => to_unsigned(32690, LUT_AMPL_WIDTH - 1),
		15668 => to_unsigned(32690, LUT_AMPL_WIDTH - 1),
		15669 => to_unsigned(32690, LUT_AMPL_WIDTH - 1),
		15670 => to_unsigned(32690, LUT_AMPL_WIDTH - 1),
		15671 => to_unsigned(32690, LUT_AMPL_WIDTH - 1),
		15672 => to_unsigned(32691, LUT_AMPL_WIDTH - 1),
		15673 => to_unsigned(32691, LUT_AMPL_WIDTH - 1),
		15674 => to_unsigned(32691, LUT_AMPL_WIDTH - 1),
		15675 => to_unsigned(32691, LUT_AMPL_WIDTH - 1),
		15676 => to_unsigned(32692, LUT_AMPL_WIDTH - 1),
		15677 => to_unsigned(32692, LUT_AMPL_WIDTH - 1),
		15678 => to_unsigned(32692, LUT_AMPL_WIDTH - 1),
		15679 => to_unsigned(32692, LUT_AMPL_WIDTH - 1),
		15680 => to_unsigned(32692, LUT_AMPL_WIDTH - 1),
		15681 => to_unsigned(32693, LUT_AMPL_WIDTH - 1),
		15682 => to_unsigned(32693, LUT_AMPL_WIDTH - 1),
		15683 => to_unsigned(32693, LUT_AMPL_WIDTH - 1),
		15684 => to_unsigned(32693, LUT_AMPL_WIDTH - 1),
		15685 => to_unsigned(32693, LUT_AMPL_WIDTH - 1),
		15686 => to_unsigned(32694, LUT_AMPL_WIDTH - 1),
		15687 => to_unsigned(32694, LUT_AMPL_WIDTH - 1),
		15688 => to_unsigned(32694, LUT_AMPL_WIDTH - 1),
		15689 => to_unsigned(32694, LUT_AMPL_WIDTH - 1),
		15690 => to_unsigned(32694, LUT_AMPL_WIDTH - 1),
		15691 => to_unsigned(32695, LUT_AMPL_WIDTH - 1),
		15692 => to_unsigned(32695, LUT_AMPL_WIDTH - 1),
		15693 => to_unsigned(32695, LUT_AMPL_WIDTH - 1),
		15694 => to_unsigned(32695, LUT_AMPL_WIDTH - 1),
		15695 => to_unsigned(32696, LUT_AMPL_WIDTH - 1),
		15696 => to_unsigned(32696, LUT_AMPL_WIDTH - 1),
		15697 => to_unsigned(32696, LUT_AMPL_WIDTH - 1),
		15698 => to_unsigned(32696, LUT_AMPL_WIDTH - 1),
		15699 => to_unsigned(32696, LUT_AMPL_WIDTH - 1),
		15700 => to_unsigned(32697, LUT_AMPL_WIDTH - 1),
		15701 => to_unsigned(32697, LUT_AMPL_WIDTH - 1),
		15702 => to_unsigned(32697, LUT_AMPL_WIDTH - 1),
		15703 => to_unsigned(32697, LUT_AMPL_WIDTH - 1),
		15704 => to_unsigned(32697, LUT_AMPL_WIDTH - 1),
		15705 => to_unsigned(32698, LUT_AMPL_WIDTH - 1),
		15706 => to_unsigned(32698, LUT_AMPL_WIDTH - 1),
		15707 => to_unsigned(32698, LUT_AMPL_WIDTH - 1),
		15708 => to_unsigned(32698, LUT_AMPL_WIDTH - 1),
		15709 => to_unsigned(32698, LUT_AMPL_WIDTH - 1),
		15710 => to_unsigned(32699, LUT_AMPL_WIDTH - 1),
		15711 => to_unsigned(32699, LUT_AMPL_WIDTH - 1),
		15712 => to_unsigned(32699, LUT_AMPL_WIDTH - 1),
		15713 => to_unsigned(32699, LUT_AMPL_WIDTH - 1),
		15714 => to_unsigned(32699, LUT_AMPL_WIDTH - 1),
		15715 => to_unsigned(32700, LUT_AMPL_WIDTH - 1),
		15716 => to_unsigned(32700, LUT_AMPL_WIDTH - 1),
		15717 => to_unsigned(32700, LUT_AMPL_WIDTH - 1),
		15718 => to_unsigned(32700, LUT_AMPL_WIDTH - 1),
		15719 => to_unsigned(32700, LUT_AMPL_WIDTH - 1),
		15720 => to_unsigned(32701, LUT_AMPL_WIDTH - 1),
		15721 => to_unsigned(32701, LUT_AMPL_WIDTH - 1),
		15722 => to_unsigned(32701, LUT_AMPL_WIDTH - 1),
		15723 => to_unsigned(32701, LUT_AMPL_WIDTH - 1),
		15724 => to_unsigned(32701, LUT_AMPL_WIDTH - 1),
		15725 => to_unsigned(32702, LUT_AMPL_WIDTH - 1),
		15726 => to_unsigned(32702, LUT_AMPL_WIDTH - 1),
		15727 => to_unsigned(32702, LUT_AMPL_WIDTH - 1),
		15728 => to_unsigned(32702, LUT_AMPL_WIDTH - 1),
		15729 => to_unsigned(32702, LUT_AMPL_WIDTH - 1),
		15730 => to_unsigned(32703, LUT_AMPL_WIDTH - 1),
		15731 => to_unsigned(32703, LUT_AMPL_WIDTH - 1),
		15732 => to_unsigned(32703, LUT_AMPL_WIDTH - 1),
		15733 => to_unsigned(32703, LUT_AMPL_WIDTH - 1),
		15734 => to_unsigned(32703, LUT_AMPL_WIDTH - 1),
		15735 => to_unsigned(32704, LUT_AMPL_WIDTH - 1),
		15736 => to_unsigned(32704, LUT_AMPL_WIDTH - 1),
		15737 => to_unsigned(32704, LUT_AMPL_WIDTH - 1),
		15738 => to_unsigned(32704, LUT_AMPL_WIDTH - 1),
		15739 => to_unsigned(32704, LUT_AMPL_WIDTH - 1),
		15740 => to_unsigned(32705, LUT_AMPL_WIDTH - 1),
		15741 => to_unsigned(32705, LUT_AMPL_WIDTH - 1),
		15742 => to_unsigned(32705, LUT_AMPL_WIDTH - 1),
		15743 => to_unsigned(32705, LUT_AMPL_WIDTH - 1),
		15744 => to_unsigned(32705, LUT_AMPL_WIDTH - 1),
		15745 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		15746 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		15747 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		15748 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		15749 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		15750 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		15751 => to_unsigned(32707, LUT_AMPL_WIDTH - 1),
		15752 => to_unsigned(32707, LUT_AMPL_WIDTH - 1),
		15753 => to_unsigned(32707, LUT_AMPL_WIDTH - 1),
		15754 => to_unsigned(32707, LUT_AMPL_WIDTH - 1),
		15755 => to_unsigned(32707, LUT_AMPL_WIDTH - 1),
		15756 => to_unsigned(32708, LUT_AMPL_WIDTH - 1),
		15757 => to_unsigned(32708, LUT_AMPL_WIDTH - 1),
		15758 => to_unsigned(32708, LUT_AMPL_WIDTH - 1),
		15759 => to_unsigned(32708, LUT_AMPL_WIDTH - 1),
		15760 => to_unsigned(32708, LUT_AMPL_WIDTH - 1),
		15761 => to_unsigned(32709, LUT_AMPL_WIDTH - 1),
		15762 => to_unsigned(32709, LUT_AMPL_WIDTH - 1),
		15763 => to_unsigned(32709, LUT_AMPL_WIDTH - 1),
		15764 => to_unsigned(32709, LUT_AMPL_WIDTH - 1),
		15765 => to_unsigned(32709, LUT_AMPL_WIDTH - 1),
		15766 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		15767 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		15768 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		15769 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		15770 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		15771 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		15772 => to_unsigned(32711, LUT_AMPL_WIDTH - 1),
		15773 => to_unsigned(32711, LUT_AMPL_WIDTH - 1),
		15774 => to_unsigned(32711, LUT_AMPL_WIDTH - 1),
		15775 => to_unsigned(32711, LUT_AMPL_WIDTH - 1),
		15776 => to_unsigned(32711, LUT_AMPL_WIDTH - 1),
		15777 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		15778 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		15779 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		15780 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		15781 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		15782 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		15783 => to_unsigned(32713, LUT_AMPL_WIDTH - 1),
		15784 => to_unsigned(32713, LUT_AMPL_WIDTH - 1),
		15785 => to_unsigned(32713, LUT_AMPL_WIDTH - 1),
		15786 => to_unsigned(32713, LUT_AMPL_WIDTH - 1),
		15787 => to_unsigned(32713, LUT_AMPL_WIDTH - 1),
		15788 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		15789 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		15790 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		15791 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		15792 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		15793 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		15794 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		15795 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		15796 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		15797 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		15798 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		15799 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		15800 => to_unsigned(32716, LUT_AMPL_WIDTH - 1),
		15801 => to_unsigned(32716, LUT_AMPL_WIDTH - 1),
		15802 => to_unsigned(32716, LUT_AMPL_WIDTH - 1),
		15803 => to_unsigned(32716, LUT_AMPL_WIDTH - 1),
		15804 => to_unsigned(32716, LUT_AMPL_WIDTH - 1),
		15805 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		15806 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		15807 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		15808 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		15809 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		15810 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		15811 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		15812 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		15813 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		15814 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		15815 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		15816 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		15817 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		15818 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		15819 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		15820 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		15821 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		15822 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		15823 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		15824 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		15825 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		15826 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		15827 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		15828 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		15829 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		15830 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		15831 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		15832 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		15833 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		15834 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		15835 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		15836 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		15837 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		15838 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		15839 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		15840 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		15841 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		15842 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		15843 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		15844 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		15845 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		15846 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		15847 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		15848 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		15849 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		15850 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		15851 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		15852 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		15853 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		15854 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		15855 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		15856 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		15857 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		15858 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		15859 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		15860 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		15861 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		15862 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		15863 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		15864 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		15865 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		15866 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		15867 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		15868 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		15869 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		15870 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		15871 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		15872 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		15873 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		15874 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		15875 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		15876 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		15877 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		15878 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		15879 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		15880 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		15881 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		15882 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		15883 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		15884 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		15885 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		15886 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		15887 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		15888 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		15889 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		15890 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		15891 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		15892 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		15893 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		15894 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		15895 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		15896 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		15897 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		15898 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		15899 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		15900 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		15901 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		15902 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		15903 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		15904 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		15905 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		15906 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		15907 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		15908 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		15909 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		15910 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		15911 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		15912 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		15913 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		15914 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		15915 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		15916 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		15917 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		15918 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		15919 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		15920 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		15921 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		15922 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		15923 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		15924 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		15925 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		15926 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		15927 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		15928 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		15929 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		15930 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		15931 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		15932 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		15933 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		15934 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		15935 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		15936 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		15937 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		15938 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		15939 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		15940 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		15941 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		15942 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		15943 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		15944 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		15945 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		15946 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		15947 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		15948 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		15949 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		15950 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		15951 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		15952 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		15953 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		15954 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		15955 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		15956 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		15957 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		15958 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		15959 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		15960 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		15961 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		15962 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		15963 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		15964 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		15965 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		15966 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		15967 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		15968 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		15969 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		15970 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		15971 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		15972 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		15973 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		15974 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		15975 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		15976 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		15977 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		15978 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		15979 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		15980 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		15981 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		15982 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		15983 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		15984 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		15985 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		15986 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		15987 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		15988 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		15989 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		15990 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		15991 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		15992 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		15993 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		15994 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		15995 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		15996 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		15997 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		15998 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		15999 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16000 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16001 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16002 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16003 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16004 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16005 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16006 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16007 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16008 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16009 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16010 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16011 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16012 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16013 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16014 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16015 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16016 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16017 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16018 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16019 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16020 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16021 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16022 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16023 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16024 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16025 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16026 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16027 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16028 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16029 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16030 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16031 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16032 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16033 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16034 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16035 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16036 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16037 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16038 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16039 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16040 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16041 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16042 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16043 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16044 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16045 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16046 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16047 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16048 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16049 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16050 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16051 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16052 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16053 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16054 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16055 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16056 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16057 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16058 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16059 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16060 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16061 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16062 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16063 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16064 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16065 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16066 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16067 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16068 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16069 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16070 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16071 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16072 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16073 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16074 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16075 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16076 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16077 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16078 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16079 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16080 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16081 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16082 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16083 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16084 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16085 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16086 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16087 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16088 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16089 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16090 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16091 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16092 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16093 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16094 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16095 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16096 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16097 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16098 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16099 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16100 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16101 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16102 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16103 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16104 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16105 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16106 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16107 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16108 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16109 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16110 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16111 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16112 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16113 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16114 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16115 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16116 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16117 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16118 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16119 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16120 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16121 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16122 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16123 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16124 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16125 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16126 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16127 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16128 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16129 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16130 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16131 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16132 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16133 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16134 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16135 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16136 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16137 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16138 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16139 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16140 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16141 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16142 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16143 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16144 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16145 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16146 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16147 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16148 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16149 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16150 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16151 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16152 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16153 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16154 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16155 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16156 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16157 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16158 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16159 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16160 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16161 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16162 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16163 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16164 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16165 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16166 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16167 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16168 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16169 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16170 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16171 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16172 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16173 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16174 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16175 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16176 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16177 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16178 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16179 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16180 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16181 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16182 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16183 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16184 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16185 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16186 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16187 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16188 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16189 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16190 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16191 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16192 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16193 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16194 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16195 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16196 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16197 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16198 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16199 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16200 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16201 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16202 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16203 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16204 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16205 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16206 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16207 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16208 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16209 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16210 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16211 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16212 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16213 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16214 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16215 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16216 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16217 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16218 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16219 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16220 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16221 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16222 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16223 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16224 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16225 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16226 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16227 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16228 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16229 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16230 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16231 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16232 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16233 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16234 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16235 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16236 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16237 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16238 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16239 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16240 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16241 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16242 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16243 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16244 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16245 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16246 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16247 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16248 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16249 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16250 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16251 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16252 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16253 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16254 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16255 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16256 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16257 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16258 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16259 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16260 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16261 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16262 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16263 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16264 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16265 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16266 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16267 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16268 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16269 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16270 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16271 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16272 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16273 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16274 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16275 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16276 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16277 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16278 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16279 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16280 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16281 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16282 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16283 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16284 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16285 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16286 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16287 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16288 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16289 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16290 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16291 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16292 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16293 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16294 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16295 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16296 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16297 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16298 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16299 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16300 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16301 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16302 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16303 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16304 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16305 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16306 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16307 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16308 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16309 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16310 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16311 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16312 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16313 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16314 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16315 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16316 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16317 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16318 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16319 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16320 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16321 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16322 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16323 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16324 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16325 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16326 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16327 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16328 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16329 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16330 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16331 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16332 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16333 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16334 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16335 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16336 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16337 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16338 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16339 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16340 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16341 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16342 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16343 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16344 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16345 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16346 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16347 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16348 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16349 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16350 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16351 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16352 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16353 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16354 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16355 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16356 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16357 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16358 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16359 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16360 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16361 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16362 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16363 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16364 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16365 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16366 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16367 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16368 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16369 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16370 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16371 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16372 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16373 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16374 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16375 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16376 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16377 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16378 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16379 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16380 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16381 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16382 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16383 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16384 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16385 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16386 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16387 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16388 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16389 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16390 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16391 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16392 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16393 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16394 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16395 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16396 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16397 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16398 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16399 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16400 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16401 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16402 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16403 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16404 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16405 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16406 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16407 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16408 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16409 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16410 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16411 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16412 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16413 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16414 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16415 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16416 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16417 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16418 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16419 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16420 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16421 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16422 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16423 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16424 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16425 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16426 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16427 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16428 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16429 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16430 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16431 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16432 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16433 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16434 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16435 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16436 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16437 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16438 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16439 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16440 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16441 => to_unsigned(32767, LUT_AMPL_WIDTH - 1),
		16442 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16443 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16444 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16445 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16446 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16447 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16448 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16449 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16450 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16451 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16452 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16453 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16454 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16455 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16456 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16457 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16458 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16459 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16460 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16461 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16462 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16463 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16464 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16465 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16466 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16467 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16468 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16469 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16470 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16471 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16472 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16473 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16474 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16475 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16476 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16477 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16478 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16479 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16480 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16481 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16482 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16483 => to_unsigned(32766, LUT_AMPL_WIDTH - 1),
		16484 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16485 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16486 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16487 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16488 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16489 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16490 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16491 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16492 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16493 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16494 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16495 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16496 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16497 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16498 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16499 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16500 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16501 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16502 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16503 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16504 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16505 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16506 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16507 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16508 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16509 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16510 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16511 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16512 => to_unsigned(32765, LUT_AMPL_WIDTH - 1),
		16513 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16514 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16515 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16516 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16517 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16518 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16519 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16520 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16521 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16522 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16523 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16524 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16525 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16526 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16527 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16528 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16529 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16530 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16531 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16532 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16533 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16534 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16535 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16536 => to_unsigned(32764, LUT_AMPL_WIDTH - 1),
		16537 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16538 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16539 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16540 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16541 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16542 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16543 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16544 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16545 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16546 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16547 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16548 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16549 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16550 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16551 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16552 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16553 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16554 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16555 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16556 => to_unsigned(32763, LUT_AMPL_WIDTH - 1),
		16557 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16558 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16559 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16560 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16561 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16562 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16563 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16564 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16565 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16566 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16567 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16568 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16569 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16570 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16571 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16572 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16573 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16574 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16575 => to_unsigned(32762, LUT_AMPL_WIDTH - 1),
		16576 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16577 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16578 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16579 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16580 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16581 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16582 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16583 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16584 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16585 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16586 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16587 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16588 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16589 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16590 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16591 => to_unsigned(32761, LUT_AMPL_WIDTH - 1),
		16592 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16593 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16594 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16595 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16596 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16597 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16598 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16599 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16600 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16601 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16602 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16603 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16604 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16605 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16606 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16607 => to_unsigned(32760, LUT_AMPL_WIDTH - 1),
		16608 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16609 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16610 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16611 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16612 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16613 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16614 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16615 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16616 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16617 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16618 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16619 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16620 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16621 => to_unsigned(32759, LUT_AMPL_WIDTH - 1),
		16622 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16623 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16624 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16625 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16626 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16627 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16628 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16629 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16630 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16631 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16632 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16633 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16634 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16635 => to_unsigned(32758, LUT_AMPL_WIDTH - 1),
		16636 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16637 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16638 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16639 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16640 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16641 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16642 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16643 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16644 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16645 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16646 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16647 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16648 => to_unsigned(32757, LUT_AMPL_WIDTH - 1),
		16649 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16650 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16651 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16652 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16653 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16654 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16655 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16656 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16657 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16658 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16659 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16660 => to_unsigned(32756, LUT_AMPL_WIDTH - 1),
		16661 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16662 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16663 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16664 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16665 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16666 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16667 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16668 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16669 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16670 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16671 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16672 => to_unsigned(32755, LUT_AMPL_WIDTH - 1),
		16673 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16674 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16675 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16676 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16677 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16678 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16679 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16680 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16681 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16682 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16683 => to_unsigned(32754, LUT_AMPL_WIDTH - 1),
		16684 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16685 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16686 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16687 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16688 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16689 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16690 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16691 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16692 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16693 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16694 => to_unsigned(32753, LUT_AMPL_WIDTH - 1),
		16695 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16696 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16697 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16698 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16699 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16700 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16701 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16702 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16703 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16704 => to_unsigned(32752, LUT_AMPL_WIDTH - 1),
		16705 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16706 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16707 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16708 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16709 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16710 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16711 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16712 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16713 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16714 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16715 => to_unsigned(32751, LUT_AMPL_WIDTH - 1),
		16716 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16717 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16718 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16719 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16720 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16721 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16722 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16723 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16724 => to_unsigned(32750, LUT_AMPL_WIDTH - 1),
		16725 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16726 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16727 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16728 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16729 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16730 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16731 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16732 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16733 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16734 => to_unsigned(32749, LUT_AMPL_WIDTH - 1),
		16735 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16736 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16737 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16738 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16739 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16740 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16741 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16742 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16743 => to_unsigned(32748, LUT_AMPL_WIDTH - 1),
		16744 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16745 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16746 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16747 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16748 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16749 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16750 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16751 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16752 => to_unsigned(32747, LUT_AMPL_WIDTH - 1),
		16753 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16754 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16755 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16756 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16757 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16758 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16759 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16760 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16761 => to_unsigned(32746, LUT_AMPL_WIDTH - 1),
		16762 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16763 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16764 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16765 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16766 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16767 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16768 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16769 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16770 => to_unsigned(32745, LUT_AMPL_WIDTH - 1),
		16771 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		16772 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		16773 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		16774 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		16775 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		16776 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		16777 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		16778 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		16779 => to_unsigned(32744, LUT_AMPL_WIDTH - 1),
		16780 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		16781 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		16782 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		16783 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		16784 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		16785 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		16786 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		16787 => to_unsigned(32743, LUT_AMPL_WIDTH - 1),
		16788 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		16789 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		16790 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		16791 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		16792 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		16793 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		16794 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		16795 => to_unsigned(32742, LUT_AMPL_WIDTH - 1),
		16796 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		16797 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		16798 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		16799 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		16800 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		16801 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		16802 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		16803 => to_unsigned(32741, LUT_AMPL_WIDTH - 1),
		16804 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		16805 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		16806 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		16807 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		16808 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		16809 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		16810 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		16811 => to_unsigned(32740, LUT_AMPL_WIDTH - 1),
		16812 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		16813 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		16814 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		16815 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		16816 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		16817 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		16818 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		16819 => to_unsigned(32739, LUT_AMPL_WIDTH - 1),
		16820 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		16821 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		16822 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		16823 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		16824 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		16825 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		16826 => to_unsigned(32738, LUT_AMPL_WIDTH - 1),
		16827 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		16828 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		16829 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		16830 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		16831 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		16832 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		16833 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		16834 => to_unsigned(32737, LUT_AMPL_WIDTH - 1),
		16835 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		16836 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		16837 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		16838 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		16839 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		16840 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		16841 => to_unsigned(32736, LUT_AMPL_WIDTH - 1),
		16842 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		16843 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		16844 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		16845 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		16846 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		16847 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		16848 => to_unsigned(32735, LUT_AMPL_WIDTH - 1),
		16849 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		16850 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		16851 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		16852 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		16853 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		16854 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		16855 => to_unsigned(32734, LUT_AMPL_WIDTH - 1),
		16856 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		16857 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		16858 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		16859 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		16860 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		16861 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		16862 => to_unsigned(32733, LUT_AMPL_WIDTH - 1),
		16863 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		16864 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		16865 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		16866 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		16867 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		16868 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		16869 => to_unsigned(32732, LUT_AMPL_WIDTH - 1),
		16870 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		16871 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		16872 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		16873 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		16874 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		16875 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		16876 => to_unsigned(32731, LUT_AMPL_WIDTH - 1),
		16877 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		16878 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		16879 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		16880 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		16881 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		16882 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		16883 => to_unsigned(32730, LUT_AMPL_WIDTH - 1),
		16884 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		16885 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		16886 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		16887 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		16888 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		16889 => to_unsigned(32729, LUT_AMPL_WIDTH - 1),
		16890 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		16891 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		16892 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		16893 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		16894 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		16895 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		16896 => to_unsigned(32728, LUT_AMPL_WIDTH - 1),
		16897 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		16898 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		16899 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		16900 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		16901 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		16902 => to_unsigned(32727, LUT_AMPL_WIDTH - 1),
		16903 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		16904 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		16905 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		16906 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		16907 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		16908 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		16909 => to_unsigned(32726, LUT_AMPL_WIDTH - 1),
		16910 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		16911 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		16912 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		16913 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		16914 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		16915 => to_unsigned(32725, LUT_AMPL_WIDTH - 1),
		16916 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		16917 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		16918 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		16919 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		16920 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		16921 => to_unsigned(32724, LUT_AMPL_WIDTH - 1),
		16922 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		16923 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		16924 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		16925 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		16926 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		16927 => to_unsigned(32723, LUT_AMPL_WIDTH - 1),
		16928 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		16929 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		16930 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		16931 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		16932 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		16933 => to_unsigned(32722, LUT_AMPL_WIDTH - 1),
		16934 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		16935 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		16936 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		16937 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		16938 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		16939 => to_unsigned(32721, LUT_AMPL_WIDTH - 1),
		16940 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		16941 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		16942 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		16943 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		16944 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		16945 => to_unsigned(32720, LUT_AMPL_WIDTH - 1),
		16946 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		16947 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		16948 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		16949 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		16950 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		16951 => to_unsigned(32719, LUT_AMPL_WIDTH - 1),
		16952 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		16953 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		16954 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		16955 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		16956 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		16957 => to_unsigned(32718, LUT_AMPL_WIDTH - 1),
		16958 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		16959 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		16960 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		16961 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		16962 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		16963 => to_unsigned(32717, LUT_AMPL_WIDTH - 1),
		16964 => to_unsigned(32716, LUT_AMPL_WIDTH - 1),
		16965 => to_unsigned(32716, LUT_AMPL_WIDTH - 1),
		16966 => to_unsigned(32716, LUT_AMPL_WIDTH - 1),
		16967 => to_unsigned(32716, LUT_AMPL_WIDTH - 1),
		16968 => to_unsigned(32716, LUT_AMPL_WIDTH - 1),
		16969 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		16970 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		16971 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		16972 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		16973 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		16974 => to_unsigned(32715, LUT_AMPL_WIDTH - 1),
		16975 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		16976 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		16977 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		16978 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		16979 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		16980 => to_unsigned(32714, LUT_AMPL_WIDTH - 1),
		16981 => to_unsigned(32713, LUT_AMPL_WIDTH - 1),
		16982 => to_unsigned(32713, LUT_AMPL_WIDTH - 1),
		16983 => to_unsigned(32713, LUT_AMPL_WIDTH - 1),
		16984 => to_unsigned(32713, LUT_AMPL_WIDTH - 1),
		16985 => to_unsigned(32713, LUT_AMPL_WIDTH - 1),
		16986 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		16987 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		16988 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		16989 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		16990 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		16991 => to_unsigned(32712, LUT_AMPL_WIDTH - 1),
		16992 => to_unsigned(32711, LUT_AMPL_WIDTH - 1),
		16993 => to_unsigned(32711, LUT_AMPL_WIDTH - 1),
		16994 => to_unsigned(32711, LUT_AMPL_WIDTH - 1),
		16995 => to_unsigned(32711, LUT_AMPL_WIDTH - 1),
		16996 => to_unsigned(32711, LUT_AMPL_WIDTH - 1),
		16997 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		16998 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		16999 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		17000 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		17001 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		17002 => to_unsigned(32710, LUT_AMPL_WIDTH - 1),
		17003 => to_unsigned(32709, LUT_AMPL_WIDTH - 1),
		17004 => to_unsigned(32709, LUT_AMPL_WIDTH - 1),
		17005 => to_unsigned(32709, LUT_AMPL_WIDTH - 1),
		17006 => to_unsigned(32709, LUT_AMPL_WIDTH - 1),
		17007 => to_unsigned(32709, LUT_AMPL_WIDTH - 1),
		17008 => to_unsigned(32708, LUT_AMPL_WIDTH - 1),
		17009 => to_unsigned(32708, LUT_AMPL_WIDTH - 1),
		17010 => to_unsigned(32708, LUT_AMPL_WIDTH - 1),
		17011 => to_unsigned(32708, LUT_AMPL_WIDTH - 1),
		17012 => to_unsigned(32708, LUT_AMPL_WIDTH - 1),
		17013 => to_unsigned(32707, LUT_AMPL_WIDTH - 1),
		17014 => to_unsigned(32707, LUT_AMPL_WIDTH - 1),
		17015 => to_unsigned(32707, LUT_AMPL_WIDTH - 1),
		17016 => to_unsigned(32707, LUT_AMPL_WIDTH - 1),
		17017 => to_unsigned(32707, LUT_AMPL_WIDTH - 1),
		17018 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		17019 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		17020 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		17021 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		17022 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		17023 => to_unsigned(32706, LUT_AMPL_WIDTH - 1),
		17024 => to_unsigned(32705, LUT_AMPL_WIDTH - 1),
		17025 => to_unsigned(32705, LUT_AMPL_WIDTH - 1),
		17026 => to_unsigned(32705, LUT_AMPL_WIDTH - 1),
		17027 => to_unsigned(32705, LUT_AMPL_WIDTH - 1),
		17028 => to_unsigned(32705, LUT_AMPL_WIDTH - 1),
		17029 => to_unsigned(32704, LUT_AMPL_WIDTH - 1),
		17030 => to_unsigned(32704, LUT_AMPL_WIDTH - 1),
		17031 => to_unsigned(32704, LUT_AMPL_WIDTH - 1),
		17032 => to_unsigned(32704, LUT_AMPL_WIDTH - 1),
		17033 => to_unsigned(32704, LUT_AMPL_WIDTH - 1),
		17034 => to_unsigned(32703, LUT_AMPL_WIDTH - 1),
		17035 => to_unsigned(32703, LUT_AMPL_WIDTH - 1),
		17036 => to_unsigned(32703, LUT_AMPL_WIDTH - 1),
		17037 => to_unsigned(32703, LUT_AMPL_WIDTH - 1),
		17038 => to_unsigned(32703, LUT_AMPL_WIDTH - 1),
		17039 => to_unsigned(32702, LUT_AMPL_WIDTH - 1),
		17040 => to_unsigned(32702, LUT_AMPL_WIDTH - 1),
		17041 => to_unsigned(32702, LUT_AMPL_WIDTH - 1),
		17042 => to_unsigned(32702, LUT_AMPL_WIDTH - 1),
		17043 => to_unsigned(32702, LUT_AMPL_WIDTH - 1),
		17044 => to_unsigned(32701, LUT_AMPL_WIDTH - 1),
		17045 => to_unsigned(32701, LUT_AMPL_WIDTH - 1),
		17046 => to_unsigned(32701, LUT_AMPL_WIDTH - 1),
		17047 => to_unsigned(32701, LUT_AMPL_WIDTH - 1),
		17048 => to_unsigned(32701, LUT_AMPL_WIDTH - 1),
		17049 => to_unsigned(32700, LUT_AMPL_WIDTH - 1),
		17050 => to_unsigned(32700, LUT_AMPL_WIDTH - 1),
		17051 => to_unsigned(32700, LUT_AMPL_WIDTH - 1),
		17052 => to_unsigned(32700, LUT_AMPL_WIDTH - 1),
		17053 => to_unsigned(32700, LUT_AMPL_WIDTH - 1),
		17054 => to_unsigned(32699, LUT_AMPL_WIDTH - 1),
		17055 => to_unsigned(32699, LUT_AMPL_WIDTH - 1),
		17056 => to_unsigned(32699, LUT_AMPL_WIDTH - 1),
		17057 => to_unsigned(32699, LUT_AMPL_WIDTH - 1),
		17058 => to_unsigned(32699, LUT_AMPL_WIDTH - 1),
		17059 => to_unsigned(32698, LUT_AMPL_WIDTH - 1),
		17060 => to_unsigned(32698, LUT_AMPL_WIDTH - 1),
		17061 => to_unsigned(32698, LUT_AMPL_WIDTH - 1),
		17062 => to_unsigned(32698, LUT_AMPL_WIDTH - 1),
		17063 => to_unsigned(32698, LUT_AMPL_WIDTH - 1),
		17064 => to_unsigned(32697, LUT_AMPL_WIDTH - 1),
		17065 => to_unsigned(32697, LUT_AMPL_WIDTH - 1),
		17066 => to_unsigned(32697, LUT_AMPL_WIDTH - 1),
		17067 => to_unsigned(32697, LUT_AMPL_WIDTH - 1),
		17068 => to_unsigned(32697, LUT_AMPL_WIDTH - 1),
		17069 => to_unsigned(32696, LUT_AMPL_WIDTH - 1),
		17070 => to_unsigned(32696, LUT_AMPL_WIDTH - 1),
		17071 => to_unsigned(32696, LUT_AMPL_WIDTH - 1),
		17072 => to_unsigned(32696, LUT_AMPL_WIDTH - 1),
		17073 => to_unsigned(32696, LUT_AMPL_WIDTH - 1),
		17074 => to_unsigned(32695, LUT_AMPL_WIDTH - 1),
		17075 => to_unsigned(32695, LUT_AMPL_WIDTH - 1),
		17076 => to_unsigned(32695, LUT_AMPL_WIDTH - 1),
		17077 => to_unsigned(32695, LUT_AMPL_WIDTH - 1),
		17078 => to_unsigned(32694, LUT_AMPL_WIDTH - 1),
		17079 => to_unsigned(32694, LUT_AMPL_WIDTH - 1),
		17080 => to_unsigned(32694, LUT_AMPL_WIDTH - 1),
		17081 => to_unsigned(32694, LUT_AMPL_WIDTH - 1),
		17082 => to_unsigned(32694, LUT_AMPL_WIDTH - 1),
		17083 => to_unsigned(32693, LUT_AMPL_WIDTH - 1),
		17084 => to_unsigned(32693, LUT_AMPL_WIDTH - 1),
		17085 => to_unsigned(32693, LUT_AMPL_WIDTH - 1),
		17086 => to_unsigned(32693, LUT_AMPL_WIDTH - 1),
		17087 => to_unsigned(32693, LUT_AMPL_WIDTH - 1),
		17088 => to_unsigned(32692, LUT_AMPL_WIDTH - 1),
		17089 => to_unsigned(32692, LUT_AMPL_WIDTH - 1),
		17090 => to_unsigned(32692, LUT_AMPL_WIDTH - 1),
		17091 => to_unsigned(32692, LUT_AMPL_WIDTH - 1),
		17092 => to_unsigned(32692, LUT_AMPL_WIDTH - 1),
		17093 => to_unsigned(32691, LUT_AMPL_WIDTH - 1),
		17094 => to_unsigned(32691, LUT_AMPL_WIDTH - 1),
		17095 => to_unsigned(32691, LUT_AMPL_WIDTH - 1),
		17096 => to_unsigned(32691, LUT_AMPL_WIDTH - 1),
		17097 => to_unsigned(32690, LUT_AMPL_WIDTH - 1),
		17098 => to_unsigned(32690, LUT_AMPL_WIDTH - 1),
		17099 => to_unsigned(32690, LUT_AMPL_WIDTH - 1),
		17100 => to_unsigned(32690, LUT_AMPL_WIDTH - 1),
		17101 => to_unsigned(32690, LUT_AMPL_WIDTH - 1),
		17102 => to_unsigned(32689, LUT_AMPL_WIDTH - 1),
		17103 => to_unsigned(32689, LUT_AMPL_WIDTH - 1),
		17104 => to_unsigned(32689, LUT_AMPL_WIDTH - 1),
		17105 => to_unsigned(32689, LUT_AMPL_WIDTH - 1),
		17106 => to_unsigned(32689, LUT_AMPL_WIDTH - 1),
		17107 => to_unsigned(32688, LUT_AMPL_WIDTH - 1),
		17108 => to_unsigned(32688, LUT_AMPL_WIDTH - 1),
		17109 => to_unsigned(32688, LUT_AMPL_WIDTH - 1),
		17110 => to_unsigned(32688, LUT_AMPL_WIDTH - 1),
		17111 => to_unsigned(32687, LUT_AMPL_WIDTH - 1),
		17112 => to_unsigned(32687, LUT_AMPL_WIDTH - 1),
		17113 => to_unsigned(32687, LUT_AMPL_WIDTH - 1),
		17114 => to_unsigned(32687, LUT_AMPL_WIDTH - 1),
		17115 => to_unsigned(32687, LUT_AMPL_WIDTH - 1),
		17116 => to_unsigned(32686, LUT_AMPL_WIDTH - 1),
		17117 => to_unsigned(32686, LUT_AMPL_WIDTH - 1),
		17118 => to_unsigned(32686, LUT_AMPL_WIDTH - 1),
		17119 => to_unsigned(32686, LUT_AMPL_WIDTH - 1),
		17120 => to_unsigned(32685, LUT_AMPL_WIDTH - 1),
		17121 => to_unsigned(32685, LUT_AMPL_WIDTH - 1),
		17122 => to_unsigned(32685, LUT_AMPL_WIDTH - 1),
		17123 => to_unsigned(32685, LUT_AMPL_WIDTH - 1),
		17124 => to_unsigned(32685, LUT_AMPL_WIDTH - 1),
		17125 => to_unsigned(32684, LUT_AMPL_WIDTH - 1),
		17126 => to_unsigned(32684, LUT_AMPL_WIDTH - 1),
		17127 => to_unsigned(32684, LUT_AMPL_WIDTH - 1),
		17128 => to_unsigned(32684, LUT_AMPL_WIDTH - 1),
		17129 => to_unsigned(32683, LUT_AMPL_WIDTH - 1),
		17130 => to_unsigned(32683, LUT_AMPL_WIDTH - 1),
		17131 => to_unsigned(32683, LUT_AMPL_WIDTH - 1),
		17132 => to_unsigned(32683, LUT_AMPL_WIDTH - 1),
		17133 => to_unsigned(32683, LUT_AMPL_WIDTH - 1),
		17134 => to_unsigned(32682, LUT_AMPL_WIDTH - 1),
		17135 => to_unsigned(32682, LUT_AMPL_WIDTH - 1),
		17136 => to_unsigned(32682, LUT_AMPL_WIDTH - 1),
		17137 => to_unsigned(32682, LUT_AMPL_WIDTH - 1),
		17138 => to_unsigned(32681, LUT_AMPL_WIDTH - 1),
		17139 => to_unsigned(32681, LUT_AMPL_WIDTH - 1),
		17140 => to_unsigned(32681, LUT_AMPL_WIDTH - 1),
		17141 => to_unsigned(32681, LUT_AMPL_WIDTH - 1),
		17142 => to_unsigned(32681, LUT_AMPL_WIDTH - 1),
		17143 => to_unsigned(32680, LUT_AMPL_WIDTH - 1),
		17144 => to_unsigned(32680, LUT_AMPL_WIDTH - 1),
		17145 => to_unsigned(32680, LUT_AMPL_WIDTH - 1),
		17146 => to_unsigned(32680, LUT_AMPL_WIDTH - 1),
		17147 => to_unsigned(32679, LUT_AMPL_WIDTH - 1),
		17148 => to_unsigned(32679, LUT_AMPL_WIDTH - 1),
		17149 => to_unsigned(32679, LUT_AMPL_WIDTH - 1),
		17150 => to_unsigned(32679, LUT_AMPL_WIDTH - 1),
		17151 => to_unsigned(32678, LUT_AMPL_WIDTH - 1),
		17152 => to_unsigned(32678, LUT_AMPL_WIDTH - 1),
		17153 => to_unsigned(32678, LUT_AMPL_WIDTH - 1),
		17154 => to_unsigned(32678, LUT_AMPL_WIDTH - 1),
		17155 => to_unsigned(32678, LUT_AMPL_WIDTH - 1),
		17156 => to_unsigned(32677, LUT_AMPL_WIDTH - 1),
		17157 => to_unsigned(32677, LUT_AMPL_WIDTH - 1),
		17158 => to_unsigned(32677, LUT_AMPL_WIDTH - 1),
		17159 => to_unsigned(32677, LUT_AMPL_WIDTH - 1),
		17160 => to_unsigned(32676, LUT_AMPL_WIDTH - 1),
		17161 => to_unsigned(32676, LUT_AMPL_WIDTH - 1),
		17162 => to_unsigned(32676, LUT_AMPL_WIDTH - 1),
		17163 => to_unsigned(32676, LUT_AMPL_WIDTH - 1),
		17164 => to_unsigned(32675, LUT_AMPL_WIDTH - 1),
		17165 => to_unsigned(32675, LUT_AMPL_WIDTH - 1),
		17166 => to_unsigned(32675, LUT_AMPL_WIDTH - 1),
		17167 => to_unsigned(32675, LUT_AMPL_WIDTH - 1),
		17168 => to_unsigned(32674, LUT_AMPL_WIDTH - 1),
		17169 => to_unsigned(32674, LUT_AMPL_WIDTH - 1),
		17170 => to_unsigned(32674, LUT_AMPL_WIDTH - 1),
		17171 => to_unsigned(32674, LUT_AMPL_WIDTH - 1),
		17172 => to_unsigned(32674, LUT_AMPL_WIDTH - 1),
		17173 => to_unsigned(32673, LUT_AMPL_WIDTH - 1),
		17174 => to_unsigned(32673, LUT_AMPL_WIDTH - 1),
		17175 => to_unsigned(32673, LUT_AMPL_WIDTH - 1),
		17176 => to_unsigned(32673, LUT_AMPL_WIDTH - 1),
		17177 => to_unsigned(32672, LUT_AMPL_WIDTH - 1),
		17178 => to_unsigned(32672, LUT_AMPL_WIDTH - 1),
		17179 => to_unsigned(32672, LUT_AMPL_WIDTH - 1),
		17180 => to_unsigned(32672, LUT_AMPL_WIDTH - 1),
		17181 => to_unsigned(32671, LUT_AMPL_WIDTH - 1),
		17182 => to_unsigned(32671, LUT_AMPL_WIDTH - 1),
		17183 => to_unsigned(32671, LUT_AMPL_WIDTH - 1),
		17184 => to_unsigned(32671, LUT_AMPL_WIDTH - 1),
		17185 => to_unsigned(32670, LUT_AMPL_WIDTH - 1),
		17186 => to_unsigned(32670, LUT_AMPL_WIDTH - 1),
		17187 => to_unsigned(32670, LUT_AMPL_WIDTH - 1),
		17188 => to_unsigned(32670, LUT_AMPL_WIDTH - 1),
		17189 => to_unsigned(32669, LUT_AMPL_WIDTH - 1),
		17190 => to_unsigned(32669, LUT_AMPL_WIDTH - 1),
		17191 => to_unsigned(32669, LUT_AMPL_WIDTH - 1),
		17192 => to_unsigned(32669, LUT_AMPL_WIDTH - 1),
		17193 => to_unsigned(32668, LUT_AMPL_WIDTH - 1),
		17194 => to_unsigned(32668, LUT_AMPL_WIDTH - 1),
		17195 => to_unsigned(32668, LUT_AMPL_WIDTH - 1),
		17196 => to_unsigned(32668, LUT_AMPL_WIDTH - 1),
		17197 => to_unsigned(32668, LUT_AMPL_WIDTH - 1),
		17198 => to_unsigned(32667, LUT_AMPL_WIDTH - 1),
		17199 => to_unsigned(32667, LUT_AMPL_WIDTH - 1),
		17200 => to_unsigned(32667, LUT_AMPL_WIDTH - 1),
		17201 => to_unsigned(32667, LUT_AMPL_WIDTH - 1),
		17202 => to_unsigned(32666, LUT_AMPL_WIDTH - 1),
		17203 => to_unsigned(32666, LUT_AMPL_WIDTH - 1),
		17204 => to_unsigned(32666, LUT_AMPL_WIDTH - 1),
		17205 => to_unsigned(32666, LUT_AMPL_WIDTH - 1),
		17206 => to_unsigned(32665, LUT_AMPL_WIDTH - 1),
		17207 => to_unsigned(32665, LUT_AMPL_WIDTH - 1),
		17208 => to_unsigned(32665, LUT_AMPL_WIDTH - 1),
		17209 => to_unsigned(32665, LUT_AMPL_WIDTH - 1),
		17210 => to_unsigned(32664, LUT_AMPL_WIDTH - 1),
		17211 => to_unsigned(32664, LUT_AMPL_WIDTH - 1),
		17212 => to_unsigned(32664, LUT_AMPL_WIDTH - 1),
		17213 => to_unsigned(32664, LUT_AMPL_WIDTH - 1),
		17214 => to_unsigned(32663, LUT_AMPL_WIDTH - 1),
		17215 => to_unsigned(32663, LUT_AMPL_WIDTH - 1),
		17216 => to_unsigned(32663, LUT_AMPL_WIDTH - 1),
		17217 => to_unsigned(32663, LUT_AMPL_WIDTH - 1),
		17218 => to_unsigned(32662, LUT_AMPL_WIDTH - 1),
		17219 => to_unsigned(32662, LUT_AMPL_WIDTH - 1),
		17220 => to_unsigned(32662, LUT_AMPL_WIDTH - 1),
		17221 => to_unsigned(32662, LUT_AMPL_WIDTH - 1),
		17222 => to_unsigned(32661, LUT_AMPL_WIDTH - 1),
		17223 => to_unsigned(32661, LUT_AMPL_WIDTH - 1),
		17224 => to_unsigned(32661, LUT_AMPL_WIDTH - 1),
		17225 => to_unsigned(32661, LUT_AMPL_WIDTH - 1),
		17226 => to_unsigned(32660, LUT_AMPL_WIDTH - 1),
		17227 => to_unsigned(32660, LUT_AMPL_WIDTH - 1),
		17228 => to_unsigned(32660, LUT_AMPL_WIDTH - 1),
		17229 => to_unsigned(32660, LUT_AMPL_WIDTH - 1),
		17230 => to_unsigned(32659, LUT_AMPL_WIDTH - 1),
		17231 => to_unsigned(32659, LUT_AMPL_WIDTH - 1),
		17232 => to_unsigned(32659, LUT_AMPL_WIDTH - 1),
		17233 => to_unsigned(32659, LUT_AMPL_WIDTH - 1),
		17234 => to_unsigned(32658, LUT_AMPL_WIDTH - 1),
		17235 => to_unsigned(32658, LUT_AMPL_WIDTH - 1),
		17236 => to_unsigned(32658, LUT_AMPL_WIDTH - 1),
		17237 => to_unsigned(32657, LUT_AMPL_WIDTH - 1),
		17238 => to_unsigned(32657, LUT_AMPL_WIDTH - 1),
		17239 => to_unsigned(32657, LUT_AMPL_WIDTH - 1),
		17240 => to_unsigned(32657, LUT_AMPL_WIDTH - 1),
		17241 => to_unsigned(32656, LUT_AMPL_WIDTH - 1),
		17242 => to_unsigned(32656, LUT_AMPL_WIDTH - 1),
		17243 => to_unsigned(32656, LUT_AMPL_WIDTH - 1),
		17244 => to_unsigned(32656, LUT_AMPL_WIDTH - 1),
		17245 => to_unsigned(32655, LUT_AMPL_WIDTH - 1),
		17246 => to_unsigned(32655, LUT_AMPL_WIDTH - 1),
		17247 => to_unsigned(32655, LUT_AMPL_WIDTH - 1),
		17248 => to_unsigned(32655, LUT_AMPL_WIDTH - 1),
		17249 => to_unsigned(32654, LUT_AMPL_WIDTH - 1),
		17250 => to_unsigned(32654, LUT_AMPL_WIDTH - 1),
		17251 => to_unsigned(32654, LUT_AMPL_WIDTH - 1),
		17252 => to_unsigned(32654, LUT_AMPL_WIDTH - 1),
		17253 => to_unsigned(32653, LUT_AMPL_WIDTH - 1),
		17254 => to_unsigned(32653, LUT_AMPL_WIDTH - 1),
		17255 => to_unsigned(32653, LUT_AMPL_WIDTH - 1),
		17256 => to_unsigned(32653, LUT_AMPL_WIDTH - 1),
		17257 => to_unsigned(32652, LUT_AMPL_WIDTH - 1),
		17258 => to_unsigned(32652, LUT_AMPL_WIDTH - 1),
		17259 => to_unsigned(32652, LUT_AMPL_WIDTH - 1),
		17260 => to_unsigned(32652, LUT_AMPL_WIDTH - 1),
		17261 => to_unsigned(32651, LUT_AMPL_WIDTH - 1),
		17262 => to_unsigned(32651, LUT_AMPL_WIDTH - 1),
		17263 => to_unsigned(32651, LUT_AMPL_WIDTH - 1),
		17264 => to_unsigned(32650, LUT_AMPL_WIDTH - 1),
		17265 => to_unsigned(32650, LUT_AMPL_WIDTH - 1),
		17266 => to_unsigned(32650, LUT_AMPL_WIDTH - 1),
		17267 => to_unsigned(32650, LUT_AMPL_WIDTH - 1),
		17268 => to_unsigned(32649, LUT_AMPL_WIDTH - 1),
		17269 => to_unsigned(32649, LUT_AMPL_WIDTH - 1),
		17270 => to_unsigned(32649, LUT_AMPL_WIDTH - 1),
		17271 => to_unsigned(32649, LUT_AMPL_WIDTH - 1),
		17272 => to_unsigned(32648, LUT_AMPL_WIDTH - 1),
		17273 => to_unsigned(32648, LUT_AMPL_WIDTH - 1),
		17274 => to_unsigned(32648, LUT_AMPL_WIDTH - 1),
		17275 => to_unsigned(32648, LUT_AMPL_WIDTH - 1),
		17276 => to_unsigned(32647, LUT_AMPL_WIDTH - 1),
		17277 => to_unsigned(32647, LUT_AMPL_WIDTH - 1),
		17278 => to_unsigned(32647, LUT_AMPL_WIDTH - 1),
		17279 => to_unsigned(32646, LUT_AMPL_WIDTH - 1),
		17280 => to_unsigned(32646, LUT_AMPL_WIDTH - 1),
		17281 => to_unsigned(32646, LUT_AMPL_WIDTH - 1),
		17282 => to_unsigned(32646, LUT_AMPL_WIDTH - 1),
		17283 => to_unsigned(32645, LUT_AMPL_WIDTH - 1),
		17284 => to_unsigned(32645, LUT_AMPL_WIDTH - 1),
		17285 => to_unsigned(32645, LUT_AMPL_WIDTH - 1),
		17286 => to_unsigned(32645, LUT_AMPL_WIDTH - 1),
		17287 => to_unsigned(32644, LUT_AMPL_WIDTH - 1),
		17288 => to_unsigned(32644, LUT_AMPL_WIDTH - 1),
		17289 => to_unsigned(32644, LUT_AMPL_WIDTH - 1),
		17290 => to_unsigned(32643, LUT_AMPL_WIDTH - 1),
		17291 => to_unsigned(32643, LUT_AMPL_WIDTH - 1),
		17292 => to_unsigned(32643, LUT_AMPL_WIDTH - 1),
		17293 => to_unsigned(32643, LUT_AMPL_WIDTH - 1),
		17294 => to_unsigned(32642, LUT_AMPL_WIDTH - 1),
		17295 => to_unsigned(32642, LUT_AMPL_WIDTH - 1),
		17296 => to_unsigned(32642, LUT_AMPL_WIDTH - 1),
		17297 => to_unsigned(32642, LUT_AMPL_WIDTH - 1),
		17298 => to_unsigned(32641, LUT_AMPL_WIDTH - 1),
		17299 => to_unsigned(32641, LUT_AMPL_WIDTH - 1),
		17300 => to_unsigned(32641, LUT_AMPL_WIDTH - 1),
		17301 => to_unsigned(32640, LUT_AMPL_WIDTH - 1),
		17302 => to_unsigned(32640, LUT_AMPL_WIDTH - 1),
		17303 => to_unsigned(32640, LUT_AMPL_WIDTH - 1),
		17304 => to_unsigned(32640, LUT_AMPL_WIDTH - 1),
		17305 => to_unsigned(32639, LUT_AMPL_WIDTH - 1),
		17306 => to_unsigned(32639, LUT_AMPL_WIDTH - 1),
		17307 => to_unsigned(32639, LUT_AMPL_WIDTH - 1),
		17308 => to_unsigned(32639, LUT_AMPL_WIDTH - 1),
		17309 => to_unsigned(32638, LUT_AMPL_WIDTH - 1),
		17310 => to_unsigned(32638, LUT_AMPL_WIDTH - 1),
		17311 => to_unsigned(32638, LUT_AMPL_WIDTH - 1),
		17312 => to_unsigned(32637, LUT_AMPL_WIDTH - 1),
		17313 => to_unsigned(32637, LUT_AMPL_WIDTH - 1),
		17314 => to_unsigned(32637, LUT_AMPL_WIDTH - 1),
		17315 => to_unsigned(32637, LUT_AMPL_WIDTH - 1),
		17316 => to_unsigned(32636, LUT_AMPL_WIDTH - 1),
		17317 => to_unsigned(32636, LUT_AMPL_WIDTH - 1),
		17318 => to_unsigned(32636, LUT_AMPL_WIDTH - 1),
		17319 => to_unsigned(32635, LUT_AMPL_WIDTH - 1),
		17320 => to_unsigned(32635, LUT_AMPL_WIDTH - 1),
		17321 => to_unsigned(32635, LUT_AMPL_WIDTH - 1),
		17322 => to_unsigned(32635, LUT_AMPL_WIDTH - 1),
		17323 => to_unsigned(32634, LUT_AMPL_WIDTH - 1),
		17324 => to_unsigned(32634, LUT_AMPL_WIDTH - 1),
		17325 => to_unsigned(32634, LUT_AMPL_WIDTH - 1),
		17326 => to_unsigned(32633, LUT_AMPL_WIDTH - 1),
		17327 => to_unsigned(32633, LUT_AMPL_WIDTH - 1),
		17328 => to_unsigned(32633, LUT_AMPL_WIDTH - 1),
		17329 => to_unsigned(32633, LUT_AMPL_WIDTH - 1),
		17330 => to_unsigned(32632, LUT_AMPL_WIDTH - 1),
		17331 => to_unsigned(32632, LUT_AMPL_WIDTH - 1),
		17332 => to_unsigned(32632, LUT_AMPL_WIDTH - 1),
		17333 => to_unsigned(32631, LUT_AMPL_WIDTH - 1),
		17334 => to_unsigned(32631, LUT_AMPL_WIDTH - 1),
		17335 => to_unsigned(32631, LUT_AMPL_WIDTH - 1),
		17336 => to_unsigned(32631, LUT_AMPL_WIDTH - 1),
		17337 => to_unsigned(32630, LUT_AMPL_WIDTH - 1),
		17338 => to_unsigned(32630, LUT_AMPL_WIDTH - 1),
		17339 => to_unsigned(32630, LUT_AMPL_WIDTH - 1),
		17340 => to_unsigned(32629, LUT_AMPL_WIDTH - 1),
		17341 => to_unsigned(32629, LUT_AMPL_WIDTH - 1),
		17342 => to_unsigned(32629, LUT_AMPL_WIDTH - 1),
		17343 => to_unsigned(32629, LUT_AMPL_WIDTH - 1),
		17344 => to_unsigned(32628, LUT_AMPL_WIDTH - 1),
		17345 => to_unsigned(32628, LUT_AMPL_WIDTH - 1),
		17346 => to_unsigned(32628, LUT_AMPL_WIDTH - 1),
		17347 => to_unsigned(32627, LUT_AMPL_WIDTH - 1),
		17348 => to_unsigned(32627, LUT_AMPL_WIDTH - 1),
		17349 => to_unsigned(32627, LUT_AMPL_WIDTH - 1),
		17350 => to_unsigned(32627, LUT_AMPL_WIDTH - 1),
		17351 => to_unsigned(32626, LUT_AMPL_WIDTH - 1),
		17352 => to_unsigned(32626, LUT_AMPL_WIDTH - 1),
		17353 => to_unsigned(32626, LUT_AMPL_WIDTH - 1),
		17354 => to_unsigned(32625, LUT_AMPL_WIDTH - 1),
		17355 => to_unsigned(32625, LUT_AMPL_WIDTH - 1),
		17356 => to_unsigned(32625, LUT_AMPL_WIDTH - 1),
		17357 => to_unsigned(32625, LUT_AMPL_WIDTH - 1),
		17358 => to_unsigned(32624, LUT_AMPL_WIDTH - 1),
		17359 => to_unsigned(32624, LUT_AMPL_WIDTH - 1),
		17360 => to_unsigned(32624, LUT_AMPL_WIDTH - 1),
		17361 => to_unsigned(32623, LUT_AMPL_WIDTH - 1),
		17362 => to_unsigned(32623, LUT_AMPL_WIDTH - 1),
		17363 => to_unsigned(32623, LUT_AMPL_WIDTH - 1),
		17364 => to_unsigned(32622, LUT_AMPL_WIDTH - 1),
		17365 => to_unsigned(32622, LUT_AMPL_WIDTH - 1),
		17366 => to_unsigned(32622, LUT_AMPL_WIDTH - 1),
		17367 => to_unsigned(32622, LUT_AMPL_WIDTH - 1),
		17368 => to_unsigned(32621, LUT_AMPL_WIDTH - 1),
		17369 => to_unsigned(32621, LUT_AMPL_WIDTH - 1),
		17370 => to_unsigned(32621, LUT_AMPL_WIDTH - 1),
		17371 => to_unsigned(32620, LUT_AMPL_WIDTH - 1),
		17372 => to_unsigned(32620, LUT_AMPL_WIDTH - 1),
		17373 => to_unsigned(32620, LUT_AMPL_WIDTH - 1),
		17374 => to_unsigned(32620, LUT_AMPL_WIDTH - 1),
		17375 => to_unsigned(32619, LUT_AMPL_WIDTH - 1),
		17376 => to_unsigned(32619, LUT_AMPL_WIDTH - 1),
		17377 => to_unsigned(32619, LUT_AMPL_WIDTH - 1),
		17378 => to_unsigned(32618, LUT_AMPL_WIDTH - 1),
		17379 => to_unsigned(32618, LUT_AMPL_WIDTH - 1),
		17380 => to_unsigned(32618, LUT_AMPL_WIDTH - 1),
		17381 => to_unsigned(32617, LUT_AMPL_WIDTH - 1),
		17382 => to_unsigned(32617, LUT_AMPL_WIDTH - 1),
		17383 => to_unsigned(32617, LUT_AMPL_WIDTH - 1),
		17384 => to_unsigned(32617, LUT_AMPL_WIDTH - 1),
		17385 => to_unsigned(32616, LUT_AMPL_WIDTH - 1),
		17386 => to_unsigned(32616, LUT_AMPL_WIDTH - 1),
		17387 => to_unsigned(32616, LUT_AMPL_WIDTH - 1),
		17388 => to_unsigned(32615, LUT_AMPL_WIDTH - 1),
		17389 => to_unsigned(32615, LUT_AMPL_WIDTH - 1),
		17390 => to_unsigned(32615, LUT_AMPL_WIDTH - 1),
		17391 => to_unsigned(32614, LUT_AMPL_WIDTH - 1),
		17392 => to_unsigned(32614, LUT_AMPL_WIDTH - 1),
		17393 => to_unsigned(32614, LUT_AMPL_WIDTH - 1),
		17394 => to_unsigned(32613, LUT_AMPL_WIDTH - 1),
		17395 => to_unsigned(32613, LUT_AMPL_WIDTH - 1),
		17396 => to_unsigned(32613, LUT_AMPL_WIDTH - 1),
		17397 => to_unsigned(32613, LUT_AMPL_WIDTH - 1),
		17398 => to_unsigned(32612, LUT_AMPL_WIDTH - 1),
		17399 => to_unsigned(32612, LUT_AMPL_WIDTH - 1),
		17400 => to_unsigned(32612, LUT_AMPL_WIDTH - 1),
		17401 => to_unsigned(32611, LUT_AMPL_WIDTH - 1),
		17402 => to_unsigned(32611, LUT_AMPL_WIDTH - 1),
		17403 => to_unsigned(32611, LUT_AMPL_WIDTH - 1),
		17404 => to_unsigned(32610, LUT_AMPL_WIDTH - 1),
		17405 => to_unsigned(32610, LUT_AMPL_WIDTH - 1),
		17406 => to_unsigned(32610, LUT_AMPL_WIDTH - 1),
		17407 => to_unsigned(32610, LUT_AMPL_WIDTH - 1),
		17408 => to_unsigned(32609, LUT_AMPL_WIDTH - 1),
		17409 => to_unsigned(32609, LUT_AMPL_WIDTH - 1),
		17410 => to_unsigned(32609, LUT_AMPL_WIDTH - 1),
		17411 => to_unsigned(32608, LUT_AMPL_WIDTH - 1),
		17412 => to_unsigned(32608, LUT_AMPL_WIDTH - 1),
		17413 => to_unsigned(32608, LUT_AMPL_WIDTH - 1),
		17414 => to_unsigned(32607, LUT_AMPL_WIDTH - 1),
		17415 => to_unsigned(32607, LUT_AMPL_WIDTH - 1),
		17416 => to_unsigned(32607, LUT_AMPL_WIDTH - 1),
		17417 => to_unsigned(32606, LUT_AMPL_WIDTH - 1),
		17418 => to_unsigned(32606, LUT_AMPL_WIDTH - 1),
		17419 => to_unsigned(32606, LUT_AMPL_WIDTH - 1),
		17420 => to_unsigned(32606, LUT_AMPL_WIDTH - 1),
		17421 => to_unsigned(32605, LUT_AMPL_WIDTH - 1),
		17422 => to_unsigned(32605, LUT_AMPL_WIDTH - 1),
		17423 => to_unsigned(32605, LUT_AMPL_WIDTH - 1),
		17424 => to_unsigned(32604, LUT_AMPL_WIDTH - 1),
		17425 => to_unsigned(32604, LUT_AMPL_WIDTH - 1),
		17426 => to_unsigned(32604, LUT_AMPL_WIDTH - 1),
		17427 => to_unsigned(32603, LUT_AMPL_WIDTH - 1),
		17428 => to_unsigned(32603, LUT_AMPL_WIDTH - 1),
		17429 => to_unsigned(32603, LUT_AMPL_WIDTH - 1),
		17430 => to_unsigned(32602, LUT_AMPL_WIDTH - 1),
		17431 => to_unsigned(32602, LUT_AMPL_WIDTH - 1),
		17432 => to_unsigned(32602, LUT_AMPL_WIDTH - 1),
		17433 => to_unsigned(32601, LUT_AMPL_WIDTH - 1),
		17434 => to_unsigned(32601, LUT_AMPL_WIDTH - 1),
		17435 => to_unsigned(32601, LUT_AMPL_WIDTH - 1),
		17436 => to_unsigned(32600, LUT_AMPL_WIDTH - 1),
		17437 => to_unsigned(32600, LUT_AMPL_WIDTH - 1),
		17438 => to_unsigned(32600, LUT_AMPL_WIDTH - 1),
		17439 => to_unsigned(32600, LUT_AMPL_WIDTH - 1),
		17440 => to_unsigned(32599, LUT_AMPL_WIDTH - 1),
		17441 => to_unsigned(32599, LUT_AMPL_WIDTH - 1),
		17442 => to_unsigned(32599, LUT_AMPL_WIDTH - 1),
		17443 => to_unsigned(32598, LUT_AMPL_WIDTH - 1),
		17444 => to_unsigned(32598, LUT_AMPL_WIDTH - 1),
		17445 => to_unsigned(32598, LUT_AMPL_WIDTH - 1),
		17446 => to_unsigned(32597, LUT_AMPL_WIDTH - 1),
		17447 => to_unsigned(32597, LUT_AMPL_WIDTH - 1),
		17448 => to_unsigned(32597, LUT_AMPL_WIDTH - 1),
		17449 => to_unsigned(32596, LUT_AMPL_WIDTH - 1),
		17450 => to_unsigned(32596, LUT_AMPL_WIDTH - 1),
		17451 => to_unsigned(32596, LUT_AMPL_WIDTH - 1),
		17452 => to_unsigned(32595, LUT_AMPL_WIDTH - 1),
		17453 => to_unsigned(32595, LUT_AMPL_WIDTH - 1),
		17454 => to_unsigned(32595, LUT_AMPL_WIDTH - 1),
		17455 => to_unsigned(32594, LUT_AMPL_WIDTH - 1),
		17456 => to_unsigned(32594, LUT_AMPL_WIDTH - 1),
		17457 => to_unsigned(32594, LUT_AMPL_WIDTH - 1),
		17458 => to_unsigned(32593, LUT_AMPL_WIDTH - 1),
		17459 => to_unsigned(32593, LUT_AMPL_WIDTH - 1),
		17460 => to_unsigned(32593, LUT_AMPL_WIDTH - 1),
		17461 => to_unsigned(32592, LUT_AMPL_WIDTH - 1),
		17462 => to_unsigned(32592, LUT_AMPL_WIDTH - 1),
		17463 => to_unsigned(32592, LUT_AMPL_WIDTH - 1),
		17464 => to_unsigned(32592, LUT_AMPL_WIDTH - 1),
		17465 => to_unsigned(32591, LUT_AMPL_WIDTH - 1),
		17466 => to_unsigned(32591, LUT_AMPL_WIDTH - 1),
		17467 => to_unsigned(32591, LUT_AMPL_WIDTH - 1),
		17468 => to_unsigned(32590, LUT_AMPL_WIDTH - 1),
		17469 => to_unsigned(32590, LUT_AMPL_WIDTH - 1),
		17470 => to_unsigned(32590, LUT_AMPL_WIDTH - 1),
		17471 => to_unsigned(32589, LUT_AMPL_WIDTH - 1),
		17472 => to_unsigned(32589, LUT_AMPL_WIDTH - 1),
		17473 => to_unsigned(32589, LUT_AMPL_WIDTH - 1),
		17474 => to_unsigned(32588, LUT_AMPL_WIDTH - 1),
		17475 => to_unsigned(32588, LUT_AMPL_WIDTH - 1),
		17476 => to_unsigned(32588, LUT_AMPL_WIDTH - 1),
		17477 => to_unsigned(32587, LUT_AMPL_WIDTH - 1),
		17478 => to_unsigned(32587, LUT_AMPL_WIDTH - 1),
		17479 => to_unsigned(32587, LUT_AMPL_WIDTH - 1),
		17480 => to_unsigned(32586, LUT_AMPL_WIDTH - 1),
		17481 => to_unsigned(32586, LUT_AMPL_WIDTH - 1),
		17482 => to_unsigned(32586, LUT_AMPL_WIDTH - 1),
		17483 => to_unsigned(32585, LUT_AMPL_WIDTH - 1),
		17484 => to_unsigned(32585, LUT_AMPL_WIDTH - 1),
		17485 => to_unsigned(32585, LUT_AMPL_WIDTH - 1),
		17486 => to_unsigned(32584, LUT_AMPL_WIDTH - 1),
		17487 => to_unsigned(32584, LUT_AMPL_WIDTH - 1),
		17488 => to_unsigned(32584, LUT_AMPL_WIDTH - 1),
		17489 => to_unsigned(32583, LUT_AMPL_WIDTH - 1),
		17490 => to_unsigned(32583, LUT_AMPL_WIDTH - 1),
		17491 => to_unsigned(32583, LUT_AMPL_WIDTH - 1),
		17492 => to_unsigned(32582, LUT_AMPL_WIDTH - 1),
		17493 => to_unsigned(32582, LUT_AMPL_WIDTH - 1),
		17494 => to_unsigned(32582, LUT_AMPL_WIDTH - 1),
		17495 => to_unsigned(32581, LUT_AMPL_WIDTH - 1),
		17496 => to_unsigned(32581, LUT_AMPL_WIDTH - 1),
		17497 => to_unsigned(32581, LUT_AMPL_WIDTH - 1),
		17498 => to_unsigned(32580, LUT_AMPL_WIDTH - 1),
		17499 => to_unsigned(32580, LUT_AMPL_WIDTH - 1),
		17500 => to_unsigned(32580, LUT_AMPL_WIDTH - 1),
		17501 => to_unsigned(32579, LUT_AMPL_WIDTH - 1),
		17502 => to_unsigned(32579, LUT_AMPL_WIDTH - 1),
		17503 => to_unsigned(32579, LUT_AMPL_WIDTH - 1),
		17504 => to_unsigned(32578, LUT_AMPL_WIDTH - 1),
		17505 => to_unsigned(32578, LUT_AMPL_WIDTH - 1),
		17506 => to_unsigned(32578, LUT_AMPL_WIDTH - 1),
		17507 => to_unsigned(32577, LUT_AMPL_WIDTH - 1),
		17508 => to_unsigned(32577, LUT_AMPL_WIDTH - 1),
		17509 => to_unsigned(32577, LUT_AMPL_WIDTH - 1),
		17510 => to_unsigned(32576, LUT_AMPL_WIDTH - 1),
		17511 => to_unsigned(32576, LUT_AMPL_WIDTH - 1),
		17512 => to_unsigned(32576, LUT_AMPL_WIDTH - 1),
		17513 => to_unsigned(32575, LUT_AMPL_WIDTH - 1),
		17514 => to_unsigned(32575, LUT_AMPL_WIDTH - 1),
		17515 => to_unsigned(32575, LUT_AMPL_WIDTH - 1),
		17516 => to_unsigned(32574, LUT_AMPL_WIDTH - 1),
		17517 => to_unsigned(32574, LUT_AMPL_WIDTH - 1),
		17518 => to_unsigned(32574, LUT_AMPL_WIDTH - 1),
		17519 => to_unsigned(32573, LUT_AMPL_WIDTH - 1),
		17520 => to_unsigned(32573, LUT_AMPL_WIDTH - 1),
		17521 => to_unsigned(32573, LUT_AMPL_WIDTH - 1),
		17522 => to_unsigned(32572, LUT_AMPL_WIDTH - 1),
		17523 => to_unsigned(32572, LUT_AMPL_WIDTH - 1),
		17524 => to_unsigned(32571, LUT_AMPL_WIDTH - 1),
		17525 => to_unsigned(32571, LUT_AMPL_WIDTH - 1),
		17526 => to_unsigned(32571, LUT_AMPL_WIDTH - 1),
		17527 => to_unsigned(32570, LUT_AMPL_WIDTH - 1),
		17528 => to_unsigned(32570, LUT_AMPL_WIDTH - 1),
		17529 => to_unsigned(32570, LUT_AMPL_WIDTH - 1),
		17530 => to_unsigned(32569, LUT_AMPL_WIDTH - 1),
		17531 => to_unsigned(32569, LUT_AMPL_WIDTH - 1),
		17532 => to_unsigned(32569, LUT_AMPL_WIDTH - 1),
		17533 => to_unsigned(32568, LUT_AMPL_WIDTH - 1),
		17534 => to_unsigned(32568, LUT_AMPL_WIDTH - 1),
		17535 => to_unsigned(32568, LUT_AMPL_WIDTH - 1),
		17536 => to_unsigned(32567, LUT_AMPL_WIDTH - 1),
		17537 => to_unsigned(32567, LUT_AMPL_WIDTH - 1),
		17538 => to_unsigned(32567, LUT_AMPL_WIDTH - 1),
		17539 => to_unsigned(32566, LUT_AMPL_WIDTH - 1),
		17540 => to_unsigned(32566, LUT_AMPL_WIDTH - 1),
		17541 => to_unsigned(32566, LUT_AMPL_WIDTH - 1),
		17542 => to_unsigned(32565, LUT_AMPL_WIDTH - 1),
		17543 => to_unsigned(32565, LUT_AMPL_WIDTH - 1),
		17544 => to_unsigned(32565, LUT_AMPL_WIDTH - 1),
		17545 => to_unsigned(32564, LUT_AMPL_WIDTH - 1),
		17546 => to_unsigned(32564, LUT_AMPL_WIDTH - 1),
		17547 => to_unsigned(32564, LUT_AMPL_WIDTH - 1),
		17548 => to_unsigned(32563, LUT_AMPL_WIDTH - 1),
		17549 => to_unsigned(32563, LUT_AMPL_WIDTH - 1),
		17550 => to_unsigned(32562, LUT_AMPL_WIDTH - 1),
		17551 => to_unsigned(32562, LUT_AMPL_WIDTH - 1),
		17552 => to_unsigned(32562, LUT_AMPL_WIDTH - 1),
		17553 => to_unsigned(32561, LUT_AMPL_WIDTH - 1),
		17554 => to_unsigned(32561, LUT_AMPL_WIDTH - 1),
		17555 => to_unsigned(32561, LUT_AMPL_WIDTH - 1),
		17556 => to_unsigned(32560, LUT_AMPL_WIDTH - 1),
		17557 => to_unsigned(32560, LUT_AMPL_WIDTH - 1),
		17558 => to_unsigned(32560, LUT_AMPL_WIDTH - 1),
		17559 => to_unsigned(32559, LUT_AMPL_WIDTH - 1),
		17560 => to_unsigned(32559, LUT_AMPL_WIDTH - 1),
		17561 => to_unsigned(32559, LUT_AMPL_WIDTH - 1),
		17562 => to_unsigned(32558, LUT_AMPL_WIDTH - 1),
		17563 => to_unsigned(32558, LUT_AMPL_WIDTH - 1),
		17564 => to_unsigned(32558, LUT_AMPL_WIDTH - 1),
		17565 => to_unsigned(32557, LUT_AMPL_WIDTH - 1),
		17566 => to_unsigned(32557, LUT_AMPL_WIDTH - 1),
		17567 => to_unsigned(32556, LUT_AMPL_WIDTH - 1),
		17568 => to_unsigned(32556, LUT_AMPL_WIDTH - 1),
		17569 => to_unsigned(32556, LUT_AMPL_WIDTH - 1),
		17570 => to_unsigned(32555, LUT_AMPL_WIDTH - 1),
		17571 => to_unsigned(32555, LUT_AMPL_WIDTH - 1),
		17572 => to_unsigned(32555, LUT_AMPL_WIDTH - 1),
		17573 => to_unsigned(32554, LUT_AMPL_WIDTH - 1),
		17574 => to_unsigned(32554, LUT_AMPL_WIDTH - 1),
		17575 => to_unsigned(32554, LUT_AMPL_WIDTH - 1),
		17576 => to_unsigned(32553, LUT_AMPL_WIDTH - 1),
		17577 => to_unsigned(32553, LUT_AMPL_WIDTH - 1),
		17578 => to_unsigned(32553, LUT_AMPL_WIDTH - 1),
		17579 => to_unsigned(32552, LUT_AMPL_WIDTH - 1),
		17580 => to_unsigned(32552, LUT_AMPL_WIDTH - 1),
		17581 => to_unsigned(32551, LUT_AMPL_WIDTH - 1),
		17582 => to_unsigned(32551, LUT_AMPL_WIDTH - 1),
		17583 => to_unsigned(32551, LUT_AMPL_WIDTH - 1),
		17584 => to_unsigned(32550, LUT_AMPL_WIDTH - 1),
		17585 => to_unsigned(32550, LUT_AMPL_WIDTH - 1),
		17586 => to_unsigned(32550, LUT_AMPL_WIDTH - 1),
		17587 => to_unsigned(32549, LUT_AMPL_WIDTH - 1),
		17588 => to_unsigned(32549, LUT_AMPL_WIDTH - 1),
		17589 => to_unsigned(32549, LUT_AMPL_WIDTH - 1),
		17590 => to_unsigned(32548, LUT_AMPL_WIDTH - 1),
		17591 => to_unsigned(32548, LUT_AMPL_WIDTH - 1),
		17592 => to_unsigned(32547, LUT_AMPL_WIDTH - 1),
		17593 => to_unsigned(32547, LUT_AMPL_WIDTH - 1),
		17594 => to_unsigned(32547, LUT_AMPL_WIDTH - 1),
		17595 => to_unsigned(32546, LUT_AMPL_WIDTH - 1),
		17596 => to_unsigned(32546, LUT_AMPL_WIDTH - 1),
		17597 => to_unsigned(32546, LUT_AMPL_WIDTH - 1),
		17598 => to_unsigned(32545, LUT_AMPL_WIDTH - 1),
		17599 => to_unsigned(32545, LUT_AMPL_WIDTH - 1),
		17600 => to_unsigned(32545, LUT_AMPL_WIDTH - 1),
		17601 => to_unsigned(32544, LUT_AMPL_WIDTH - 1),
		17602 => to_unsigned(32544, LUT_AMPL_WIDTH - 1),
		17603 => to_unsigned(32543, LUT_AMPL_WIDTH - 1),
		17604 => to_unsigned(32543, LUT_AMPL_WIDTH - 1),
		17605 => to_unsigned(32543, LUT_AMPL_WIDTH - 1),
		17606 => to_unsigned(32542, LUT_AMPL_WIDTH - 1),
		17607 => to_unsigned(32542, LUT_AMPL_WIDTH - 1),
		17608 => to_unsigned(32542, LUT_AMPL_WIDTH - 1),
		17609 => to_unsigned(32541, LUT_AMPL_WIDTH - 1),
		17610 => to_unsigned(32541, LUT_AMPL_WIDTH - 1),
		17611 => to_unsigned(32541, LUT_AMPL_WIDTH - 1),
		17612 => to_unsigned(32540, LUT_AMPL_WIDTH - 1),
		17613 => to_unsigned(32540, LUT_AMPL_WIDTH - 1),
		17614 => to_unsigned(32539, LUT_AMPL_WIDTH - 1),
		17615 => to_unsigned(32539, LUT_AMPL_WIDTH - 1),
		17616 => to_unsigned(32539, LUT_AMPL_WIDTH - 1),
		17617 => to_unsigned(32538, LUT_AMPL_WIDTH - 1),
		17618 => to_unsigned(32538, LUT_AMPL_WIDTH - 1),
		17619 => to_unsigned(32538, LUT_AMPL_WIDTH - 1),
		17620 => to_unsigned(32537, LUT_AMPL_WIDTH - 1),
		17621 => to_unsigned(32537, LUT_AMPL_WIDTH - 1),
		17622 => to_unsigned(32536, LUT_AMPL_WIDTH - 1),
		17623 => to_unsigned(32536, LUT_AMPL_WIDTH - 1),
		17624 => to_unsigned(32536, LUT_AMPL_WIDTH - 1),
		17625 => to_unsigned(32535, LUT_AMPL_WIDTH - 1),
		17626 => to_unsigned(32535, LUT_AMPL_WIDTH - 1),
		17627 => to_unsigned(32535, LUT_AMPL_WIDTH - 1),
		17628 => to_unsigned(32534, LUT_AMPL_WIDTH - 1),
		17629 => to_unsigned(32534, LUT_AMPL_WIDTH - 1),
		17630 => to_unsigned(32533, LUT_AMPL_WIDTH - 1),
		17631 => to_unsigned(32533, LUT_AMPL_WIDTH - 1),
		17632 => to_unsigned(32533, LUT_AMPL_WIDTH - 1),
		17633 => to_unsigned(32532, LUT_AMPL_WIDTH - 1),
		17634 => to_unsigned(32532, LUT_AMPL_WIDTH - 1),
		17635 => to_unsigned(32532, LUT_AMPL_WIDTH - 1),
		17636 => to_unsigned(32531, LUT_AMPL_WIDTH - 1),
		17637 => to_unsigned(32531, LUT_AMPL_WIDTH - 1),
		17638 => to_unsigned(32530, LUT_AMPL_WIDTH - 1),
		17639 => to_unsigned(32530, LUT_AMPL_WIDTH - 1),
		17640 => to_unsigned(32530, LUT_AMPL_WIDTH - 1),
		17641 => to_unsigned(32529, LUT_AMPL_WIDTH - 1),
		17642 => to_unsigned(32529, LUT_AMPL_WIDTH - 1),
		17643 => to_unsigned(32529, LUT_AMPL_WIDTH - 1),
		17644 => to_unsigned(32528, LUT_AMPL_WIDTH - 1),
		17645 => to_unsigned(32528, LUT_AMPL_WIDTH - 1),
		17646 => to_unsigned(32527, LUT_AMPL_WIDTH - 1),
		17647 => to_unsigned(32527, LUT_AMPL_WIDTH - 1),
		17648 => to_unsigned(32527, LUT_AMPL_WIDTH - 1),
		17649 => to_unsigned(32526, LUT_AMPL_WIDTH - 1),
		17650 => to_unsigned(32526, LUT_AMPL_WIDTH - 1),
		17651 => to_unsigned(32526, LUT_AMPL_WIDTH - 1),
		17652 => to_unsigned(32525, LUT_AMPL_WIDTH - 1),
		17653 => to_unsigned(32525, LUT_AMPL_WIDTH - 1),
		17654 => to_unsigned(32524, LUT_AMPL_WIDTH - 1),
		17655 => to_unsigned(32524, LUT_AMPL_WIDTH - 1),
		17656 => to_unsigned(32524, LUT_AMPL_WIDTH - 1),
		17657 => to_unsigned(32523, LUT_AMPL_WIDTH - 1),
		17658 => to_unsigned(32523, LUT_AMPL_WIDTH - 1),
		17659 => to_unsigned(32522, LUT_AMPL_WIDTH - 1),
		17660 => to_unsigned(32522, LUT_AMPL_WIDTH - 1),
		17661 => to_unsigned(32522, LUT_AMPL_WIDTH - 1),
		17662 => to_unsigned(32521, LUT_AMPL_WIDTH - 1),
		17663 => to_unsigned(32521, LUT_AMPL_WIDTH - 1),
		17664 => to_unsigned(32521, LUT_AMPL_WIDTH - 1),
		17665 => to_unsigned(32520, LUT_AMPL_WIDTH - 1),
		17666 => to_unsigned(32520, LUT_AMPL_WIDTH - 1),
		17667 => to_unsigned(32519, LUT_AMPL_WIDTH - 1),
		17668 => to_unsigned(32519, LUT_AMPL_WIDTH - 1),
		17669 => to_unsigned(32519, LUT_AMPL_WIDTH - 1),
		17670 => to_unsigned(32518, LUT_AMPL_WIDTH - 1),
		17671 => to_unsigned(32518, LUT_AMPL_WIDTH - 1),
		17672 => to_unsigned(32517, LUT_AMPL_WIDTH - 1),
		17673 => to_unsigned(32517, LUT_AMPL_WIDTH - 1),
		17674 => to_unsigned(32517, LUT_AMPL_WIDTH - 1),
		17675 => to_unsigned(32516, LUT_AMPL_WIDTH - 1),
		17676 => to_unsigned(32516, LUT_AMPL_WIDTH - 1),
		17677 => to_unsigned(32516, LUT_AMPL_WIDTH - 1),
		17678 => to_unsigned(32515, LUT_AMPL_WIDTH - 1),
		17679 => to_unsigned(32515, LUT_AMPL_WIDTH - 1),
		17680 => to_unsigned(32514, LUT_AMPL_WIDTH - 1),
		17681 => to_unsigned(32514, LUT_AMPL_WIDTH - 1),
		17682 => to_unsigned(32514, LUT_AMPL_WIDTH - 1),
		17683 => to_unsigned(32513, LUT_AMPL_WIDTH - 1),
		17684 => to_unsigned(32513, LUT_AMPL_WIDTH - 1),
		17685 => to_unsigned(32512, LUT_AMPL_WIDTH - 1),
		17686 => to_unsigned(32512, LUT_AMPL_WIDTH - 1),
		17687 => to_unsigned(32512, LUT_AMPL_WIDTH - 1),
		17688 => to_unsigned(32511, LUT_AMPL_WIDTH - 1),
		17689 => to_unsigned(32511, LUT_AMPL_WIDTH - 1),
		17690 => to_unsigned(32510, LUT_AMPL_WIDTH - 1),
		17691 => to_unsigned(32510, LUT_AMPL_WIDTH - 1),
		17692 => to_unsigned(32510, LUT_AMPL_WIDTH - 1),
		17693 => to_unsigned(32509, LUT_AMPL_WIDTH - 1),
		17694 => to_unsigned(32509, LUT_AMPL_WIDTH - 1),
		17695 => to_unsigned(32509, LUT_AMPL_WIDTH - 1),
		17696 => to_unsigned(32508, LUT_AMPL_WIDTH - 1),
		17697 => to_unsigned(32508, LUT_AMPL_WIDTH - 1),
		17698 => to_unsigned(32507, LUT_AMPL_WIDTH - 1),
		17699 => to_unsigned(32507, LUT_AMPL_WIDTH - 1),
		17700 => to_unsigned(32507, LUT_AMPL_WIDTH - 1),
		17701 => to_unsigned(32506, LUT_AMPL_WIDTH - 1),
		17702 => to_unsigned(32506, LUT_AMPL_WIDTH - 1),
		17703 => to_unsigned(32505, LUT_AMPL_WIDTH - 1),
		17704 => to_unsigned(32505, LUT_AMPL_WIDTH - 1),
		17705 => to_unsigned(32505, LUT_AMPL_WIDTH - 1),
		17706 => to_unsigned(32504, LUT_AMPL_WIDTH - 1),
		17707 => to_unsigned(32504, LUT_AMPL_WIDTH - 1),
		17708 => to_unsigned(32503, LUT_AMPL_WIDTH - 1),
		17709 => to_unsigned(32503, LUT_AMPL_WIDTH - 1),
		17710 => to_unsigned(32503, LUT_AMPL_WIDTH - 1),
		17711 => to_unsigned(32502, LUT_AMPL_WIDTH - 1),
		17712 => to_unsigned(32502, LUT_AMPL_WIDTH - 1),
		17713 => to_unsigned(32501, LUT_AMPL_WIDTH - 1),
		17714 => to_unsigned(32501, LUT_AMPL_WIDTH - 1),
		17715 => to_unsigned(32501, LUT_AMPL_WIDTH - 1),
		17716 => to_unsigned(32500, LUT_AMPL_WIDTH - 1),
		17717 => to_unsigned(32500, LUT_AMPL_WIDTH - 1),
		17718 => to_unsigned(32499, LUT_AMPL_WIDTH - 1),
		17719 => to_unsigned(32499, LUT_AMPL_WIDTH - 1),
		17720 => to_unsigned(32499, LUT_AMPL_WIDTH - 1),
		17721 => to_unsigned(32498, LUT_AMPL_WIDTH - 1),
		17722 => to_unsigned(32498, LUT_AMPL_WIDTH - 1),
		17723 => to_unsigned(32497, LUT_AMPL_WIDTH - 1),
		17724 => to_unsigned(32497, LUT_AMPL_WIDTH - 1),
		17725 => to_unsigned(32497, LUT_AMPL_WIDTH - 1),
		17726 => to_unsigned(32496, LUT_AMPL_WIDTH - 1),
		17727 => to_unsigned(32496, LUT_AMPL_WIDTH - 1),
		17728 => to_unsigned(32495, LUT_AMPL_WIDTH - 1),
		17729 => to_unsigned(32495, LUT_AMPL_WIDTH - 1),
		17730 => to_unsigned(32495, LUT_AMPL_WIDTH - 1),
		17731 => to_unsigned(32494, LUT_AMPL_WIDTH - 1),
		17732 => to_unsigned(32494, LUT_AMPL_WIDTH - 1),
		17733 => to_unsigned(32493, LUT_AMPL_WIDTH - 1),
		17734 => to_unsigned(32493, LUT_AMPL_WIDTH - 1),
		17735 => to_unsigned(32493, LUT_AMPL_WIDTH - 1),
		17736 => to_unsigned(32492, LUT_AMPL_WIDTH - 1),
		17737 => to_unsigned(32492, LUT_AMPL_WIDTH - 1),
		17738 => to_unsigned(32491, LUT_AMPL_WIDTH - 1),
		17739 => to_unsigned(32491, LUT_AMPL_WIDTH - 1),
		17740 => to_unsigned(32490, LUT_AMPL_WIDTH - 1),
		17741 => to_unsigned(32490, LUT_AMPL_WIDTH - 1),
		17742 => to_unsigned(32490, LUT_AMPL_WIDTH - 1),
		17743 => to_unsigned(32489, LUT_AMPL_WIDTH - 1),
		17744 => to_unsigned(32489, LUT_AMPL_WIDTH - 1),
		17745 => to_unsigned(32488, LUT_AMPL_WIDTH - 1),
		17746 => to_unsigned(32488, LUT_AMPL_WIDTH - 1),
		17747 => to_unsigned(32488, LUT_AMPL_WIDTH - 1),
		17748 => to_unsigned(32487, LUT_AMPL_WIDTH - 1),
		17749 => to_unsigned(32487, LUT_AMPL_WIDTH - 1),
		17750 => to_unsigned(32486, LUT_AMPL_WIDTH - 1),
		17751 => to_unsigned(32486, LUT_AMPL_WIDTH - 1),
		17752 => to_unsigned(32486, LUT_AMPL_WIDTH - 1),
		17753 => to_unsigned(32485, LUT_AMPL_WIDTH - 1),
		17754 => to_unsigned(32485, LUT_AMPL_WIDTH - 1),
		17755 => to_unsigned(32484, LUT_AMPL_WIDTH - 1),
		17756 => to_unsigned(32484, LUT_AMPL_WIDTH - 1),
		17757 => to_unsigned(32484, LUT_AMPL_WIDTH - 1),
		17758 => to_unsigned(32483, LUT_AMPL_WIDTH - 1),
		17759 => to_unsigned(32483, LUT_AMPL_WIDTH - 1),
		17760 => to_unsigned(32482, LUT_AMPL_WIDTH - 1),
		17761 => to_unsigned(32482, LUT_AMPL_WIDTH - 1),
		17762 => to_unsigned(32481, LUT_AMPL_WIDTH - 1),
		17763 => to_unsigned(32481, LUT_AMPL_WIDTH - 1),
		17764 => to_unsigned(32481, LUT_AMPL_WIDTH - 1),
		17765 => to_unsigned(32480, LUT_AMPL_WIDTH - 1),
		17766 => to_unsigned(32480, LUT_AMPL_WIDTH - 1),
		17767 => to_unsigned(32479, LUT_AMPL_WIDTH - 1),
		17768 => to_unsigned(32479, LUT_AMPL_WIDTH - 1),
		17769 => to_unsigned(32479, LUT_AMPL_WIDTH - 1),
		17770 => to_unsigned(32478, LUT_AMPL_WIDTH - 1),
		17771 => to_unsigned(32478, LUT_AMPL_WIDTH - 1),
		17772 => to_unsigned(32477, LUT_AMPL_WIDTH - 1),
		17773 => to_unsigned(32477, LUT_AMPL_WIDTH - 1),
		17774 => to_unsigned(32476, LUT_AMPL_WIDTH - 1),
		17775 => to_unsigned(32476, LUT_AMPL_WIDTH - 1),
		17776 => to_unsigned(32476, LUT_AMPL_WIDTH - 1),
		17777 => to_unsigned(32475, LUT_AMPL_WIDTH - 1),
		17778 => to_unsigned(32475, LUT_AMPL_WIDTH - 1),
		17779 => to_unsigned(32474, LUT_AMPL_WIDTH - 1),
		17780 => to_unsigned(32474, LUT_AMPL_WIDTH - 1),
		17781 => to_unsigned(32474, LUT_AMPL_WIDTH - 1),
		17782 => to_unsigned(32473, LUT_AMPL_WIDTH - 1),
		17783 => to_unsigned(32473, LUT_AMPL_WIDTH - 1),
		17784 => to_unsigned(32472, LUT_AMPL_WIDTH - 1),
		17785 => to_unsigned(32472, LUT_AMPL_WIDTH - 1),
		17786 => to_unsigned(32471, LUT_AMPL_WIDTH - 1),
		17787 => to_unsigned(32471, LUT_AMPL_WIDTH - 1),
		17788 => to_unsigned(32471, LUT_AMPL_WIDTH - 1),
		17789 => to_unsigned(32470, LUT_AMPL_WIDTH - 1),
		17790 => to_unsigned(32470, LUT_AMPL_WIDTH - 1),
		17791 => to_unsigned(32469, LUT_AMPL_WIDTH - 1),
		17792 => to_unsigned(32469, LUT_AMPL_WIDTH - 1),
		17793 => to_unsigned(32468, LUT_AMPL_WIDTH - 1),
		17794 => to_unsigned(32468, LUT_AMPL_WIDTH - 1),
		17795 => to_unsigned(32468, LUT_AMPL_WIDTH - 1),
		17796 => to_unsigned(32467, LUT_AMPL_WIDTH - 1),
		17797 => to_unsigned(32467, LUT_AMPL_WIDTH - 1),
		17798 => to_unsigned(32466, LUT_AMPL_WIDTH - 1),
		17799 => to_unsigned(32466, LUT_AMPL_WIDTH - 1),
		17800 => to_unsigned(32466, LUT_AMPL_WIDTH - 1),
		17801 => to_unsigned(32465, LUT_AMPL_WIDTH - 1),
		17802 => to_unsigned(32465, LUT_AMPL_WIDTH - 1),
		17803 => to_unsigned(32464, LUT_AMPL_WIDTH - 1),
		17804 => to_unsigned(32464, LUT_AMPL_WIDTH - 1),
		17805 => to_unsigned(32463, LUT_AMPL_WIDTH - 1),
		17806 => to_unsigned(32463, LUT_AMPL_WIDTH - 1),
		17807 => to_unsigned(32463, LUT_AMPL_WIDTH - 1),
		17808 => to_unsigned(32462, LUT_AMPL_WIDTH - 1),
		17809 => to_unsigned(32462, LUT_AMPL_WIDTH - 1),
		17810 => to_unsigned(32461, LUT_AMPL_WIDTH - 1),
		17811 => to_unsigned(32461, LUT_AMPL_WIDTH - 1),
		17812 => to_unsigned(32460, LUT_AMPL_WIDTH - 1),
		17813 => to_unsigned(32460, LUT_AMPL_WIDTH - 1),
		17814 => to_unsigned(32460, LUT_AMPL_WIDTH - 1),
		17815 => to_unsigned(32459, LUT_AMPL_WIDTH - 1),
		17816 => to_unsigned(32459, LUT_AMPL_WIDTH - 1),
		17817 => to_unsigned(32458, LUT_AMPL_WIDTH - 1),
		17818 => to_unsigned(32458, LUT_AMPL_WIDTH - 1),
		17819 => to_unsigned(32457, LUT_AMPL_WIDTH - 1),
		17820 => to_unsigned(32457, LUT_AMPL_WIDTH - 1),
		17821 => to_unsigned(32457, LUT_AMPL_WIDTH - 1),
		17822 => to_unsigned(32456, LUT_AMPL_WIDTH - 1),
		17823 => to_unsigned(32456, LUT_AMPL_WIDTH - 1),
		17824 => to_unsigned(32455, LUT_AMPL_WIDTH - 1),
		17825 => to_unsigned(32455, LUT_AMPL_WIDTH - 1),
		17826 => to_unsigned(32454, LUT_AMPL_WIDTH - 1),
		17827 => to_unsigned(32454, LUT_AMPL_WIDTH - 1),
		17828 => to_unsigned(32453, LUT_AMPL_WIDTH - 1),
		17829 => to_unsigned(32453, LUT_AMPL_WIDTH - 1),
		17830 => to_unsigned(32453, LUT_AMPL_WIDTH - 1),
		17831 => to_unsigned(32452, LUT_AMPL_WIDTH - 1),
		17832 => to_unsigned(32452, LUT_AMPL_WIDTH - 1),
		17833 => to_unsigned(32451, LUT_AMPL_WIDTH - 1),
		17834 => to_unsigned(32451, LUT_AMPL_WIDTH - 1),
		17835 => to_unsigned(32450, LUT_AMPL_WIDTH - 1),
		17836 => to_unsigned(32450, LUT_AMPL_WIDTH - 1),
		17837 => to_unsigned(32450, LUT_AMPL_WIDTH - 1),
		17838 => to_unsigned(32449, LUT_AMPL_WIDTH - 1),
		17839 => to_unsigned(32449, LUT_AMPL_WIDTH - 1),
		17840 => to_unsigned(32448, LUT_AMPL_WIDTH - 1),
		17841 => to_unsigned(32448, LUT_AMPL_WIDTH - 1),
		17842 => to_unsigned(32447, LUT_AMPL_WIDTH - 1),
		17843 => to_unsigned(32447, LUT_AMPL_WIDTH - 1),
		17844 => to_unsigned(32447, LUT_AMPL_WIDTH - 1),
		17845 => to_unsigned(32446, LUT_AMPL_WIDTH - 1),
		17846 => to_unsigned(32446, LUT_AMPL_WIDTH - 1),
		17847 => to_unsigned(32445, LUT_AMPL_WIDTH - 1),
		17848 => to_unsigned(32445, LUT_AMPL_WIDTH - 1),
		17849 => to_unsigned(32444, LUT_AMPL_WIDTH - 1),
		17850 => to_unsigned(32444, LUT_AMPL_WIDTH - 1),
		17851 => to_unsigned(32443, LUT_AMPL_WIDTH - 1),
		17852 => to_unsigned(32443, LUT_AMPL_WIDTH - 1),
		17853 => to_unsigned(32443, LUT_AMPL_WIDTH - 1),
		17854 => to_unsigned(32442, LUT_AMPL_WIDTH - 1),
		17855 => to_unsigned(32442, LUT_AMPL_WIDTH - 1),
		17856 => to_unsigned(32441, LUT_AMPL_WIDTH - 1),
		17857 => to_unsigned(32441, LUT_AMPL_WIDTH - 1),
		17858 => to_unsigned(32440, LUT_AMPL_WIDTH - 1),
		17859 => to_unsigned(32440, LUT_AMPL_WIDTH - 1),
		17860 => to_unsigned(32439, LUT_AMPL_WIDTH - 1),
		17861 => to_unsigned(32439, LUT_AMPL_WIDTH - 1),
		17862 => to_unsigned(32439, LUT_AMPL_WIDTH - 1),
		17863 => to_unsigned(32438, LUT_AMPL_WIDTH - 1),
		17864 => to_unsigned(32438, LUT_AMPL_WIDTH - 1),
		17865 => to_unsigned(32437, LUT_AMPL_WIDTH - 1),
		17866 => to_unsigned(32437, LUT_AMPL_WIDTH - 1),
		17867 => to_unsigned(32436, LUT_AMPL_WIDTH - 1),
		17868 => to_unsigned(32436, LUT_AMPL_WIDTH - 1),
		17869 => to_unsigned(32435, LUT_AMPL_WIDTH - 1),
		17870 => to_unsigned(32435, LUT_AMPL_WIDTH - 1),
		17871 => to_unsigned(32435, LUT_AMPL_WIDTH - 1),
		17872 => to_unsigned(32434, LUT_AMPL_WIDTH - 1),
		17873 => to_unsigned(32434, LUT_AMPL_WIDTH - 1),
		17874 => to_unsigned(32433, LUT_AMPL_WIDTH - 1),
		17875 => to_unsigned(32433, LUT_AMPL_WIDTH - 1),
		17876 => to_unsigned(32432, LUT_AMPL_WIDTH - 1),
		17877 => to_unsigned(32432, LUT_AMPL_WIDTH - 1),
		17878 => to_unsigned(32431, LUT_AMPL_WIDTH - 1),
		17879 => to_unsigned(32431, LUT_AMPL_WIDTH - 1),
		17880 => to_unsigned(32431, LUT_AMPL_WIDTH - 1),
		17881 => to_unsigned(32430, LUT_AMPL_WIDTH - 1),
		17882 => to_unsigned(32430, LUT_AMPL_WIDTH - 1),
		17883 => to_unsigned(32429, LUT_AMPL_WIDTH - 1),
		17884 => to_unsigned(32429, LUT_AMPL_WIDTH - 1),
		17885 => to_unsigned(32428, LUT_AMPL_WIDTH - 1),
		17886 => to_unsigned(32428, LUT_AMPL_WIDTH - 1),
		17887 => to_unsigned(32427, LUT_AMPL_WIDTH - 1),
		17888 => to_unsigned(32427, LUT_AMPL_WIDTH - 1),
		17889 => to_unsigned(32426, LUT_AMPL_WIDTH - 1),
		17890 => to_unsigned(32426, LUT_AMPL_WIDTH - 1),
		17891 => to_unsigned(32426, LUT_AMPL_WIDTH - 1),
		17892 => to_unsigned(32425, LUT_AMPL_WIDTH - 1),
		17893 => to_unsigned(32425, LUT_AMPL_WIDTH - 1),
		17894 => to_unsigned(32424, LUT_AMPL_WIDTH - 1),
		17895 => to_unsigned(32424, LUT_AMPL_WIDTH - 1),
		17896 => to_unsigned(32423, LUT_AMPL_WIDTH - 1),
		17897 => to_unsigned(32423, LUT_AMPL_WIDTH - 1),
		17898 => to_unsigned(32422, LUT_AMPL_WIDTH - 1),
		17899 => to_unsigned(32422, LUT_AMPL_WIDTH - 1),
		17900 => to_unsigned(32422, LUT_AMPL_WIDTH - 1),
		17901 => to_unsigned(32421, LUT_AMPL_WIDTH - 1),
		17902 => to_unsigned(32421, LUT_AMPL_WIDTH - 1),
		17903 => to_unsigned(32420, LUT_AMPL_WIDTH - 1),
		17904 => to_unsigned(32420, LUT_AMPL_WIDTH - 1),
		17905 => to_unsigned(32419, LUT_AMPL_WIDTH - 1),
		17906 => to_unsigned(32419, LUT_AMPL_WIDTH - 1),
		17907 => to_unsigned(32418, LUT_AMPL_WIDTH - 1),
		17908 => to_unsigned(32418, LUT_AMPL_WIDTH - 1),
		17909 => to_unsigned(32417, LUT_AMPL_WIDTH - 1),
		17910 => to_unsigned(32417, LUT_AMPL_WIDTH - 1),
		17911 => to_unsigned(32416, LUT_AMPL_WIDTH - 1),
		17912 => to_unsigned(32416, LUT_AMPL_WIDTH - 1),
		17913 => to_unsigned(32416, LUT_AMPL_WIDTH - 1),
		17914 => to_unsigned(32415, LUT_AMPL_WIDTH - 1),
		17915 => to_unsigned(32415, LUT_AMPL_WIDTH - 1),
		17916 => to_unsigned(32414, LUT_AMPL_WIDTH - 1),
		17917 => to_unsigned(32414, LUT_AMPL_WIDTH - 1),
		17918 => to_unsigned(32413, LUT_AMPL_WIDTH - 1),
		17919 => to_unsigned(32413, LUT_AMPL_WIDTH - 1),
		17920 => to_unsigned(32412, LUT_AMPL_WIDTH - 1),
		17921 => to_unsigned(32412, LUT_AMPL_WIDTH - 1),
		17922 => to_unsigned(32411, LUT_AMPL_WIDTH - 1),
		17923 => to_unsigned(32411, LUT_AMPL_WIDTH - 1),
		17924 => to_unsigned(32411, LUT_AMPL_WIDTH - 1),
		17925 => to_unsigned(32410, LUT_AMPL_WIDTH - 1),
		17926 => to_unsigned(32410, LUT_AMPL_WIDTH - 1),
		17927 => to_unsigned(32409, LUT_AMPL_WIDTH - 1),
		17928 => to_unsigned(32409, LUT_AMPL_WIDTH - 1),
		17929 => to_unsigned(32408, LUT_AMPL_WIDTH - 1),
		17930 => to_unsigned(32408, LUT_AMPL_WIDTH - 1),
		17931 => to_unsigned(32407, LUT_AMPL_WIDTH - 1),
		17932 => to_unsigned(32407, LUT_AMPL_WIDTH - 1),
		17933 => to_unsigned(32406, LUT_AMPL_WIDTH - 1),
		17934 => to_unsigned(32406, LUT_AMPL_WIDTH - 1),
		17935 => to_unsigned(32405, LUT_AMPL_WIDTH - 1),
		17936 => to_unsigned(32405, LUT_AMPL_WIDTH - 1),
		17937 => to_unsigned(32404, LUT_AMPL_WIDTH - 1),
		17938 => to_unsigned(32404, LUT_AMPL_WIDTH - 1),
		17939 => to_unsigned(32404, LUT_AMPL_WIDTH - 1),
		17940 => to_unsigned(32403, LUT_AMPL_WIDTH - 1),
		17941 => to_unsigned(32403, LUT_AMPL_WIDTH - 1),
		17942 => to_unsigned(32402, LUT_AMPL_WIDTH - 1),
		17943 => to_unsigned(32402, LUT_AMPL_WIDTH - 1),
		17944 => to_unsigned(32401, LUT_AMPL_WIDTH - 1),
		17945 => to_unsigned(32401, LUT_AMPL_WIDTH - 1),
		17946 => to_unsigned(32400, LUT_AMPL_WIDTH - 1),
		17947 => to_unsigned(32400, LUT_AMPL_WIDTH - 1),
		17948 => to_unsigned(32399, LUT_AMPL_WIDTH - 1),
		17949 => to_unsigned(32399, LUT_AMPL_WIDTH - 1),
		17950 => to_unsigned(32398, LUT_AMPL_WIDTH - 1),
		17951 => to_unsigned(32398, LUT_AMPL_WIDTH - 1),
		17952 => to_unsigned(32397, LUT_AMPL_WIDTH - 1),
		17953 => to_unsigned(32397, LUT_AMPL_WIDTH - 1),
		17954 => to_unsigned(32397, LUT_AMPL_WIDTH - 1),
		17955 => to_unsigned(32396, LUT_AMPL_WIDTH - 1),
		17956 => to_unsigned(32396, LUT_AMPL_WIDTH - 1),
		17957 => to_unsigned(32395, LUT_AMPL_WIDTH - 1),
		17958 => to_unsigned(32395, LUT_AMPL_WIDTH - 1),
		17959 => to_unsigned(32394, LUT_AMPL_WIDTH - 1),
		17960 => to_unsigned(32394, LUT_AMPL_WIDTH - 1),
		17961 => to_unsigned(32393, LUT_AMPL_WIDTH - 1),
		17962 => to_unsigned(32393, LUT_AMPL_WIDTH - 1),
		17963 => to_unsigned(32392, LUT_AMPL_WIDTH - 1),
		17964 => to_unsigned(32392, LUT_AMPL_WIDTH - 1),
		17965 => to_unsigned(32391, LUT_AMPL_WIDTH - 1),
		17966 => to_unsigned(32391, LUT_AMPL_WIDTH - 1),
		17967 => to_unsigned(32390, LUT_AMPL_WIDTH - 1),
		17968 => to_unsigned(32390, LUT_AMPL_WIDTH - 1),
		17969 => to_unsigned(32389, LUT_AMPL_WIDTH - 1),
		17970 => to_unsigned(32389, LUT_AMPL_WIDTH - 1),
		17971 => to_unsigned(32388, LUT_AMPL_WIDTH - 1),
		17972 => to_unsigned(32388, LUT_AMPL_WIDTH - 1),
		17973 => to_unsigned(32387, LUT_AMPL_WIDTH - 1),
		17974 => to_unsigned(32387, LUT_AMPL_WIDTH - 1),
		17975 => to_unsigned(32387, LUT_AMPL_WIDTH - 1),
		17976 => to_unsigned(32386, LUT_AMPL_WIDTH - 1),
		17977 => to_unsigned(32386, LUT_AMPL_WIDTH - 1),
		17978 => to_unsigned(32385, LUT_AMPL_WIDTH - 1),
		17979 => to_unsigned(32385, LUT_AMPL_WIDTH - 1),
		17980 => to_unsigned(32384, LUT_AMPL_WIDTH - 1),
		17981 => to_unsigned(32384, LUT_AMPL_WIDTH - 1),
		17982 => to_unsigned(32383, LUT_AMPL_WIDTH - 1),
		17983 => to_unsigned(32383, LUT_AMPL_WIDTH - 1),
		17984 => to_unsigned(32382, LUT_AMPL_WIDTH - 1),
		17985 => to_unsigned(32382, LUT_AMPL_WIDTH - 1),
		17986 => to_unsigned(32381, LUT_AMPL_WIDTH - 1),
		17987 => to_unsigned(32381, LUT_AMPL_WIDTH - 1),
		17988 => to_unsigned(32380, LUT_AMPL_WIDTH - 1),
		17989 => to_unsigned(32380, LUT_AMPL_WIDTH - 1),
		17990 => to_unsigned(32379, LUT_AMPL_WIDTH - 1),
		17991 => to_unsigned(32379, LUT_AMPL_WIDTH - 1),
		17992 => to_unsigned(32378, LUT_AMPL_WIDTH - 1),
		17993 => to_unsigned(32378, LUT_AMPL_WIDTH - 1),
		17994 => to_unsigned(32377, LUT_AMPL_WIDTH - 1),
		17995 => to_unsigned(32377, LUT_AMPL_WIDTH - 1),
		17996 => to_unsigned(32376, LUT_AMPL_WIDTH - 1),
		17997 => to_unsigned(32376, LUT_AMPL_WIDTH - 1),
		17998 => to_unsigned(32375, LUT_AMPL_WIDTH - 1),
		17999 => to_unsigned(32375, LUT_AMPL_WIDTH - 1),
		18000 => to_unsigned(32375, LUT_AMPL_WIDTH - 1),
		18001 => to_unsigned(32374, LUT_AMPL_WIDTH - 1),
		18002 => to_unsigned(32374, LUT_AMPL_WIDTH - 1),
		18003 => to_unsigned(32373, LUT_AMPL_WIDTH - 1),
		18004 => to_unsigned(32373, LUT_AMPL_WIDTH - 1),
		18005 => to_unsigned(32372, LUT_AMPL_WIDTH - 1),
		18006 => to_unsigned(32372, LUT_AMPL_WIDTH - 1),
		18007 => to_unsigned(32371, LUT_AMPL_WIDTH - 1),
		18008 => to_unsigned(32371, LUT_AMPL_WIDTH - 1),
		18009 => to_unsigned(32370, LUT_AMPL_WIDTH - 1),
		18010 => to_unsigned(32370, LUT_AMPL_WIDTH - 1),
		18011 => to_unsigned(32369, LUT_AMPL_WIDTH - 1),
		18012 => to_unsigned(32369, LUT_AMPL_WIDTH - 1),
		18013 => to_unsigned(32368, LUT_AMPL_WIDTH - 1),
		18014 => to_unsigned(32368, LUT_AMPL_WIDTH - 1),
		18015 => to_unsigned(32367, LUT_AMPL_WIDTH - 1),
		18016 => to_unsigned(32367, LUT_AMPL_WIDTH - 1),
		18017 => to_unsigned(32366, LUT_AMPL_WIDTH - 1),
		18018 => to_unsigned(32366, LUT_AMPL_WIDTH - 1),
		18019 => to_unsigned(32365, LUT_AMPL_WIDTH - 1),
		18020 => to_unsigned(32365, LUT_AMPL_WIDTH - 1),
		18021 => to_unsigned(32364, LUT_AMPL_WIDTH - 1),
		18022 => to_unsigned(32364, LUT_AMPL_WIDTH - 1),
		18023 => to_unsigned(32363, LUT_AMPL_WIDTH - 1),
		18024 => to_unsigned(32363, LUT_AMPL_WIDTH - 1),
		18025 => to_unsigned(32362, LUT_AMPL_WIDTH - 1),
		18026 => to_unsigned(32362, LUT_AMPL_WIDTH - 1),
		18027 => to_unsigned(32361, LUT_AMPL_WIDTH - 1),
		18028 => to_unsigned(32361, LUT_AMPL_WIDTH - 1),
		18029 => to_unsigned(32360, LUT_AMPL_WIDTH - 1),
		18030 => to_unsigned(32360, LUT_AMPL_WIDTH - 1),
		18031 => to_unsigned(32359, LUT_AMPL_WIDTH - 1),
		18032 => to_unsigned(32359, LUT_AMPL_WIDTH - 1),
		18033 => to_unsigned(32358, LUT_AMPL_WIDTH - 1),
		18034 => to_unsigned(32358, LUT_AMPL_WIDTH - 1),
		18035 => to_unsigned(32357, LUT_AMPL_WIDTH - 1),
		18036 => to_unsigned(32357, LUT_AMPL_WIDTH - 1),
		18037 => to_unsigned(32356, LUT_AMPL_WIDTH - 1),
		18038 => to_unsigned(32356, LUT_AMPL_WIDTH - 1),
		18039 => to_unsigned(32355, LUT_AMPL_WIDTH - 1),
		18040 => to_unsigned(32355, LUT_AMPL_WIDTH - 1),
		18041 => to_unsigned(32354, LUT_AMPL_WIDTH - 1),
		18042 => to_unsigned(32354, LUT_AMPL_WIDTH - 1),
		18043 => to_unsigned(32353, LUT_AMPL_WIDTH - 1),
		18044 => to_unsigned(32353, LUT_AMPL_WIDTH - 1),
		18045 => to_unsigned(32352, LUT_AMPL_WIDTH - 1),
		18046 => to_unsigned(32352, LUT_AMPL_WIDTH - 1),
		18047 => to_unsigned(32351, LUT_AMPL_WIDTH - 1),
		18048 => to_unsigned(32351, LUT_AMPL_WIDTH - 1),
		18049 => to_unsigned(32350, LUT_AMPL_WIDTH - 1),
		18050 => to_unsigned(32350, LUT_AMPL_WIDTH - 1),
		18051 => to_unsigned(32349, LUT_AMPL_WIDTH - 1),
		18052 => to_unsigned(32349, LUT_AMPL_WIDTH - 1),
		18053 => to_unsigned(32348, LUT_AMPL_WIDTH - 1),
		18054 => to_unsigned(32348, LUT_AMPL_WIDTH - 1),
		18055 => to_unsigned(32347, LUT_AMPL_WIDTH - 1),
		18056 => to_unsigned(32347, LUT_AMPL_WIDTH - 1),
		18057 => to_unsigned(32346, LUT_AMPL_WIDTH - 1),
		18058 => to_unsigned(32346, LUT_AMPL_WIDTH - 1),
		18059 => to_unsigned(32345, LUT_AMPL_WIDTH - 1),
		18060 => to_unsigned(32345, LUT_AMPL_WIDTH - 1),
		18061 => to_unsigned(32344, LUT_AMPL_WIDTH - 1),
		18062 => to_unsigned(32344, LUT_AMPL_WIDTH - 1),
		18063 => to_unsigned(32343, LUT_AMPL_WIDTH - 1),
		18064 => to_unsigned(32343, LUT_AMPL_WIDTH - 1),
		18065 => to_unsigned(32342, LUT_AMPL_WIDTH - 1),
		18066 => to_unsigned(32342, LUT_AMPL_WIDTH - 1),
		18067 => to_unsigned(32341, LUT_AMPL_WIDTH - 1),
		18068 => to_unsigned(32341, LUT_AMPL_WIDTH - 1),
		18069 => to_unsigned(32340, LUT_AMPL_WIDTH - 1),
		18070 => to_unsigned(32340, LUT_AMPL_WIDTH - 1),
		18071 => to_unsigned(32339, LUT_AMPL_WIDTH - 1),
		18072 => to_unsigned(32339, LUT_AMPL_WIDTH - 1),
		18073 => to_unsigned(32338, LUT_AMPL_WIDTH - 1),
		18074 => to_unsigned(32338, LUT_AMPL_WIDTH - 1),
		18075 => to_unsigned(32337, LUT_AMPL_WIDTH - 1),
		18076 => to_unsigned(32337, LUT_AMPL_WIDTH - 1),
		18077 => to_unsigned(32336, LUT_AMPL_WIDTH - 1),
		18078 => to_unsigned(32336, LUT_AMPL_WIDTH - 1),
		18079 => to_unsigned(32335, LUT_AMPL_WIDTH - 1),
		18080 => to_unsigned(32335, LUT_AMPL_WIDTH - 1),
		18081 => to_unsigned(32334, LUT_AMPL_WIDTH - 1),
		18082 => to_unsigned(32334, LUT_AMPL_WIDTH - 1),
		18083 => to_unsigned(32333, LUT_AMPL_WIDTH - 1),
		18084 => to_unsigned(32333, LUT_AMPL_WIDTH - 1),
		18085 => to_unsigned(32332, LUT_AMPL_WIDTH - 1),
		18086 => to_unsigned(32332, LUT_AMPL_WIDTH - 1),
		18087 => to_unsigned(32331, LUT_AMPL_WIDTH - 1),
		18088 => to_unsigned(32331, LUT_AMPL_WIDTH - 1),
		18089 => to_unsigned(32330, LUT_AMPL_WIDTH - 1),
		18090 => to_unsigned(32330, LUT_AMPL_WIDTH - 1),
		18091 => to_unsigned(32329, LUT_AMPL_WIDTH - 1),
		18092 => to_unsigned(32329, LUT_AMPL_WIDTH - 1),
		18093 => to_unsigned(32328, LUT_AMPL_WIDTH - 1),
		18094 => to_unsigned(32328, LUT_AMPL_WIDTH - 1),
		18095 => to_unsigned(32327, LUT_AMPL_WIDTH - 1),
		18096 => to_unsigned(32327, LUT_AMPL_WIDTH - 1),
		18097 => to_unsigned(32326, LUT_AMPL_WIDTH - 1),
		18098 => to_unsigned(32326, LUT_AMPL_WIDTH - 1),
		18099 => to_unsigned(32325, LUT_AMPL_WIDTH - 1),
		18100 => to_unsigned(32325, LUT_AMPL_WIDTH - 1),
		18101 => to_unsigned(32324, LUT_AMPL_WIDTH - 1),
		18102 => to_unsigned(32324, LUT_AMPL_WIDTH - 1),
		18103 => to_unsigned(32323, LUT_AMPL_WIDTH - 1),
		18104 => to_unsigned(32322, LUT_AMPL_WIDTH - 1),
		18105 => to_unsigned(32322, LUT_AMPL_WIDTH - 1),
		18106 => to_unsigned(32321, LUT_AMPL_WIDTH - 1),
		18107 => to_unsigned(32321, LUT_AMPL_WIDTH - 1),
		18108 => to_unsigned(32320, LUT_AMPL_WIDTH - 1),
		18109 => to_unsigned(32320, LUT_AMPL_WIDTH - 1),
		18110 => to_unsigned(32319, LUT_AMPL_WIDTH - 1),
		18111 => to_unsigned(32319, LUT_AMPL_WIDTH - 1),
		18112 => to_unsigned(32318, LUT_AMPL_WIDTH - 1),
		18113 => to_unsigned(32318, LUT_AMPL_WIDTH - 1),
		18114 => to_unsigned(32317, LUT_AMPL_WIDTH - 1),
		18115 => to_unsigned(32317, LUT_AMPL_WIDTH - 1),
		18116 => to_unsigned(32316, LUT_AMPL_WIDTH - 1),
		18117 => to_unsigned(32316, LUT_AMPL_WIDTH - 1),
		18118 => to_unsigned(32315, LUT_AMPL_WIDTH - 1),
		18119 => to_unsigned(32315, LUT_AMPL_WIDTH - 1),
		18120 => to_unsigned(32314, LUT_AMPL_WIDTH - 1),
		18121 => to_unsigned(32314, LUT_AMPL_WIDTH - 1),
		18122 => to_unsigned(32313, LUT_AMPL_WIDTH - 1),
		18123 => to_unsigned(32313, LUT_AMPL_WIDTH - 1),
		18124 => to_unsigned(32312, LUT_AMPL_WIDTH - 1),
		18125 => to_unsigned(32312, LUT_AMPL_WIDTH - 1),
		18126 => to_unsigned(32311, LUT_AMPL_WIDTH - 1),
		18127 => to_unsigned(32311, LUT_AMPL_WIDTH - 1),
		18128 => to_unsigned(32310, LUT_AMPL_WIDTH - 1),
		18129 => to_unsigned(32310, LUT_AMPL_WIDTH - 1),
		18130 => to_unsigned(32309, LUT_AMPL_WIDTH - 1),
		18131 => to_unsigned(32308, LUT_AMPL_WIDTH - 1),
		18132 => to_unsigned(32308, LUT_AMPL_WIDTH - 1),
		18133 => to_unsigned(32307, LUT_AMPL_WIDTH - 1),
		18134 => to_unsigned(32307, LUT_AMPL_WIDTH - 1),
		18135 => to_unsigned(32306, LUT_AMPL_WIDTH - 1),
		18136 => to_unsigned(32306, LUT_AMPL_WIDTH - 1),
		18137 => to_unsigned(32305, LUT_AMPL_WIDTH - 1),
		18138 => to_unsigned(32305, LUT_AMPL_WIDTH - 1),
		18139 => to_unsigned(32304, LUT_AMPL_WIDTH - 1),
		18140 => to_unsigned(32304, LUT_AMPL_WIDTH - 1),
		18141 => to_unsigned(32303, LUT_AMPL_WIDTH - 1),
		18142 => to_unsigned(32303, LUT_AMPL_WIDTH - 1),
		18143 => to_unsigned(32302, LUT_AMPL_WIDTH - 1),
		18144 => to_unsigned(32302, LUT_AMPL_WIDTH - 1),
		18145 => to_unsigned(32301, LUT_AMPL_WIDTH - 1),
		18146 => to_unsigned(32301, LUT_AMPL_WIDTH - 1),
		18147 => to_unsigned(32300, LUT_AMPL_WIDTH - 1),
		18148 => to_unsigned(32300, LUT_AMPL_WIDTH - 1),
		18149 => to_unsigned(32299, LUT_AMPL_WIDTH - 1),
		18150 => to_unsigned(32298, LUT_AMPL_WIDTH - 1),
		18151 => to_unsigned(32298, LUT_AMPL_WIDTH - 1),
		18152 => to_unsigned(32297, LUT_AMPL_WIDTH - 1),
		18153 => to_unsigned(32297, LUT_AMPL_WIDTH - 1),
		18154 => to_unsigned(32296, LUT_AMPL_WIDTH - 1),
		18155 => to_unsigned(32296, LUT_AMPL_WIDTH - 1),
		18156 => to_unsigned(32295, LUT_AMPL_WIDTH - 1),
		18157 => to_unsigned(32295, LUT_AMPL_WIDTH - 1),
		18158 => to_unsigned(32294, LUT_AMPL_WIDTH - 1),
		18159 => to_unsigned(32294, LUT_AMPL_WIDTH - 1),
		18160 => to_unsigned(32293, LUT_AMPL_WIDTH - 1),
		18161 => to_unsigned(32293, LUT_AMPL_WIDTH - 1),
		18162 => to_unsigned(32292, LUT_AMPL_WIDTH - 1),
		18163 => to_unsigned(32292, LUT_AMPL_WIDTH - 1),
		18164 => to_unsigned(32291, LUT_AMPL_WIDTH - 1),
		18165 => to_unsigned(32290, LUT_AMPL_WIDTH - 1),
		18166 => to_unsigned(32290, LUT_AMPL_WIDTH - 1),
		18167 => to_unsigned(32289, LUT_AMPL_WIDTH - 1),
		18168 => to_unsigned(32289, LUT_AMPL_WIDTH - 1),
		18169 => to_unsigned(32288, LUT_AMPL_WIDTH - 1),
		18170 => to_unsigned(32288, LUT_AMPL_WIDTH - 1),
		18171 => to_unsigned(32287, LUT_AMPL_WIDTH - 1),
		18172 => to_unsigned(32287, LUT_AMPL_WIDTH - 1),
		18173 => to_unsigned(32286, LUT_AMPL_WIDTH - 1),
		18174 => to_unsigned(32286, LUT_AMPL_WIDTH - 1),
		18175 => to_unsigned(32285, LUT_AMPL_WIDTH - 1),
		18176 => to_unsigned(32285, LUT_AMPL_WIDTH - 1),
		18177 => to_unsigned(32284, LUT_AMPL_WIDTH - 1),
		18178 => to_unsigned(32284, LUT_AMPL_WIDTH - 1),
		18179 => to_unsigned(32283, LUT_AMPL_WIDTH - 1),
		18180 => to_unsigned(32282, LUT_AMPL_WIDTH - 1),
		18181 => to_unsigned(32282, LUT_AMPL_WIDTH - 1),
		18182 => to_unsigned(32281, LUT_AMPL_WIDTH - 1),
		18183 => to_unsigned(32281, LUT_AMPL_WIDTH - 1),
		18184 => to_unsigned(32280, LUT_AMPL_WIDTH - 1),
		18185 => to_unsigned(32280, LUT_AMPL_WIDTH - 1),
		18186 => to_unsigned(32279, LUT_AMPL_WIDTH - 1),
		18187 => to_unsigned(32279, LUT_AMPL_WIDTH - 1),
		18188 => to_unsigned(32278, LUT_AMPL_WIDTH - 1),
		18189 => to_unsigned(32278, LUT_AMPL_WIDTH - 1),
		18190 => to_unsigned(32277, LUT_AMPL_WIDTH - 1),
		18191 => to_unsigned(32277, LUT_AMPL_WIDTH - 1),
		18192 => to_unsigned(32276, LUT_AMPL_WIDTH - 1),
		18193 => to_unsigned(32275, LUT_AMPL_WIDTH - 1),
		18194 => to_unsigned(32275, LUT_AMPL_WIDTH - 1),
		18195 => to_unsigned(32274, LUT_AMPL_WIDTH - 1),
		18196 => to_unsigned(32274, LUT_AMPL_WIDTH - 1),
		18197 => to_unsigned(32273, LUT_AMPL_WIDTH - 1),
		18198 => to_unsigned(32273, LUT_AMPL_WIDTH - 1),
		18199 => to_unsigned(32272, LUT_AMPL_WIDTH - 1),
		18200 => to_unsigned(32272, LUT_AMPL_WIDTH - 1),
		18201 => to_unsigned(32271, LUT_AMPL_WIDTH - 1),
		18202 => to_unsigned(32271, LUT_AMPL_WIDTH - 1),
		18203 => to_unsigned(32270, LUT_AMPL_WIDTH - 1),
		18204 => to_unsigned(32269, LUT_AMPL_WIDTH - 1),
		18205 => to_unsigned(32269, LUT_AMPL_WIDTH - 1),
		18206 => to_unsigned(32268, LUT_AMPL_WIDTH - 1),
		18207 => to_unsigned(32268, LUT_AMPL_WIDTH - 1),
		18208 => to_unsigned(32267, LUT_AMPL_WIDTH - 1),
		18209 => to_unsigned(32267, LUT_AMPL_WIDTH - 1),
		18210 => to_unsigned(32266, LUT_AMPL_WIDTH - 1),
		18211 => to_unsigned(32266, LUT_AMPL_WIDTH - 1),
		18212 => to_unsigned(32265, LUT_AMPL_WIDTH - 1),
		18213 => to_unsigned(32265, LUT_AMPL_WIDTH - 1),
		18214 => to_unsigned(32264, LUT_AMPL_WIDTH - 1),
		18215 => to_unsigned(32263, LUT_AMPL_WIDTH - 1),
		18216 => to_unsigned(32263, LUT_AMPL_WIDTH - 1),
		18217 => to_unsigned(32262, LUT_AMPL_WIDTH - 1),
		18218 => to_unsigned(32262, LUT_AMPL_WIDTH - 1),
		18219 => to_unsigned(32261, LUT_AMPL_WIDTH - 1),
		18220 => to_unsigned(32261, LUT_AMPL_WIDTH - 1),
		18221 => to_unsigned(32260, LUT_AMPL_WIDTH - 1),
		18222 => to_unsigned(32260, LUT_AMPL_WIDTH - 1),
		18223 => to_unsigned(32259, LUT_AMPL_WIDTH - 1),
		18224 => to_unsigned(32258, LUT_AMPL_WIDTH - 1),
		18225 => to_unsigned(32258, LUT_AMPL_WIDTH - 1),
		18226 => to_unsigned(32257, LUT_AMPL_WIDTH - 1),
		18227 => to_unsigned(32257, LUT_AMPL_WIDTH - 1),
		18228 => to_unsigned(32256, LUT_AMPL_WIDTH - 1),
		18229 => to_unsigned(32256, LUT_AMPL_WIDTH - 1),
		18230 => to_unsigned(32255, LUT_AMPL_WIDTH - 1),
		18231 => to_unsigned(32255, LUT_AMPL_WIDTH - 1),
		18232 => to_unsigned(32254, LUT_AMPL_WIDTH - 1),
		18233 => to_unsigned(32253, LUT_AMPL_WIDTH - 1),
		18234 => to_unsigned(32253, LUT_AMPL_WIDTH - 1),
		18235 => to_unsigned(32252, LUT_AMPL_WIDTH - 1),
		18236 => to_unsigned(32252, LUT_AMPL_WIDTH - 1),
		18237 => to_unsigned(32251, LUT_AMPL_WIDTH - 1),
		18238 => to_unsigned(32251, LUT_AMPL_WIDTH - 1),
		18239 => to_unsigned(32250, LUT_AMPL_WIDTH - 1),
		18240 => to_unsigned(32250, LUT_AMPL_WIDTH - 1),
		18241 => to_unsigned(32249, LUT_AMPL_WIDTH - 1),
		18242 => to_unsigned(32248, LUT_AMPL_WIDTH - 1),
		18243 => to_unsigned(32248, LUT_AMPL_WIDTH - 1),
		18244 => to_unsigned(32247, LUT_AMPL_WIDTH - 1),
		18245 => to_unsigned(32247, LUT_AMPL_WIDTH - 1),
		18246 => to_unsigned(32246, LUT_AMPL_WIDTH - 1),
		18247 => to_unsigned(32246, LUT_AMPL_WIDTH - 1),
		18248 => to_unsigned(32245, LUT_AMPL_WIDTH - 1),
		18249 => to_unsigned(32245, LUT_AMPL_WIDTH - 1),
		18250 => to_unsigned(32244, LUT_AMPL_WIDTH - 1),
		18251 => to_unsigned(32243, LUT_AMPL_WIDTH - 1),
		18252 => to_unsigned(32243, LUT_AMPL_WIDTH - 1),
		18253 => to_unsigned(32242, LUT_AMPL_WIDTH - 1),
		18254 => to_unsigned(32242, LUT_AMPL_WIDTH - 1),
		18255 => to_unsigned(32241, LUT_AMPL_WIDTH - 1),
		18256 => to_unsigned(32241, LUT_AMPL_WIDTH - 1),
		18257 => to_unsigned(32240, LUT_AMPL_WIDTH - 1),
		18258 => to_unsigned(32240, LUT_AMPL_WIDTH - 1),
		18259 => to_unsigned(32239, LUT_AMPL_WIDTH - 1),
		18260 => to_unsigned(32238, LUT_AMPL_WIDTH - 1),
		18261 => to_unsigned(32238, LUT_AMPL_WIDTH - 1),
		18262 => to_unsigned(32237, LUT_AMPL_WIDTH - 1),
		18263 => to_unsigned(32237, LUT_AMPL_WIDTH - 1),
		18264 => to_unsigned(32236, LUT_AMPL_WIDTH - 1),
		18265 => to_unsigned(32236, LUT_AMPL_WIDTH - 1),
		18266 => to_unsigned(32235, LUT_AMPL_WIDTH - 1),
		18267 => to_unsigned(32234, LUT_AMPL_WIDTH - 1),
		18268 => to_unsigned(32234, LUT_AMPL_WIDTH - 1),
		18269 => to_unsigned(32233, LUT_AMPL_WIDTH - 1),
		18270 => to_unsigned(32233, LUT_AMPL_WIDTH - 1),
		18271 => to_unsigned(32232, LUT_AMPL_WIDTH - 1),
		18272 => to_unsigned(32232, LUT_AMPL_WIDTH - 1),
		18273 => to_unsigned(32231, LUT_AMPL_WIDTH - 1),
		18274 => to_unsigned(32231, LUT_AMPL_WIDTH - 1),
		18275 => to_unsigned(32230, LUT_AMPL_WIDTH - 1),
		18276 => to_unsigned(32229, LUT_AMPL_WIDTH - 1),
		18277 => to_unsigned(32229, LUT_AMPL_WIDTH - 1),
		18278 => to_unsigned(32228, LUT_AMPL_WIDTH - 1),
		18279 => to_unsigned(32228, LUT_AMPL_WIDTH - 1),
		18280 => to_unsigned(32227, LUT_AMPL_WIDTH - 1),
		18281 => to_unsigned(32227, LUT_AMPL_WIDTH - 1),
		18282 => to_unsigned(32226, LUT_AMPL_WIDTH - 1),
		18283 => to_unsigned(32225, LUT_AMPL_WIDTH - 1),
		18284 => to_unsigned(32225, LUT_AMPL_WIDTH - 1),
		18285 => to_unsigned(32224, LUT_AMPL_WIDTH - 1),
		18286 => to_unsigned(32224, LUT_AMPL_WIDTH - 1),
		18287 => to_unsigned(32223, LUT_AMPL_WIDTH - 1),
		18288 => to_unsigned(32223, LUT_AMPL_WIDTH - 1),
		18289 => to_unsigned(32222, LUT_AMPL_WIDTH - 1),
		18290 => to_unsigned(32221, LUT_AMPL_WIDTH - 1),
		18291 => to_unsigned(32221, LUT_AMPL_WIDTH - 1),
		18292 => to_unsigned(32220, LUT_AMPL_WIDTH - 1),
		18293 => to_unsigned(32220, LUT_AMPL_WIDTH - 1),
		18294 => to_unsigned(32219, LUT_AMPL_WIDTH - 1),
		18295 => to_unsigned(32219, LUT_AMPL_WIDTH - 1),
		18296 => to_unsigned(32218, LUT_AMPL_WIDTH - 1),
		18297 => to_unsigned(32217, LUT_AMPL_WIDTH - 1),
		18298 => to_unsigned(32217, LUT_AMPL_WIDTH - 1),
		18299 => to_unsigned(32216, LUT_AMPL_WIDTH - 1),
		18300 => to_unsigned(32216, LUT_AMPL_WIDTH - 1),
		18301 => to_unsigned(32215, LUT_AMPL_WIDTH - 1),
		18302 => to_unsigned(32215, LUT_AMPL_WIDTH - 1),
		18303 => to_unsigned(32214, LUT_AMPL_WIDTH - 1),
		18304 => to_unsigned(32213, LUT_AMPL_WIDTH - 1),
		18305 => to_unsigned(32213, LUT_AMPL_WIDTH - 1),
		18306 => to_unsigned(32212, LUT_AMPL_WIDTH - 1),
		18307 => to_unsigned(32212, LUT_AMPL_WIDTH - 1),
		18308 => to_unsigned(32211, LUT_AMPL_WIDTH - 1),
		18309 => to_unsigned(32211, LUT_AMPL_WIDTH - 1),
		18310 => to_unsigned(32210, LUT_AMPL_WIDTH - 1),
		18311 => to_unsigned(32209, LUT_AMPL_WIDTH - 1),
		18312 => to_unsigned(32209, LUT_AMPL_WIDTH - 1),
		18313 => to_unsigned(32208, LUT_AMPL_WIDTH - 1),
		18314 => to_unsigned(32208, LUT_AMPL_WIDTH - 1),
		18315 => to_unsigned(32207, LUT_AMPL_WIDTH - 1),
		18316 => to_unsigned(32206, LUT_AMPL_WIDTH - 1),
		18317 => to_unsigned(32206, LUT_AMPL_WIDTH - 1),
		18318 => to_unsigned(32205, LUT_AMPL_WIDTH - 1),
		18319 => to_unsigned(32205, LUT_AMPL_WIDTH - 1),
		18320 => to_unsigned(32204, LUT_AMPL_WIDTH - 1),
		18321 => to_unsigned(32204, LUT_AMPL_WIDTH - 1),
		18322 => to_unsigned(32203, LUT_AMPL_WIDTH - 1),
		18323 => to_unsigned(32202, LUT_AMPL_WIDTH - 1),
		18324 => to_unsigned(32202, LUT_AMPL_WIDTH - 1),
		18325 => to_unsigned(32201, LUT_AMPL_WIDTH - 1),
		18326 => to_unsigned(32201, LUT_AMPL_WIDTH - 1),
		18327 => to_unsigned(32200, LUT_AMPL_WIDTH - 1),
		18328 => to_unsigned(32200, LUT_AMPL_WIDTH - 1),
		18329 => to_unsigned(32199, LUT_AMPL_WIDTH - 1),
		18330 => to_unsigned(32198, LUT_AMPL_WIDTH - 1),
		18331 => to_unsigned(32198, LUT_AMPL_WIDTH - 1),
		18332 => to_unsigned(32197, LUT_AMPL_WIDTH - 1),
		18333 => to_unsigned(32197, LUT_AMPL_WIDTH - 1),
		18334 => to_unsigned(32196, LUT_AMPL_WIDTH - 1),
		18335 => to_unsigned(32195, LUT_AMPL_WIDTH - 1),
		18336 => to_unsigned(32195, LUT_AMPL_WIDTH - 1),
		18337 => to_unsigned(32194, LUT_AMPL_WIDTH - 1),
		18338 => to_unsigned(32194, LUT_AMPL_WIDTH - 1),
		18339 => to_unsigned(32193, LUT_AMPL_WIDTH - 1),
		18340 => to_unsigned(32193, LUT_AMPL_WIDTH - 1),
		18341 => to_unsigned(32192, LUT_AMPL_WIDTH - 1),
		18342 => to_unsigned(32191, LUT_AMPL_WIDTH - 1),
		18343 => to_unsigned(32191, LUT_AMPL_WIDTH - 1),
		18344 => to_unsigned(32190, LUT_AMPL_WIDTH - 1),
		18345 => to_unsigned(32190, LUT_AMPL_WIDTH - 1),
		18346 => to_unsigned(32189, LUT_AMPL_WIDTH - 1),
		18347 => to_unsigned(32188, LUT_AMPL_WIDTH - 1),
		18348 => to_unsigned(32188, LUT_AMPL_WIDTH - 1),
		18349 => to_unsigned(32187, LUT_AMPL_WIDTH - 1),
		18350 => to_unsigned(32187, LUT_AMPL_WIDTH - 1),
		18351 => to_unsigned(32186, LUT_AMPL_WIDTH - 1),
		18352 => to_unsigned(32185, LUT_AMPL_WIDTH - 1),
		18353 => to_unsigned(32185, LUT_AMPL_WIDTH - 1),
		18354 => to_unsigned(32184, LUT_AMPL_WIDTH - 1),
		18355 => to_unsigned(32184, LUT_AMPL_WIDTH - 1),
		18356 => to_unsigned(32183, LUT_AMPL_WIDTH - 1),
		18357 => to_unsigned(32183, LUT_AMPL_WIDTH - 1),
		18358 => to_unsigned(32182, LUT_AMPL_WIDTH - 1),
		18359 => to_unsigned(32181, LUT_AMPL_WIDTH - 1),
		18360 => to_unsigned(32181, LUT_AMPL_WIDTH - 1),
		18361 => to_unsigned(32180, LUT_AMPL_WIDTH - 1),
		18362 => to_unsigned(32180, LUT_AMPL_WIDTH - 1),
		18363 => to_unsigned(32179, LUT_AMPL_WIDTH - 1),
		18364 => to_unsigned(32178, LUT_AMPL_WIDTH - 1),
		18365 => to_unsigned(32178, LUT_AMPL_WIDTH - 1),
		18366 => to_unsigned(32177, LUT_AMPL_WIDTH - 1),
		18367 => to_unsigned(32177, LUT_AMPL_WIDTH - 1),
		18368 => to_unsigned(32176, LUT_AMPL_WIDTH - 1),
		18369 => to_unsigned(32175, LUT_AMPL_WIDTH - 1),
		18370 => to_unsigned(32175, LUT_AMPL_WIDTH - 1),
		18371 => to_unsigned(32174, LUT_AMPL_WIDTH - 1),
		18372 => to_unsigned(32174, LUT_AMPL_WIDTH - 1),
		18373 => to_unsigned(32173, LUT_AMPL_WIDTH - 1),
		18374 => to_unsigned(32172, LUT_AMPL_WIDTH - 1),
		18375 => to_unsigned(32172, LUT_AMPL_WIDTH - 1),
		18376 => to_unsigned(32171, LUT_AMPL_WIDTH - 1),
		18377 => to_unsigned(32171, LUT_AMPL_WIDTH - 1),
		18378 => to_unsigned(32170, LUT_AMPL_WIDTH - 1),
		18379 => to_unsigned(32169, LUT_AMPL_WIDTH - 1),
		18380 => to_unsigned(32169, LUT_AMPL_WIDTH - 1),
		18381 => to_unsigned(32168, LUT_AMPL_WIDTH - 1),
		18382 => to_unsigned(32168, LUT_AMPL_WIDTH - 1),
		18383 => to_unsigned(32167, LUT_AMPL_WIDTH - 1),
		18384 => to_unsigned(32166, LUT_AMPL_WIDTH - 1),
		18385 => to_unsigned(32166, LUT_AMPL_WIDTH - 1),
		18386 => to_unsigned(32165, LUT_AMPL_WIDTH - 1),
		18387 => to_unsigned(32165, LUT_AMPL_WIDTH - 1),
		18388 => to_unsigned(32164, LUT_AMPL_WIDTH - 1),
		18389 => to_unsigned(32163, LUT_AMPL_WIDTH - 1),
		18390 => to_unsigned(32163, LUT_AMPL_WIDTH - 1),
		18391 => to_unsigned(32162, LUT_AMPL_WIDTH - 1),
		18392 => to_unsigned(32162, LUT_AMPL_WIDTH - 1),
		18393 => to_unsigned(32161, LUT_AMPL_WIDTH - 1),
		18394 => to_unsigned(32160, LUT_AMPL_WIDTH - 1),
		18395 => to_unsigned(32160, LUT_AMPL_WIDTH - 1),
		18396 => to_unsigned(32159, LUT_AMPL_WIDTH - 1),
		18397 => to_unsigned(32159, LUT_AMPL_WIDTH - 1),
		18398 => to_unsigned(32158, LUT_AMPL_WIDTH - 1),
		18399 => to_unsigned(32157, LUT_AMPL_WIDTH - 1),
		18400 => to_unsigned(32157, LUT_AMPL_WIDTH - 1),
		18401 => to_unsigned(32156, LUT_AMPL_WIDTH - 1),
		18402 => to_unsigned(32156, LUT_AMPL_WIDTH - 1),
		18403 => to_unsigned(32155, LUT_AMPL_WIDTH - 1),
		18404 => to_unsigned(32154, LUT_AMPL_WIDTH - 1),
		18405 => to_unsigned(32154, LUT_AMPL_WIDTH - 1),
		18406 => to_unsigned(32153, LUT_AMPL_WIDTH - 1),
		18407 => to_unsigned(32153, LUT_AMPL_WIDTH - 1),
		18408 => to_unsigned(32152, LUT_AMPL_WIDTH - 1),
		18409 => to_unsigned(32151, LUT_AMPL_WIDTH - 1),
		18410 => to_unsigned(32151, LUT_AMPL_WIDTH - 1),
		18411 => to_unsigned(32150, LUT_AMPL_WIDTH - 1),
		18412 => to_unsigned(32150, LUT_AMPL_WIDTH - 1),
		18413 => to_unsigned(32149, LUT_AMPL_WIDTH - 1),
		18414 => to_unsigned(32148, LUT_AMPL_WIDTH - 1),
		18415 => to_unsigned(32148, LUT_AMPL_WIDTH - 1),
		18416 => to_unsigned(32147, LUT_AMPL_WIDTH - 1),
		18417 => to_unsigned(32147, LUT_AMPL_WIDTH - 1),
		18418 => to_unsigned(32146, LUT_AMPL_WIDTH - 1),
		18419 => to_unsigned(32145, LUT_AMPL_WIDTH - 1),
		18420 => to_unsigned(32145, LUT_AMPL_WIDTH - 1),
		18421 => to_unsigned(32144, LUT_AMPL_WIDTH - 1),
		18422 => to_unsigned(32144, LUT_AMPL_WIDTH - 1),
		18423 => to_unsigned(32143, LUT_AMPL_WIDTH - 1),
		18424 => to_unsigned(32142, LUT_AMPL_WIDTH - 1),
		18425 => to_unsigned(32142, LUT_AMPL_WIDTH - 1),
		18426 => to_unsigned(32141, LUT_AMPL_WIDTH - 1),
		18427 => to_unsigned(32140, LUT_AMPL_WIDTH - 1),
		18428 => to_unsigned(32140, LUT_AMPL_WIDTH - 1),
		18429 => to_unsigned(32139, LUT_AMPL_WIDTH - 1),
		18430 => to_unsigned(32139, LUT_AMPL_WIDTH - 1),
		18431 => to_unsigned(32138, LUT_AMPL_WIDTH - 1),
		18432 => to_unsigned(32137, LUT_AMPL_WIDTH - 1),
		18433 => to_unsigned(32137, LUT_AMPL_WIDTH - 1),
		18434 => to_unsigned(32136, LUT_AMPL_WIDTH - 1),
		18435 => to_unsigned(32136, LUT_AMPL_WIDTH - 1),
		18436 => to_unsigned(32135, LUT_AMPL_WIDTH - 1),
		18437 => to_unsigned(32134, LUT_AMPL_WIDTH - 1),
		18438 => to_unsigned(32134, LUT_AMPL_WIDTH - 1),
		18439 => to_unsigned(32133, LUT_AMPL_WIDTH - 1),
		18440 => to_unsigned(32132, LUT_AMPL_WIDTH - 1),
		18441 => to_unsigned(32132, LUT_AMPL_WIDTH - 1),
		18442 => to_unsigned(32131, LUT_AMPL_WIDTH - 1),
		18443 => to_unsigned(32131, LUT_AMPL_WIDTH - 1),
		18444 => to_unsigned(32130, LUT_AMPL_WIDTH - 1),
		18445 => to_unsigned(32129, LUT_AMPL_WIDTH - 1),
		18446 => to_unsigned(32129, LUT_AMPL_WIDTH - 1),
		18447 => to_unsigned(32128, LUT_AMPL_WIDTH - 1),
		18448 => to_unsigned(32128, LUT_AMPL_WIDTH - 1),
		18449 => to_unsigned(32127, LUT_AMPL_WIDTH - 1),
		18450 => to_unsigned(32126, LUT_AMPL_WIDTH - 1),
		18451 => to_unsigned(32126, LUT_AMPL_WIDTH - 1),
		18452 => to_unsigned(32125, LUT_AMPL_WIDTH - 1),
		18453 => to_unsigned(32124, LUT_AMPL_WIDTH - 1),
		18454 => to_unsigned(32124, LUT_AMPL_WIDTH - 1),
		18455 => to_unsigned(32123, LUT_AMPL_WIDTH - 1),
		18456 => to_unsigned(32123, LUT_AMPL_WIDTH - 1),
		18457 => to_unsigned(32122, LUT_AMPL_WIDTH - 1),
		18458 => to_unsigned(32121, LUT_AMPL_WIDTH - 1),
		18459 => to_unsigned(32121, LUT_AMPL_WIDTH - 1),
		18460 => to_unsigned(32120, LUT_AMPL_WIDTH - 1),
		18461 => to_unsigned(32119, LUT_AMPL_WIDTH - 1),
		18462 => to_unsigned(32119, LUT_AMPL_WIDTH - 1),
		18463 => to_unsigned(32118, LUT_AMPL_WIDTH - 1),
		18464 => to_unsigned(32118, LUT_AMPL_WIDTH - 1),
		18465 => to_unsigned(32117, LUT_AMPL_WIDTH - 1),
		18466 => to_unsigned(32116, LUT_AMPL_WIDTH - 1),
		18467 => to_unsigned(32116, LUT_AMPL_WIDTH - 1),
		18468 => to_unsigned(32115, LUT_AMPL_WIDTH - 1),
		18469 => to_unsigned(32115, LUT_AMPL_WIDTH - 1),
		18470 => to_unsigned(32114, LUT_AMPL_WIDTH - 1),
		18471 => to_unsigned(32113, LUT_AMPL_WIDTH - 1),
		18472 => to_unsigned(32113, LUT_AMPL_WIDTH - 1),
		18473 => to_unsigned(32112, LUT_AMPL_WIDTH - 1),
		18474 => to_unsigned(32111, LUT_AMPL_WIDTH - 1),
		18475 => to_unsigned(32111, LUT_AMPL_WIDTH - 1),
		18476 => to_unsigned(32110, LUT_AMPL_WIDTH - 1),
		18477 => to_unsigned(32110, LUT_AMPL_WIDTH - 1),
		18478 => to_unsigned(32109, LUT_AMPL_WIDTH - 1),
		18479 => to_unsigned(32108, LUT_AMPL_WIDTH - 1),
		18480 => to_unsigned(32108, LUT_AMPL_WIDTH - 1),
		18481 => to_unsigned(32107, LUT_AMPL_WIDTH - 1),
		18482 => to_unsigned(32106, LUT_AMPL_WIDTH - 1),
		18483 => to_unsigned(32106, LUT_AMPL_WIDTH - 1),
		18484 => to_unsigned(32105, LUT_AMPL_WIDTH - 1),
		18485 => to_unsigned(32104, LUT_AMPL_WIDTH - 1),
		18486 => to_unsigned(32104, LUT_AMPL_WIDTH - 1),
		18487 => to_unsigned(32103, LUT_AMPL_WIDTH - 1),
		18488 => to_unsigned(32103, LUT_AMPL_WIDTH - 1),
		18489 => to_unsigned(32102, LUT_AMPL_WIDTH - 1),
		18490 => to_unsigned(32101, LUT_AMPL_WIDTH - 1),
		18491 => to_unsigned(32101, LUT_AMPL_WIDTH - 1),
		18492 => to_unsigned(32100, LUT_AMPL_WIDTH - 1),
		18493 => to_unsigned(32099, LUT_AMPL_WIDTH - 1),
		18494 => to_unsigned(32099, LUT_AMPL_WIDTH - 1),
		18495 => to_unsigned(32098, LUT_AMPL_WIDTH - 1),
		18496 => to_unsigned(32098, LUT_AMPL_WIDTH - 1),
		18497 => to_unsigned(32097, LUT_AMPL_WIDTH - 1),
		18498 => to_unsigned(32096, LUT_AMPL_WIDTH - 1),
		18499 => to_unsigned(32096, LUT_AMPL_WIDTH - 1),
		18500 => to_unsigned(32095, LUT_AMPL_WIDTH - 1),
		18501 => to_unsigned(32094, LUT_AMPL_WIDTH - 1),
		18502 => to_unsigned(32094, LUT_AMPL_WIDTH - 1),
		18503 => to_unsigned(32093, LUT_AMPL_WIDTH - 1),
		18504 => to_unsigned(32092, LUT_AMPL_WIDTH - 1),
		18505 => to_unsigned(32092, LUT_AMPL_WIDTH - 1),
		18506 => to_unsigned(32091, LUT_AMPL_WIDTH - 1),
		18507 => to_unsigned(32091, LUT_AMPL_WIDTH - 1),
		18508 => to_unsigned(32090, LUT_AMPL_WIDTH - 1),
		18509 => to_unsigned(32089, LUT_AMPL_WIDTH - 1),
		18510 => to_unsigned(32089, LUT_AMPL_WIDTH - 1),
		18511 => to_unsigned(32088, LUT_AMPL_WIDTH - 1),
		18512 => to_unsigned(32087, LUT_AMPL_WIDTH - 1),
		18513 => to_unsigned(32087, LUT_AMPL_WIDTH - 1),
		18514 => to_unsigned(32086, LUT_AMPL_WIDTH - 1),
		18515 => to_unsigned(32086, LUT_AMPL_WIDTH - 1),
		18516 => to_unsigned(32085, LUT_AMPL_WIDTH - 1),
		18517 => to_unsigned(32084, LUT_AMPL_WIDTH - 1),
		18518 => to_unsigned(32084, LUT_AMPL_WIDTH - 1),
		18519 => to_unsigned(32083, LUT_AMPL_WIDTH - 1),
		18520 => to_unsigned(32082, LUT_AMPL_WIDTH - 1),
		18521 => to_unsigned(32082, LUT_AMPL_WIDTH - 1),
		18522 => to_unsigned(32081, LUT_AMPL_WIDTH - 1),
		18523 => to_unsigned(32080, LUT_AMPL_WIDTH - 1),
		18524 => to_unsigned(32080, LUT_AMPL_WIDTH - 1),
		18525 => to_unsigned(32079, LUT_AMPL_WIDTH - 1),
		18526 => to_unsigned(32078, LUT_AMPL_WIDTH - 1),
		18527 => to_unsigned(32078, LUT_AMPL_WIDTH - 1),
		18528 => to_unsigned(32077, LUT_AMPL_WIDTH - 1),
		18529 => to_unsigned(32077, LUT_AMPL_WIDTH - 1),
		18530 => to_unsigned(32076, LUT_AMPL_WIDTH - 1),
		18531 => to_unsigned(32075, LUT_AMPL_WIDTH - 1),
		18532 => to_unsigned(32075, LUT_AMPL_WIDTH - 1),
		18533 => to_unsigned(32074, LUT_AMPL_WIDTH - 1),
		18534 => to_unsigned(32073, LUT_AMPL_WIDTH - 1),
		18535 => to_unsigned(32073, LUT_AMPL_WIDTH - 1),
		18536 => to_unsigned(32072, LUT_AMPL_WIDTH - 1),
		18537 => to_unsigned(32071, LUT_AMPL_WIDTH - 1),
		18538 => to_unsigned(32071, LUT_AMPL_WIDTH - 1),
		18539 => to_unsigned(32070, LUT_AMPL_WIDTH - 1),
		18540 => to_unsigned(32069, LUT_AMPL_WIDTH - 1),
		18541 => to_unsigned(32069, LUT_AMPL_WIDTH - 1),
		18542 => to_unsigned(32068, LUT_AMPL_WIDTH - 1),
		18543 => to_unsigned(32068, LUT_AMPL_WIDTH - 1),
		18544 => to_unsigned(32067, LUT_AMPL_WIDTH - 1),
		18545 => to_unsigned(32066, LUT_AMPL_WIDTH - 1),
		18546 => to_unsigned(32066, LUT_AMPL_WIDTH - 1),
		18547 => to_unsigned(32065, LUT_AMPL_WIDTH - 1),
		18548 => to_unsigned(32064, LUT_AMPL_WIDTH - 1),
		18549 => to_unsigned(32064, LUT_AMPL_WIDTH - 1),
		18550 => to_unsigned(32063, LUT_AMPL_WIDTH - 1),
		18551 => to_unsigned(32062, LUT_AMPL_WIDTH - 1),
		18552 => to_unsigned(32062, LUT_AMPL_WIDTH - 1),
		18553 => to_unsigned(32061, LUT_AMPL_WIDTH - 1),
		18554 => to_unsigned(32060, LUT_AMPL_WIDTH - 1),
		18555 => to_unsigned(32060, LUT_AMPL_WIDTH - 1),
		18556 => to_unsigned(32059, LUT_AMPL_WIDTH - 1),
		18557 => to_unsigned(32058, LUT_AMPL_WIDTH - 1),
		18558 => to_unsigned(32058, LUT_AMPL_WIDTH - 1),
		18559 => to_unsigned(32057, LUT_AMPL_WIDTH - 1),
		18560 => to_unsigned(32057, LUT_AMPL_WIDTH - 1),
		18561 => to_unsigned(32056, LUT_AMPL_WIDTH - 1),
		18562 => to_unsigned(32055, LUT_AMPL_WIDTH - 1),
		18563 => to_unsigned(32055, LUT_AMPL_WIDTH - 1),
		18564 => to_unsigned(32054, LUT_AMPL_WIDTH - 1),
		18565 => to_unsigned(32053, LUT_AMPL_WIDTH - 1),
		18566 => to_unsigned(32053, LUT_AMPL_WIDTH - 1),
		18567 => to_unsigned(32052, LUT_AMPL_WIDTH - 1),
		18568 => to_unsigned(32051, LUT_AMPL_WIDTH - 1),
		18569 => to_unsigned(32051, LUT_AMPL_WIDTH - 1),
		18570 => to_unsigned(32050, LUT_AMPL_WIDTH - 1),
		18571 => to_unsigned(32049, LUT_AMPL_WIDTH - 1),
		18572 => to_unsigned(32049, LUT_AMPL_WIDTH - 1),
		18573 => to_unsigned(32048, LUT_AMPL_WIDTH - 1),
		18574 => to_unsigned(32047, LUT_AMPL_WIDTH - 1),
		18575 => to_unsigned(32047, LUT_AMPL_WIDTH - 1),
		18576 => to_unsigned(32046, LUT_AMPL_WIDTH - 1),
		18577 => to_unsigned(32045, LUT_AMPL_WIDTH - 1),
		18578 => to_unsigned(32045, LUT_AMPL_WIDTH - 1),
		18579 => to_unsigned(32044, LUT_AMPL_WIDTH - 1),
		18580 => to_unsigned(32043, LUT_AMPL_WIDTH - 1),
		18581 => to_unsigned(32043, LUT_AMPL_WIDTH - 1),
		18582 => to_unsigned(32042, LUT_AMPL_WIDTH - 1),
		18583 => to_unsigned(32041, LUT_AMPL_WIDTH - 1),
		18584 => to_unsigned(32041, LUT_AMPL_WIDTH - 1),
		18585 => to_unsigned(32040, LUT_AMPL_WIDTH - 1),
		18586 => to_unsigned(32040, LUT_AMPL_WIDTH - 1),
		18587 => to_unsigned(32039, LUT_AMPL_WIDTH - 1),
		18588 => to_unsigned(32038, LUT_AMPL_WIDTH - 1),
		18589 => to_unsigned(32038, LUT_AMPL_WIDTH - 1),
		18590 => to_unsigned(32037, LUT_AMPL_WIDTH - 1),
		18591 => to_unsigned(32036, LUT_AMPL_WIDTH - 1),
		18592 => to_unsigned(32036, LUT_AMPL_WIDTH - 1),
		18593 => to_unsigned(32035, LUT_AMPL_WIDTH - 1),
		18594 => to_unsigned(32034, LUT_AMPL_WIDTH - 1),
		18595 => to_unsigned(32034, LUT_AMPL_WIDTH - 1),
		18596 => to_unsigned(32033, LUT_AMPL_WIDTH - 1),
		18597 => to_unsigned(32032, LUT_AMPL_WIDTH - 1),
		18598 => to_unsigned(32032, LUT_AMPL_WIDTH - 1),
		18599 => to_unsigned(32031, LUT_AMPL_WIDTH - 1),
		18600 => to_unsigned(32030, LUT_AMPL_WIDTH - 1),
		18601 => to_unsigned(32030, LUT_AMPL_WIDTH - 1),
		18602 => to_unsigned(32029, LUT_AMPL_WIDTH - 1),
		18603 => to_unsigned(32028, LUT_AMPL_WIDTH - 1),
		18604 => to_unsigned(32028, LUT_AMPL_WIDTH - 1),
		18605 => to_unsigned(32027, LUT_AMPL_WIDTH - 1),
		18606 => to_unsigned(32026, LUT_AMPL_WIDTH - 1),
		18607 => to_unsigned(32026, LUT_AMPL_WIDTH - 1),
		18608 => to_unsigned(32025, LUT_AMPL_WIDTH - 1),
		18609 => to_unsigned(32024, LUT_AMPL_WIDTH - 1),
		18610 => to_unsigned(32024, LUT_AMPL_WIDTH - 1),
		18611 => to_unsigned(32023, LUT_AMPL_WIDTH - 1),
		18612 => to_unsigned(32022, LUT_AMPL_WIDTH - 1),
		18613 => to_unsigned(32022, LUT_AMPL_WIDTH - 1),
		18614 => to_unsigned(32021, LUT_AMPL_WIDTH - 1),
		18615 => to_unsigned(32020, LUT_AMPL_WIDTH - 1),
		18616 => to_unsigned(32020, LUT_AMPL_WIDTH - 1),
		18617 => to_unsigned(32019, LUT_AMPL_WIDTH - 1),
		18618 => to_unsigned(32018, LUT_AMPL_WIDTH - 1),
		18619 => to_unsigned(32018, LUT_AMPL_WIDTH - 1),
		18620 => to_unsigned(32017, LUT_AMPL_WIDTH - 1),
		18621 => to_unsigned(32016, LUT_AMPL_WIDTH - 1),
		18622 => to_unsigned(32016, LUT_AMPL_WIDTH - 1),
		18623 => to_unsigned(32015, LUT_AMPL_WIDTH - 1),
		18624 => to_unsigned(32014, LUT_AMPL_WIDTH - 1),
		18625 => to_unsigned(32014, LUT_AMPL_WIDTH - 1),
		18626 => to_unsigned(32013, LUT_AMPL_WIDTH - 1),
		18627 => to_unsigned(32012, LUT_AMPL_WIDTH - 1),
		18628 => to_unsigned(32012, LUT_AMPL_WIDTH - 1),
		18629 => to_unsigned(32011, LUT_AMPL_WIDTH - 1),
		18630 => to_unsigned(32010, LUT_AMPL_WIDTH - 1),
		18631 => to_unsigned(32010, LUT_AMPL_WIDTH - 1),
		18632 => to_unsigned(32009, LUT_AMPL_WIDTH - 1),
		18633 => to_unsigned(32008, LUT_AMPL_WIDTH - 1),
		18634 => to_unsigned(32008, LUT_AMPL_WIDTH - 1),
		18635 => to_unsigned(32007, LUT_AMPL_WIDTH - 1),
		18636 => to_unsigned(32006, LUT_AMPL_WIDTH - 1),
		18637 => to_unsigned(32006, LUT_AMPL_WIDTH - 1),
		18638 => to_unsigned(32005, LUT_AMPL_WIDTH - 1),
		18639 => to_unsigned(32004, LUT_AMPL_WIDTH - 1),
		18640 => to_unsigned(32004, LUT_AMPL_WIDTH - 1),
		18641 => to_unsigned(32003, LUT_AMPL_WIDTH - 1),
		18642 => to_unsigned(32002, LUT_AMPL_WIDTH - 1),
		18643 => to_unsigned(32002, LUT_AMPL_WIDTH - 1),
		18644 => to_unsigned(32001, LUT_AMPL_WIDTH - 1),
		18645 => to_unsigned(32000, LUT_AMPL_WIDTH - 1),
		18646 => to_unsigned(31999, LUT_AMPL_WIDTH - 1),
		18647 => to_unsigned(31999, LUT_AMPL_WIDTH - 1),
		18648 => to_unsigned(31998, LUT_AMPL_WIDTH - 1),
		18649 => to_unsigned(31997, LUT_AMPL_WIDTH - 1),
		18650 => to_unsigned(31997, LUT_AMPL_WIDTH - 1),
		18651 => to_unsigned(31996, LUT_AMPL_WIDTH - 1),
		18652 => to_unsigned(31995, LUT_AMPL_WIDTH - 1),
		18653 => to_unsigned(31995, LUT_AMPL_WIDTH - 1),
		18654 => to_unsigned(31994, LUT_AMPL_WIDTH - 1),
		18655 => to_unsigned(31993, LUT_AMPL_WIDTH - 1),
		18656 => to_unsigned(31993, LUT_AMPL_WIDTH - 1),
		18657 => to_unsigned(31992, LUT_AMPL_WIDTH - 1),
		18658 => to_unsigned(31991, LUT_AMPL_WIDTH - 1),
		18659 => to_unsigned(31991, LUT_AMPL_WIDTH - 1),
		18660 => to_unsigned(31990, LUT_AMPL_WIDTH - 1),
		18661 => to_unsigned(31989, LUT_AMPL_WIDTH - 1),
		18662 => to_unsigned(31989, LUT_AMPL_WIDTH - 1),
		18663 => to_unsigned(31988, LUT_AMPL_WIDTH - 1),
		18664 => to_unsigned(31987, LUT_AMPL_WIDTH - 1),
		18665 => to_unsigned(31987, LUT_AMPL_WIDTH - 1),
		18666 => to_unsigned(31986, LUT_AMPL_WIDTH - 1),
		18667 => to_unsigned(31985, LUT_AMPL_WIDTH - 1),
		18668 => to_unsigned(31985, LUT_AMPL_WIDTH - 1),
		18669 => to_unsigned(31984, LUT_AMPL_WIDTH - 1),
		18670 => to_unsigned(31983, LUT_AMPL_WIDTH - 1),
		18671 => to_unsigned(31982, LUT_AMPL_WIDTH - 1),
		18672 => to_unsigned(31982, LUT_AMPL_WIDTH - 1),
		18673 => to_unsigned(31981, LUT_AMPL_WIDTH - 1),
		18674 => to_unsigned(31980, LUT_AMPL_WIDTH - 1),
		18675 => to_unsigned(31980, LUT_AMPL_WIDTH - 1),
		18676 => to_unsigned(31979, LUT_AMPL_WIDTH - 1),
		18677 => to_unsigned(31978, LUT_AMPL_WIDTH - 1),
		18678 => to_unsigned(31978, LUT_AMPL_WIDTH - 1),
		18679 => to_unsigned(31977, LUT_AMPL_WIDTH - 1),
		18680 => to_unsigned(31976, LUT_AMPL_WIDTH - 1),
		18681 => to_unsigned(31976, LUT_AMPL_WIDTH - 1),
		18682 => to_unsigned(31975, LUT_AMPL_WIDTH - 1),
		18683 => to_unsigned(31974, LUT_AMPL_WIDTH - 1),
		18684 => to_unsigned(31974, LUT_AMPL_WIDTH - 1),
		18685 => to_unsigned(31973, LUT_AMPL_WIDTH - 1),
		18686 => to_unsigned(31972, LUT_AMPL_WIDTH - 1),
		18687 => to_unsigned(31972, LUT_AMPL_WIDTH - 1),
		18688 => to_unsigned(31971, LUT_AMPL_WIDTH - 1),
		18689 => to_unsigned(31970, LUT_AMPL_WIDTH - 1),
		18690 => to_unsigned(31969, LUT_AMPL_WIDTH - 1),
		18691 => to_unsigned(31969, LUT_AMPL_WIDTH - 1),
		18692 => to_unsigned(31968, LUT_AMPL_WIDTH - 1),
		18693 => to_unsigned(31967, LUT_AMPL_WIDTH - 1),
		18694 => to_unsigned(31967, LUT_AMPL_WIDTH - 1),
		18695 => to_unsigned(31966, LUT_AMPL_WIDTH - 1),
		18696 => to_unsigned(31965, LUT_AMPL_WIDTH - 1),
		18697 => to_unsigned(31965, LUT_AMPL_WIDTH - 1),
		18698 => to_unsigned(31964, LUT_AMPL_WIDTH - 1),
		18699 => to_unsigned(31963, LUT_AMPL_WIDTH - 1),
		18700 => to_unsigned(31963, LUT_AMPL_WIDTH - 1),
		18701 => to_unsigned(31962, LUT_AMPL_WIDTH - 1),
		18702 => to_unsigned(31961, LUT_AMPL_WIDTH - 1),
		18703 => to_unsigned(31960, LUT_AMPL_WIDTH - 1),
		18704 => to_unsigned(31960, LUT_AMPL_WIDTH - 1),
		18705 => to_unsigned(31959, LUT_AMPL_WIDTH - 1),
		18706 => to_unsigned(31958, LUT_AMPL_WIDTH - 1),
		18707 => to_unsigned(31958, LUT_AMPL_WIDTH - 1),
		18708 => to_unsigned(31957, LUT_AMPL_WIDTH - 1),
		18709 => to_unsigned(31956, LUT_AMPL_WIDTH - 1),
		18710 => to_unsigned(31956, LUT_AMPL_WIDTH - 1),
		18711 => to_unsigned(31955, LUT_AMPL_WIDTH - 1),
		18712 => to_unsigned(31954, LUT_AMPL_WIDTH - 1),
		18713 => to_unsigned(31954, LUT_AMPL_WIDTH - 1),
		18714 => to_unsigned(31953, LUT_AMPL_WIDTH - 1),
		18715 => to_unsigned(31952, LUT_AMPL_WIDTH - 1),
		18716 => to_unsigned(31951, LUT_AMPL_WIDTH - 1),
		18717 => to_unsigned(31951, LUT_AMPL_WIDTH - 1),
		18718 => to_unsigned(31950, LUT_AMPL_WIDTH - 1),
		18719 => to_unsigned(31949, LUT_AMPL_WIDTH - 1),
		18720 => to_unsigned(31949, LUT_AMPL_WIDTH - 1),
		18721 => to_unsigned(31948, LUT_AMPL_WIDTH - 1),
		18722 => to_unsigned(31947, LUT_AMPL_WIDTH - 1),
		18723 => to_unsigned(31947, LUT_AMPL_WIDTH - 1),
		18724 => to_unsigned(31946, LUT_AMPL_WIDTH - 1),
		18725 => to_unsigned(31945, LUT_AMPL_WIDTH - 1),
		18726 => to_unsigned(31944, LUT_AMPL_WIDTH - 1),
		18727 => to_unsigned(31944, LUT_AMPL_WIDTH - 1),
		18728 => to_unsigned(31943, LUT_AMPL_WIDTH - 1),
		18729 => to_unsigned(31942, LUT_AMPL_WIDTH - 1),
		18730 => to_unsigned(31942, LUT_AMPL_WIDTH - 1),
		18731 => to_unsigned(31941, LUT_AMPL_WIDTH - 1),
		18732 => to_unsigned(31940, LUT_AMPL_WIDTH - 1),
		18733 => to_unsigned(31940, LUT_AMPL_WIDTH - 1),
		18734 => to_unsigned(31939, LUT_AMPL_WIDTH - 1),
		18735 => to_unsigned(31938, LUT_AMPL_WIDTH - 1),
		18736 => to_unsigned(31937, LUT_AMPL_WIDTH - 1),
		18737 => to_unsigned(31937, LUT_AMPL_WIDTH - 1),
		18738 => to_unsigned(31936, LUT_AMPL_WIDTH - 1),
		18739 => to_unsigned(31935, LUT_AMPL_WIDTH - 1),
		18740 => to_unsigned(31935, LUT_AMPL_WIDTH - 1),
		18741 => to_unsigned(31934, LUT_AMPL_WIDTH - 1),
		18742 => to_unsigned(31933, LUT_AMPL_WIDTH - 1),
		18743 => to_unsigned(31933, LUT_AMPL_WIDTH - 1),
		18744 => to_unsigned(31932, LUT_AMPL_WIDTH - 1),
		18745 => to_unsigned(31931, LUT_AMPL_WIDTH - 1),
		18746 => to_unsigned(31930, LUT_AMPL_WIDTH - 1),
		18747 => to_unsigned(31930, LUT_AMPL_WIDTH - 1),
		18748 => to_unsigned(31929, LUT_AMPL_WIDTH - 1),
		18749 => to_unsigned(31928, LUT_AMPL_WIDTH - 1),
		18750 => to_unsigned(31928, LUT_AMPL_WIDTH - 1),
		18751 => to_unsigned(31927, LUT_AMPL_WIDTH - 1),
		18752 => to_unsigned(31926, LUT_AMPL_WIDTH - 1),
		18753 => to_unsigned(31925, LUT_AMPL_WIDTH - 1),
		18754 => to_unsigned(31925, LUT_AMPL_WIDTH - 1),
		18755 => to_unsigned(31924, LUT_AMPL_WIDTH - 1),
		18756 => to_unsigned(31923, LUT_AMPL_WIDTH - 1),
		18757 => to_unsigned(31923, LUT_AMPL_WIDTH - 1),
		18758 => to_unsigned(31922, LUT_AMPL_WIDTH - 1),
		18759 => to_unsigned(31921, LUT_AMPL_WIDTH - 1),
		18760 => to_unsigned(31921, LUT_AMPL_WIDTH - 1),
		18761 => to_unsigned(31920, LUT_AMPL_WIDTH - 1),
		18762 => to_unsigned(31919, LUT_AMPL_WIDTH - 1),
		18763 => to_unsigned(31918, LUT_AMPL_WIDTH - 1),
		18764 => to_unsigned(31918, LUT_AMPL_WIDTH - 1),
		18765 => to_unsigned(31917, LUT_AMPL_WIDTH - 1),
		18766 => to_unsigned(31916, LUT_AMPL_WIDTH - 1),
		18767 => to_unsigned(31916, LUT_AMPL_WIDTH - 1),
		18768 => to_unsigned(31915, LUT_AMPL_WIDTH - 1),
		18769 => to_unsigned(31914, LUT_AMPL_WIDTH - 1),
		18770 => to_unsigned(31913, LUT_AMPL_WIDTH - 1),
		18771 => to_unsigned(31913, LUT_AMPL_WIDTH - 1),
		18772 => to_unsigned(31912, LUT_AMPL_WIDTH - 1),
		18773 => to_unsigned(31911, LUT_AMPL_WIDTH - 1),
		18774 => to_unsigned(31911, LUT_AMPL_WIDTH - 1),
		18775 => to_unsigned(31910, LUT_AMPL_WIDTH - 1),
		18776 => to_unsigned(31909, LUT_AMPL_WIDTH - 1),
		18777 => to_unsigned(31908, LUT_AMPL_WIDTH - 1),
		18778 => to_unsigned(31908, LUT_AMPL_WIDTH - 1),
		18779 => to_unsigned(31907, LUT_AMPL_WIDTH - 1),
		18780 => to_unsigned(31906, LUT_AMPL_WIDTH - 1),
		18781 => to_unsigned(31906, LUT_AMPL_WIDTH - 1),
		18782 => to_unsigned(31905, LUT_AMPL_WIDTH - 1),
		18783 => to_unsigned(31904, LUT_AMPL_WIDTH - 1),
		18784 => to_unsigned(31903, LUT_AMPL_WIDTH - 1),
		18785 => to_unsigned(31903, LUT_AMPL_WIDTH - 1),
		18786 => to_unsigned(31902, LUT_AMPL_WIDTH - 1),
		18787 => to_unsigned(31901, LUT_AMPL_WIDTH - 1),
		18788 => to_unsigned(31901, LUT_AMPL_WIDTH - 1),
		18789 => to_unsigned(31900, LUT_AMPL_WIDTH - 1),
		18790 => to_unsigned(31899, LUT_AMPL_WIDTH - 1),
		18791 => to_unsigned(31898, LUT_AMPL_WIDTH - 1),
		18792 => to_unsigned(31898, LUT_AMPL_WIDTH - 1),
		18793 => to_unsigned(31897, LUT_AMPL_WIDTH - 1),
		18794 => to_unsigned(31896, LUT_AMPL_WIDTH - 1),
		18795 => to_unsigned(31896, LUT_AMPL_WIDTH - 1),
		18796 => to_unsigned(31895, LUT_AMPL_WIDTH - 1),
		18797 => to_unsigned(31894, LUT_AMPL_WIDTH - 1),
		18798 => to_unsigned(31893, LUT_AMPL_WIDTH - 1),
		18799 => to_unsigned(31893, LUT_AMPL_WIDTH - 1),
		18800 => to_unsigned(31892, LUT_AMPL_WIDTH - 1),
		18801 => to_unsigned(31891, LUT_AMPL_WIDTH - 1),
		18802 => to_unsigned(31890, LUT_AMPL_WIDTH - 1),
		18803 => to_unsigned(31890, LUT_AMPL_WIDTH - 1),
		18804 => to_unsigned(31889, LUT_AMPL_WIDTH - 1),
		18805 => to_unsigned(31888, LUT_AMPL_WIDTH - 1),
		18806 => to_unsigned(31888, LUT_AMPL_WIDTH - 1),
		18807 => to_unsigned(31887, LUT_AMPL_WIDTH - 1),
		18808 => to_unsigned(31886, LUT_AMPL_WIDTH - 1),
		18809 => to_unsigned(31885, LUT_AMPL_WIDTH - 1),
		18810 => to_unsigned(31885, LUT_AMPL_WIDTH - 1),
		18811 => to_unsigned(31884, LUT_AMPL_WIDTH - 1),
		18812 => to_unsigned(31883, LUT_AMPL_WIDTH - 1),
		18813 => to_unsigned(31882, LUT_AMPL_WIDTH - 1),
		18814 => to_unsigned(31882, LUT_AMPL_WIDTH - 1),
		18815 => to_unsigned(31881, LUT_AMPL_WIDTH - 1),
		18816 => to_unsigned(31880, LUT_AMPL_WIDTH - 1),
		18817 => to_unsigned(31880, LUT_AMPL_WIDTH - 1),
		18818 => to_unsigned(31879, LUT_AMPL_WIDTH - 1),
		18819 => to_unsigned(31878, LUT_AMPL_WIDTH - 1),
		18820 => to_unsigned(31877, LUT_AMPL_WIDTH - 1),
		18821 => to_unsigned(31877, LUT_AMPL_WIDTH - 1),
		18822 => to_unsigned(31876, LUT_AMPL_WIDTH - 1),
		18823 => to_unsigned(31875, LUT_AMPL_WIDTH - 1),
		18824 => to_unsigned(31875, LUT_AMPL_WIDTH - 1),
		18825 => to_unsigned(31874, LUT_AMPL_WIDTH - 1),
		18826 => to_unsigned(31873, LUT_AMPL_WIDTH - 1),
		18827 => to_unsigned(31872, LUT_AMPL_WIDTH - 1),
		18828 => to_unsigned(31872, LUT_AMPL_WIDTH - 1),
		18829 => to_unsigned(31871, LUT_AMPL_WIDTH - 1),
		18830 => to_unsigned(31870, LUT_AMPL_WIDTH - 1),
		18831 => to_unsigned(31869, LUT_AMPL_WIDTH - 1),
		18832 => to_unsigned(31869, LUT_AMPL_WIDTH - 1),
		18833 => to_unsigned(31868, LUT_AMPL_WIDTH - 1),
		18834 => to_unsigned(31867, LUT_AMPL_WIDTH - 1),
		18835 => to_unsigned(31866, LUT_AMPL_WIDTH - 1),
		18836 => to_unsigned(31866, LUT_AMPL_WIDTH - 1),
		18837 => to_unsigned(31865, LUT_AMPL_WIDTH - 1),
		18838 => to_unsigned(31864, LUT_AMPL_WIDTH - 1),
		18839 => to_unsigned(31864, LUT_AMPL_WIDTH - 1),
		18840 => to_unsigned(31863, LUT_AMPL_WIDTH - 1),
		18841 => to_unsigned(31862, LUT_AMPL_WIDTH - 1),
		18842 => to_unsigned(31861, LUT_AMPL_WIDTH - 1),
		18843 => to_unsigned(31861, LUT_AMPL_WIDTH - 1),
		18844 => to_unsigned(31860, LUT_AMPL_WIDTH - 1),
		18845 => to_unsigned(31859, LUT_AMPL_WIDTH - 1),
		18846 => to_unsigned(31858, LUT_AMPL_WIDTH - 1),
		18847 => to_unsigned(31858, LUT_AMPL_WIDTH - 1),
		18848 => to_unsigned(31857, LUT_AMPL_WIDTH - 1),
		18849 => to_unsigned(31856, LUT_AMPL_WIDTH - 1),
		18850 => to_unsigned(31855, LUT_AMPL_WIDTH - 1),
		18851 => to_unsigned(31855, LUT_AMPL_WIDTH - 1),
		18852 => to_unsigned(31854, LUT_AMPL_WIDTH - 1),
		18853 => to_unsigned(31853, LUT_AMPL_WIDTH - 1),
		18854 => to_unsigned(31853, LUT_AMPL_WIDTH - 1),
		18855 => to_unsigned(31852, LUT_AMPL_WIDTH - 1),
		18856 => to_unsigned(31851, LUT_AMPL_WIDTH - 1),
		18857 => to_unsigned(31850, LUT_AMPL_WIDTH - 1),
		18858 => to_unsigned(31850, LUT_AMPL_WIDTH - 1),
		18859 => to_unsigned(31849, LUT_AMPL_WIDTH - 1),
		18860 => to_unsigned(31848, LUT_AMPL_WIDTH - 1),
		18861 => to_unsigned(31847, LUT_AMPL_WIDTH - 1),
		18862 => to_unsigned(31847, LUT_AMPL_WIDTH - 1),
		18863 => to_unsigned(31846, LUT_AMPL_WIDTH - 1),
		18864 => to_unsigned(31845, LUT_AMPL_WIDTH - 1),
		18865 => to_unsigned(31844, LUT_AMPL_WIDTH - 1),
		18866 => to_unsigned(31844, LUT_AMPL_WIDTH - 1),
		18867 => to_unsigned(31843, LUT_AMPL_WIDTH - 1),
		18868 => to_unsigned(31842, LUT_AMPL_WIDTH - 1),
		18869 => to_unsigned(31841, LUT_AMPL_WIDTH - 1),
		18870 => to_unsigned(31841, LUT_AMPL_WIDTH - 1),
		18871 => to_unsigned(31840, LUT_AMPL_WIDTH - 1),
		18872 => to_unsigned(31839, LUT_AMPL_WIDTH - 1),
		18873 => to_unsigned(31838, LUT_AMPL_WIDTH - 1),
		18874 => to_unsigned(31838, LUT_AMPL_WIDTH - 1),
		18875 => to_unsigned(31837, LUT_AMPL_WIDTH - 1),
		18876 => to_unsigned(31836, LUT_AMPL_WIDTH - 1),
		18877 => to_unsigned(31836, LUT_AMPL_WIDTH - 1),
		18878 => to_unsigned(31835, LUT_AMPL_WIDTH - 1),
		18879 => to_unsigned(31834, LUT_AMPL_WIDTH - 1),
		18880 => to_unsigned(31833, LUT_AMPL_WIDTH - 1),
		18881 => to_unsigned(31833, LUT_AMPL_WIDTH - 1),
		18882 => to_unsigned(31832, LUT_AMPL_WIDTH - 1),
		18883 => to_unsigned(31831, LUT_AMPL_WIDTH - 1),
		18884 => to_unsigned(31830, LUT_AMPL_WIDTH - 1),
		18885 => to_unsigned(31830, LUT_AMPL_WIDTH - 1),
		18886 => to_unsigned(31829, LUT_AMPL_WIDTH - 1),
		18887 => to_unsigned(31828, LUT_AMPL_WIDTH - 1),
		18888 => to_unsigned(31827, LUT_AMPL_WIDTH - 1),
		18889 => to_unsigned(31827, LUT_AMPL_WIDTH - 1),
		18890 => to_unsigned(31826, LUT_AMPL_WIDTH - 1),
		18891 => to_unsigned(31825, LUT_AMPL_WIDTH - 1),
		18892 => to_unsigned(31824, LUT_AMPL_WIDTH - 1),
		18893 => to_unsigned(31824, LUT_AMPL_WIDTH - 1),
		18894 => to_unsigned(31823, LUT_AMPL_WIDTH - 1),
		18895 => to_unsigned(31822, LUT_AMPL_WIDTH - 1),
		18896 => to_unsigned(31821, LUT_AMPL_WIDTH - 1),
		18897 => to_unsigned(31821, LUT_AMPL_WIDTH - 1),
		18898 => to_unsigned(31820, LUT_AMPL_WIDTH - 1),
		18899 => to_unsigned(31819, LUT_AMPL_WIDTH - 1),
		18900 => to_unsigned(31818, LUT_AMPL_WIDTH - 1),
		18901 => to_unsigned(31818, LUT_AMPL_WIDTH - 1),
		18902 => to_unsigned(31817, LUT_AMPL_WIDTH - 1),
		18903 => to_unsigned(31816, LUT_AMPL_WIDTH - 1),
		18904 => to_unsigned(31815, LUT_AMPL_WIDTH - 1),
		18905 => to_unsigned(31815, LUT_AMPL_WIDTH - 1),
		18906 => to_unsigned(31814, LUT_AMPL_WIDTH - 1),
		18907 => to_unsigned(31813, LUT_AMPL_WIDTH - 1),
		18908 => to_unsigned(31812, LUT_AMPL_WIDTH - 1),
		18909 => to_unsigned(31812, LUT_AMPL_WIDTH - 1),
		18910 => to_unsigned(31811, LUT_AMPL_WIDTH - 1),
		18911 => to_unsigned(31810, LUT_AMPL_WIDTH - 1),
		18912 => to_unsigned(31809, LUT_AMPL_WIDTH - 1),
		18913 => to_unsigned(31809, LUT_AMPL_WIDTH - 1),
		18914 => to_unsigned(31808, LUT_AMPL_WIDTH - 1),
		18915 => to_unsigned(31807, LUT_AMPL_WIDTH - 1),
		18916 => to_unsigned(31806, LUT_AMPL_WIDTH - 1),
		18917 => to_unsigned(31806, LUT_AMPL_WIDTH - 1),
		18918 => to_unsigned(31805, LUT_AMPL_WIDTH - 1),
		18919 => to_unsigned(31804, LUT_AMPL_WIDTH - 1),
		18920 => to_unsigned(31803, LUT_AMPL_WIDTH - 1),
		18921 => to_unsigned(31802, LUT_AMPL_WIDTH - 1),
		18922 => to_unsigned(31802, LUT_AMPL_WIDTH - 1),
		18923 => to_unsigned(31801, LUT_AMPL_WIDTH - 1),
		18924 => to_unsigned(31800, LUT_AMPL_WIDTH - 1),
		18925 => to_unsigned(31799, LUT_AMPL_WIDTH - 1),
		18926 => to_unsigned(31799, LUT_AMPL_WIDTH - 1),
		18927 => to_unsigned(31798, LUT_AMPL_WIDTH - 1),
		18928 => to_unsigned(31797, LUT_AMPL_WIDTH - 1),
		18929 => to_unsigned(31796, LUT_AMPL_WIDTH - 1),
		18930 => to_unsigned(31796, LUT_AMPL_WIDTH - 1),
		18931 => to_unsigned(31795, LUT_AMPL_WIDTH - 1),
		18932 => to_unsigned(31794, LUT_AMPL_WIDTH - 1),
		18933 => to_unsigned(31793, LUT_AMPL_WIDTH - 1),
		18934 => to_unsigned(31793, LUT_AMPL_WIDTH - 1),
		18935 => to_unsigned(31792, LUT_AMPL_WIDTH - 1),
		18936 => to_unsigned(31791, LUT_AMPL_WIDTH - 1),
		18937 => to_unsigned(31790, LUT_AMPL_WIDTH - 1),
		18938 => to_unsigned(31790, LUT_AMPL_WIDTH - 1),
		18939 => to_unsigned(31789, LUT_AMPL_WIDTH - 1),
		18940 => to_unsigned(31788, LUT_AMPL_WIDTH - 1),
		18941 => to_unsigned(31787, LUT_AMPL_WIDTH - 1),
		18942 => to_unsigned(31787, LUT_AMPL_WIDTH - 1),
		18943 => to_unsigned(31786, LUT_AMPL_WIDTH - 1),
		18944 => to_unsigned(31785, LUT_AMPL_WIDTH - 1),
		18945 => to_unsigned(31784, LUT_AMPL_WIDTH - 1),
		18946 => to_unsigned(31783, LUT_AMPL_WIDTH - 1),
		18947 => to_unsigned(31783, LUT_AMPL_WIDTH - 1),
		18948 => to_unsigned(31782, LUT_AMPL_WIDTH - 1),
		18949 => to_unsigned(31781, LUT_AMPL_WIDTH - 1),
		18950 => to_unsigned(31780, LUT_AMPL_WIDTH - 1),
		18951 => to_unsigned(31780, LUT_AMPL_WIDTH - 1),
		18952 => to_unsigned(31779, LUT_AMPL_WIDTH - 1),
		18953 => to_unsigned(31778, LUT_AMPL_WIDTH - 1),
		18954 => to_unsigned(31777, LUT_AMPL_WIDTH - 1),
		18955 => to_unsigned(31777, LUT_AMPL_WIDTH - 1),
		18956 => to_unsigned(31776, LUT_AMPL_WIDTH - 1),
		18957 => to_unsigned(31775, LUT_AMPL_WIDTH - 1),
		18958 => to_unsigned(31774, LUT_AMPL_WIDTH - 1),
		18959 => to_unsigned(31774, LUT_AMPL_WIDTH - 1),
		18960 => to_unsigned(31773, LUT_AMPL_WIDTH - 1),
		18961 => to_unsigned(31772, LUT_AMPL_WIDTH - 1),
		18962 => to_unsigned(31771, LUT_AMPL_WIDTH - 1),
		18963 => to_unsigned(31770, LUT_AMPL_WIDTH - 1),
		18964 => to_unsigned(31770, LUT_AMPL_WIDTH - 1),
		18965 => to_unsigned(31769, LUT_AMPL_WIDTH - 1),
		18966 => to_unsigned(31768, LUT_AMPL_WIDTH - 1),
		18967 => to_unsigned(31767, LUT_AMPL_WIDTH - 1),
		18968 => to_unsigned(31767, LUT_AMPL_WIDTH - 1),
		18969 => to_unsigned(31766, LUT_AMPL_WIDTH - 1),
		18970 => to_unsigned(31765, LUT_AMPL_WIDTH - 1),
		18971 => to_unsigned(31764, LUT_AMPL_WIDTH - 1),
		18972 => to_unsigned(31764, LUT_AMPL_WIDTH - 1),
		18973 => to_unsigned(31763, LUT_AMPL_WIDTH - 1),
		18974 => to_unsigned(31762, LUT_AMPL_WIDTH - 1),
		18975 => to_unsigned(31761, LUT_AMPL_WIDTH - 1),
		18976 => to_unsigned(31760, LUT_AMPL_WIDTH - 1),
		18977 => to_unsigned(31760, LUT_AMPL_WIDTH - 1),
		18978 => to_unsigned(31759, LUT_AMPL_WIDTH - 1),
		18979 => to_unsigned(31758, LUT_AMPL_WIDTH - 1),
		18980 => to_unsigned(31757, LUT_AMPL_WIDTH - 1),
		18981 => to_unsigned(31757, LUT_AMPL_WIDTH - 1),
		18982 => to_unsigned(31756, LUT_AMPL_WIDTH - 1),
		18983 => to_unsigned(31755, LUT_AMPL_WIDTH - 1),
		18984 => to_unsigned(31754, LUT_AMPL_WIDTH - 1),
		18985 => to_unsigned(31753, LUT_AMPL_WIDTH - 1),
		18986 => to_unsigned(31753, LUT_AMPL_WIDTH - 1),
		18987 => to_unsigned(31752, LUT_AMPL_WIDTH - 1),
		18988 => to_unsigned(31751, LUT_AMPL_WIDTH - 1),
		18989 => to_unsigned(31750, LUT_AMPL_WIDTH - 1),
		18990 => to_unsigned(31750, LUT_AMPL_WIDTH - 1),
		18991 => to_unsigned(31749, LUT_AMPL_WIDTH - 1),
		18992 => to_unsigned(31748, LUT_AMPL_WIDTH - 1),
		18993 => to_unsigned(31747, LUT_AMPL_WIDTH - 1),
		18994 => to_unsigned(31746, LUT_AMPL_WIDTH - 1),
		18995 => to_unsigned(31746, LUT_AMPL_WIDTH - 1),
		18996 => to_unsigned(31745, LUT_AMPL_WIDTH - 1),
		18997 => to_unsigned(31744, LUT_AMPL_WIDTH - 1),
		18998 => to_unsigned(31743, LUT_AMPL_WIDTH - 1),
		18999 => to_unsigned(31743, LUT_AMPL_WIDTH - 1),
		19000 => to_unsigned(31742, LUT_AMPL_WIDTH - 1),
		19001 => to_unsigned(31741, LUT_AMPL_WIDTH - 1),
		19002 => to_unsigned(31740, LUT_AMPL_WIDTH - 1),
		19003 => to_unsigned(31739, LUT_AMPL_WIDTH - 1),
		19004 => to_unsigned(31739, LUT_AMPL_WIDTH - 1),
		19005 => to_unsigned(31738, LUT_AMPL_WIDTH - 1),
		19006 => to_unsigned(31737, LUT_AMPL_WIDTH - 1),
		19007 => to_unsigned(31736, LUT_AMPL_WIDTH - 1),
		19008 => to_unsigned(31736, LUT_AMPL_WIDTH - 1),
		19009 => to_unsigned(31735, LUT_AMPL_WIDTH - 1),
		19010 => to_unsigned(31734, LUT_AMPL_WIDTH - 1),
		19011 => to_unsigned(31733, LUT_AMPL_WIDTH - 1),
		19012 => to_unsigned(31732, LUT_AMPL_WIDTH - 1),
		19013 => to_unsigned(31732, LUT_AMPL_WIDTH - 1),
		19014 => to_unsigned(31731, LUT_AMPL_WIDTH - 1),
		19015 => to_unsigned(31730, LUT_AMPL_WIDTH - 1),
		19016 => to_unsigned(31729, LUT_AMPL_WIDTH - 1),
		19017 => to_unsigned(31729, LUT_AMPL_WIDTH - 1),
		19018 => to_unsigned(31728, LUT_AMPL_WIDTH - 1),
		19019 => to_unsigned(31727, LUT_AMPL_WIDTH - 1),
		19020 => to_unsigned(31726, LUT_AMPL_WIDTH - 1),
		19021 => to_unsigned(31725, LUT_AMPL_WIDTH - 1),
		19022 => to_unsigned(31725, LUT_AMPL_WIDTH - 1),
		19023 => to_unsigned(31724, LUT_AMPL_WIDTH - 1),
		19024 => to_unsigned(31723, LUT_AMPL_WIDTH - 1),
		19025 => to_unsigned(31722, LUT_AMPL_WIDTH - 1),
		19026 => to_unsigned(31721, LUT_AMPL_WIDTH - 1),
		19027 => to_unsigned(31721, LUT_AMPL_WIDTH - 1),
		19028 => to_unsigned(31720, LUT_AMPL_WIDTH - 1),
		19029 => to_unsigned(31719, LUT_AMPL_WIDTH - 1),
		19030 => to_unsigned(31718, LUT_AMPL_WIDTH - 1),
		19031 => to_unsigned(31718, LUT_AMPL_WIDTH - 1),
		19032 => to_unsigned(31717, LUT_AMPL_WIDTH - 1),
		19033 => to_unsigned(31716, LUT_AMPL_WIDTH - 1),
		19034 => to_unsigned(31715, LUT_AMPL_WIDTH - 1),
		19035 => to_unsigned(31714, LUT_AMPL_WIDTH - 1),
		19036 => to_unsigned(31714, LUT_AMPL_WIDTH - 1),
		19037 => to_unsigned(31713, LUT_AMPL_WIDTH - 1),
		19038 => to_unsigned(31712, LUT_AMPL_WIDTH - 1),
		19039 => to_unsigned(31711, LUT_AMPL_WIDTH - 1),
		19040 => to_unsigned(31710, LUT_AMPL_WIDTH - 1),
		19041 => to_unsigned(31710, LUT_AMPL_WIDTH - 1),
		19042 => to_unsigned(31709, LUT_AMPL_WIDTH - 1),
		19043 => to_unsigned(31708, LUT_AMPL_WIDTH - 1),
		19044 => to_unsigned(31707, LUT_AMPL_WIDTH - 1),
		19045 => to_unsigned(31706, LUT_AMPL_WIDTH - 1),
		19046 => to_unsigned(31706, LUT_AMPL_WIDTH - 1),
		19047 => to_unsigned(31705, LUT_AMPL_WIDTH - 1),
		19048 => to_unsigned(31704, LUT_AMPL_WIDTH - 1),
		19049 => to_unsigned(31703, LUT_AMPL_WIDTH - 1),
		19050 => to_unsigned(31702, LUT_AMPL_WIDTH - 1),
		19051 => to_unsigned(31702, LUT_AMPL_WIDTH - 1),
		19052 => to_unsigned(31701, LUT_AMPL_WIDTH - 1),
		19053 => to_unsigned(31700, LUT_AMPL_WIDTH - 1),
		19054 => to_unsigned(31699, LUT_AMPL_WIDTH - 1),
		19055 => to_unsigned(31698, LUT_AMPL_WIDTH - 1),
		19056 => to_unsigned(31698, LUT_AMPL_WIDTH - 1),
		19057 => to_unsigned(31697, LUT_AMPL_WIDTH - 1),
		19058 => to_unsigned(31696, LUT_AMPL_WIDTH - 1),
		19059 => to_unsigned(31695, LUT_AMPL_WIDTH - 1),
		19060 => to_unsigned(31695, LUT_AMPL_WIDTH - 1),
		19061 => to_unsigned(31694, LUT_AMPL_WIDTH - 1),
		19062 => to_unsigned(31693, LUT_AMPL_WIDTH - 1),
		19063 => to_unsigned(31692, LUT_AMPL_WIDTH - 1),
		19064 => to_unsigned(31691, LUT_AMPL_WIDTH - 1),
		19065 => to_unsigned(31691, LUT_AMPL_WIDTH - 1),
		19066 => to_unsigned(31690, LUT_AMPL_WIDTH - 1),
		19067 => to_unsigned(31689, LUT_AMPL_WIDTH - 1),
		19068 => to_unsigned(31688, LUT_AMPL_WIDTH - 1),
		19069 => to_unsigned(31687, LUT_AMPL_WIDTH - 1),
		19070 => to_unsigned(31687, LUT_AMPL_WIDTH - 1),
		19071 => to_unsigned(31686, LUT_AMPL_WIDTH - 1),
		19072 => to_unsigned(31685, LUT_AMPL_WIDTH - 1),
		19073 => to_unsigned(31684, LUT_AMPL_WIDTH - 1),
		19074 => to_unsigned(31683, LUT_AMPL_WIDTH - 1),
		19075 => to_unsigned(31683, LUT_AMPL_WIDTH - 1),
		19076 => to_unsigned(31682, LUT_AMPL_WIDTH - 1),
		19077 => to_unsigned(31681, LUT_AMPL_WIDTH - 1),
		19078 => to_unsigned(31680, LUT_AMPL_WIDTH - 1),
		19079 => to_unsigned(31679, LUT_AMPL_WIDTH - 1),
		19080 => to_unsigned(31679, LUT_AMPL_WIDTH - 1),
		19081 => to_unsigned(31678, LUT_AMPL_WIDTH - 1),
		19082 => to_unsigned(31677, LUT_AMPL_WIDTH - 1),
		19083 => to_unsigned(31676, LUT_AMPL_WIDTH - 1),
		19084 => to_unsigned(31675, LUT_AMPL_WIDTH - 1),
		19085 => to_unsigned(31674, LUT_AMPL_WIDTH - 1),
		19086 => to_unsigned(31674, LUT_AMPL_WIDTH - 1),
		19087 => to_unsigned(31673, LUT_AMPL_WIDTH - 1),
		19088 => to_unsigned(31672, LUT_AMPL_WIDTH - 1),
		19089 => to_unsigned(31671, LUT_AMPL_WIDTH - 1),
		19090 => to_unsigned(31670, LUT_AMPL_WIDTH - 1),
		19091 => to_unsigned(31670, LUT_AMPL_WIDTH - 1),
		19092 => to_unsigned(31669, LUT_AMPL_WIDTH - 1),
		19093 => to_unsigned(31668, LUT_AMPL_WIDTH - 1),
		19094 => to_unsigned(31667, LUT_AMPL_WIDTH - 1),
		19095 => to_unsigned(31666, LUT_AMPL_WIDTH - 1),
		19096 => to_unsigned(31666, LUT_AMPL_WIDTH - 1),
		19097 => to_unsigned(31665, LUT_AMPL_WIDTH - 1),
		19098 => to_unsigned(31664, LUT_AMPL_WIDTH - 1),
		19099 => to_unsigned(31663, LUT_AMPL_WIDTH - 1),
		19100 => to_unsigned(31662, LUT_AMPL_WIDTH - 1),
		19101 => to_unsigned(31662, LUT_AMPL_WIDTH - 1),
		19102 => to_unsigned(31661, LUT_AMPL_WIDTH - 1),
		19103 => to_unsigned(31660, LUT_AMPL_WIDTH - 1),
		19104 => to_unsigned(31659, LUT_AMPL_WIDTH - 1),
		19105 => to_unsigned(31658, LUT_AMPL_WIDTH - 1),
		19106 => to_unsigned(31658, LUT_AMPL_WIDTH - 1),
		19107 => to_unsigned(31657, LUT_AMPL_WIDTH - 1),
		19108 => to_unsigned(31656, LUT_AMPL_WIDTH - 1),
		19109 => to_unsigned(31655, LUT_AMPL_WIDTH - 1),
		19110 => to_unsigned(31654, LUT_AMPL_WIDTH - 1),
		19111 => to_unsigned(31653, LUT_AMPL_WIDTH - 1),
		19112 => to_unsigned(31653, LUT_AMPL_WIDTH - 1),
		19113 => to_unsigned(31652, LUT_AMPL_WIDTH - 1),
		19114 => to_unsigned(31651, LUT_AMPL_WIDTH - 1),
		19115 => to_unsigned(31650, LUT_AMPL_WIDTH - 1),
		19116 => to_unsigned(31649, LUT_AMPL_WIDTH - 1),
		19117 => to_unsigned(31649, LUT_AMPL_WIDTH - 1),
		19118 => to_unsigned(31648, LUT_AMPL_WIDTH - 1),
		19119 => to_unsigned(31647, LUT_AMPL_WIDTH - 1),
		19120 => to_unsigned(31646, LUT_AMPL_WIDTH - 1),
		19121 => to_unsigned(31645, LUT_AMPL_WIDTH - 1),
		19122 => to_unsigned(31645, LUT_AMPL_WIDTH - 1),
		19123 => to_unsigned(31644, LUT_AMPL_WIDTH - 1),
		19124 => to_unsigned(31643, LUT_AMPL_WIDTH - 1),
		19125 => to_unsigned(31642, LUT_AMPL_WIDTH - 1),
		19126 => to_unsigned(31641, LUT_AMPL_WIDTH - 1),
		19127 => to_unsigned(31640, LUT_AMPL_WIDTH - 1),
		19128 => to_unsigned(31640, LUT_AMPL_WIDTH - 1),
		19129 => to_unsigned(31639, LUT_AMPL_WIDTH - 1),
		19130 => to_unsigned(31638, LUT_AMPL_WIDTH - 1),
		19131 => to_unsigned(31637, LUT_AMPL_WIDTH - 1),
		19132 => to_unsigned(31636, LUT_AMPL_WIDTH - 1),
		19133 => to_unsigned(31636, LUT_AMPL_WIDTH - 1),
		19134 => to_unsigned(31635, LUT_AMPL_WIDTH - 1),
		19135 => to_unsigned(31634, LUT_AMPL_WIDTH - 1),
		19136 => to_unsigned(31633, LUT_AMPL_WIDTH - 1),
		19137 => to_unsigned(31632, LUT_AMPL_WIDTH - 1),
		19138 => to_unsigned(31631, LUT_AMPL_WIDTH - 1),
		19139 => to_unsigned(31631, LUT_AMPL_WIDTH - 1),
		19140 => to_unsigned(31630, LUT_AMPL_WIDTH - 1),
		19141 => to_unsigned(31629, LUT_AMPL_WIDTH - 1),
		19142 => to_unsigned(31628, LUT_AMPL_WIDTH - 1),
		19143 => to_unsigned(31627, LUT_AMPL_WIDTH - 1),
		19144 => to_unsigned(31627, LUT_AMPL_WIDTH - 1),
		19145 => to_unsigned(31626, LUT_AMPL_WIDTH - 1),
		19146 => to_unsigned(31625, LUT_AMPL_WIDTH - 1),
		19147 => to_unsigned(31624, LUT_AMPL_WIDTH - 1),
		19148 => to_unsigned(31623, LUT_AMPL_WIDTH - 1),
		19149 => to_unsigned(31622, LUT_AMPL_WIDTH - 1),
		19150 => to_unsigned(31622, LUT_AMPL_WIDTH - 1),
		19151 => to_unsigned(31621, LUT_AMPL_WIDTH - 1),
		19152 => to_unsigned(31620, LUT_AMPL_WIDTH - 1),
		19153 => to_unsigned(31619, LUT_AMPL_WIDTH - 1),
		19154 => to_unsigned(31618, LUT_AMPL_WIDTH - 1),
		19155 => to_unsigned(31617, LUT_AMPL_WIDTH - 1),
		19156 => to_unsigned(31617, LUT_AMPL_WIDTH - 1),
		19157 => to_unsigned(31616, LUT_AMPL_WIDTH - 1),
		19158 => to_unsigned(31615, LUT_AMPL_WIDTH - 1),
		19159 => to_unsigned(31614, LUT_AMPL_WIDTH - 1),
		19160 => to_unsigned(31613, LUT_AMPL_WIDTH - 1),
		19161 => to_unsigned(31613, LUT_AMPL_WIDTH - 1),
		19162 => to_unsigned(31612, LUT_AMPL_WIDTH - 1),
		19163 => to_unsigned(31611, LUT_AMPL_WIDTH - 1),
		19164 => to_unsigned(31610, LUT_AMPL_WIDTH - 1),
		19165 => to_unsigned(31609, LUT_AMPL_WIDTH - 1),
		19166 => to_unsigned(31608, LUT_AMPL_WIDTH - 1),
		19167 => to_unsigned(31608, LUT_AMPL_WIDTH - 1),
		19168 => to_unsigned(31607, LUT_AMPL_WIDTH - 1),
		19169 => to_unsigned(31606, LUT_AMPL_WIDTH - 1),
		19170 => to_unsigned(31605, LUT_AMPL_WIDTH - 1),
		19171 => to_unsigned(31604, LUT_AMPL_WIDTH - 1),
		19172 => to_unsigned(31603, LUT_AMPL_WIDTH - 1),
		19173 => to_unsigned(31603, LUT_AMPL_WIDTH - 1),
		19174 => to_unsigned(31602, LUT_AMPL_WIDTH - 1),
		19175 => to_unsigned(31601, LUT_AMPL_WIDTH - 1),
		19176 => to_unsigned(31600, LUT_AMPL_WIDTH - 1),
		19177 => to_unsigned(31599, LUT_AMPL_WIDTH - 1),
		19178 => to_unsigned(31598, LUT_AMPL_WIDTH - 1),
		19179 => to_unsigned(31598, LUT_AMPL_WIDTH - 1),
		19180 => to_unsigned(31597, LUT_AMPL_WIDTH - 1),
		19181 => to_unsigned(31596, LUT_AMPL_WIDTH - 1),
		19182 => to_unsigned(31595, LUT_AMPL_WIDTH - 1),
		19183 => to_unsigned(31594, LUT_AMPL_WIDTH - 1),
		19184 => to_unsigned(31593, LUT_AMPL_WIDTH - 1),
		19185 => to_unsigned(31593, LUT_AMPL_WIDTH - 1),
		19186 => to_unsigned(31592, LUT_AMPL_WIDTH - 1),
		19187 => to_unsigned(31591, LUT_AMPL_WIDTH - 1),
		19188 => to_unsigned(31590, LUT_AMPL_WIDTH - 1),
		19189 => to_unsigned(31589, LUT_AMPL_WIDTH - 1),
		19190 => to_unsigned(31588, LUT_AMPL_WIDTH - 1),
		19191 => to_unsigned(31588, LUT_AMPL_WIDTH - 1),
		19192 => to_unsigned(31587, LUT_AMPL_WIDTH - 1),
		19193 => to_unsigned(31586, LUT_AMPL_WIDTH - 1),
		19194 => to_unsigned(31585, LUT_AMPL_WIDTH - 1),
		19195 => to_unsigned(31584, LUT_AMPL_WIDTH - 1),
		19196 => to_unsigned(31583, LUT_AMPL_WIDTH - 1),
		19197 => to_unsigned(31583, LUT_AMPL_WIDTH - 1),
		19198 => to_unsigned(31582, LUT_AMPL_WIDTH - 1),
		19199 => to_unsigned(31581, LUT_AMPL_WIDTH - 1),
		19200 => to_unsigned(31580, LUT_AMPL_WIDTH - 1),
		19201 => to_unsigned(31579, LUT_AMPL_WIDTH - 1),
		19202 => to_unsigned(31578, LUT_AMPL_WIDTH - 1),
		19203 => to_unsigned(31578, LUT_AMPL_WIDTH - 1),
		19204 => to_unsigned(31577, LUT_AMPL_WIDTH - 1),
		19205 => to_unsigned(31576, LUT_AMPL_WIDTH - 1),
		19206 => to_unsigned(31575, LUT_AMPL_WIDTH - 1),
		19207 => to_unsigned(31574, LUT_AMPL_WIDTH - 1),
		19208 => to_unsigned(31573, LUT_AMPL_WIDTH - 1),
		19209 => to_unsigned(31572, LUT_AMPL_WIDTH - 1),
		19210 => to_unsigned(31572, LUT_AMPL_WIDTH - 1),
		19211 => to_unsigned(31571, LUT_AMPL_WIDTH - 1),
		19212 => to_unsigned(31570, LUT_AMPL_WIDTH - 1),
		19213 => to_unsigned(31569, LUT_AMPL_WIDTH - 1),
		19214 => to_unsigned(31568, LUT_AMPL_WIDTH - 1),
		19215 => to_unsigned(31567, LUT_AMPL_WIDTH - 1),
		19216 => to_unsigned(31567, LUT_AMPL_WIDTH - 1),
		19217 => to_unsigned(31566, LUT_AMPL_WIDTH - 1),
		19218 => to_unsigned(31565, LUT_AMPL_WIDTH - 1),
		19219 => to_unsigned(31564, LUT_AMPL_WIDTH - 1),
		19220 => to_unsigned(31563, LUT_AMPL_WIDTH - 1),
		19221 => to_unsigned(31562, LUT_AMPL_WIDTH - 1),
		19222 => to_unsigned(31562, LUT_AMPL_WIDTH - 1),
		19223 => to_unsigned(31561, LUT_AMPL_WIDTH - 1),
		19224 => to_unsigned(31560, LUT_AMPL_WIDTH - 1),
		19225 => to_unsigned(31559, LUT_AMPL_WIDTH - 1),
		19226 => to_unsigned(31558, LUT_AMPL_WIDTH - 1),
		19227 => to_unsigned(31557, LUT_AMPL_WIDTH - 1),
		19228 => to_unsigned(31556, LUT_AMPL_WIDTH - 1),
		19229 => to_unsigned(31556, LUT_AMPL_WIDTH - 1),
		19230 => to_unsigned(31555, LUT_AMPL_WIDTH - 1),
		19231 => to_unsigned(31554, LUT_AMPL_WIDTH - 1),
		19232 => to_unsigned(31553, LUT_AMPL_WIDTH - 1),
		19233 => to_unsigned(31552, LUT_AMPL_WIDTH - 1),
		19234 => to_unsigned(31551, LUT_AMPL_WIDTH - 1),
		19235 => to_unsigned(31551, LUT_AMPL_WIDTH - 1),
		19236 => to_unsigned(31550, LUT_AMPL_WIDTH - 1),
		19237 => to_unsigned(31549, LUT_AMPL_WIDTH - 1),
		19238 => to_unsigned(31548, LUT_AMPL_WIDTH - 1),
		19239 => to_unsigned(31547, LUT_AMPL_WIDTH - 1),
		19240 => to_unsigned(31546, LUT_AMPL_WIDTH - 1),
		19241 => to_unsigned(31545, LUT_AMPL_WIDTH - 1),
		19242 => to_unsigned(31545, LUT_AMPL_WIDTH - 1),
		19243 => to_unsigned(31544, LUT_AMPL_WIDTH - 1),
		19244 => to_unsigned(31543, LUT_AMPL_WIDTH - 1),
		19245 => to_unsigned(31542, LUT_AMPL_WIDTH - 1),
		19246 => to_unsigned(31541, LUT_AMPL_WIDTH - 1),
		19247 => to_unsigned(31540, LUT_AMPL_WIDTH - 1),
		19248 => to_unsigned(31539, LUT_AMPL_WIDTH - 1),
		19249 => to_unsigned(31539, LUT_AMPL_WIDTH - 1),
		19250 => to_unsigned(31538, LUT_AMPL_WIDTH - 1),
		19251 => to_unsigned(31537, LUT_AMPL_WIDTH - 1),
		19252 => to_unsigned(31536, LUT_AMPL_WIDTH - 1),
		19253 => to_unsigned(31535, LUT_AMPL_WIDTH - 1),
		19254 => to_unsigned(31534, LUT_AMPL_WIDTH - 1),
		19255 => to_unsigned(31534, LUT_AMPL_WIDTH - 1),
		19256 => to_unsigned(31533, LUT_AMPL_WIDTH - 1),
		19257 => to_unsigned(31532, LUT_AMPL_WIDTH - 1),
		19258 => to_unsigned(31531, LUT_AMPL_WIDTH - 1),
		19259 => to_unsigned(31530, LUT_AMPL_WIDTH - 1),
		19260 => to_unsigned(31529, LUT_AMPL_WIDTH - 1),
		19261 => to_unsigned(31528, LUT_AMPL_WIDTH - 1),
		19262 => to_unsigned(31528, LUT_AMPL_WIDTH - 1),
		19263 => to_unsigned(31527, LUT_AMPL_WIDTH - 1),
		19264 => to_unsigned(31526, LUT_AMPL_WIDTH - 1),
		19265 => to_unsigned(31525, LUT_AMPL_WIDTH - 1),
		19266 => to_unsigned(31524, LUT_AMPL_WIDTH - 1),
		19267 => to_unsigned(31523, LUT_AMPL_WIDTH - 1),
		19268 => to_unsigned(31522, LUT_AMPL_WIDTH - 1),
		19269 => to_unsigned(31522, LUT_AMPL_WIDTH - 1),
		19270 => to_unsigned(31521, LUT_AMPL_WIDTH - 1),
		19271 => to_unsigned(31520, LUT_AMPL_WIDTH - 1),
		19272 => to_unsigned(31519, LUT_AMPL_WIDTH - 1),
		19273 => to_unsigned(31518, LUT_AMPL_WIDTH - 1),
		19274 => to_unsigned(31517, LUT_AMPL_WIDTH - 1),
		19275 => to_unsigned(31516, LUT_AMPL_WIDTH - 1),
		19276 => to_unsigned(31516, LUT_AMPL_WIDTH - 1),
		19277 => to_unsigned(31515, LUT_AMPL_WIDTH - 1),
		19278 => to_unsigned(31514, LUT_AMPL_WIDTH - 1),
		19279 => to_unsigned(31513, LUT_AMPL_WIDTH - 1),
		19280 => to_unsigned(31512, LUT_AMPL_WIDTH - 1),
		19281 => to_unsigned(31511, LUT_AMPL_WIDTH - 1),
		19282 => to_unsigned(31510, LUT_AMPL_WIDTH - 1),
		19283 => to_unsigned(31510, LUT_AMPL_WIDTH - 1),
		19284 => to_unsigned(31509, LUT_AMPL_WIDTH - 1),
		19285 => to_unsigned(31508, LUT_AMPL_WIDTH - 1),
		19286 => to_unsigned(31507, LUT_AMPL_WIDTH - 1),
		19287 => to_unsigned(31506, LUT_AMPL_WIDTH - 1),
		19288 => to_unsigned(31505, LUT_AMPL_WIDTH - 1),
		19289 => to_unsigned(31504, LUT_AMPL_WIDTH - 1),
		19290 => to_unsigned(31503, LUT_AMPL_WIDTH - 1),
		19291 => to_unsigned(31503, LUT_AMPL_WIDTH - 1),
		19292 => to_unsigned(31502, LUT_AMPL_WIDTH - 1),
		19293 => to_unsigned(31501, LUT_AMPL_WIDTH - 1),
		19294 => to_unsigned(31500, LUT_AMPL_WIDTH - 1),
		19295 => to_unsigned(31499, LUT_AMPL_WIDTH - 1),
		19296 => to_unsigned(31498, LUT_AMPL_WIDTH - 1),
		19297 => to_unsigned(31497, LUT_AMPL_WIDTH - 1),
		19298 => to_unsigned(31497, LUT_AMPL_WIDTH - 1),
		19299 => to_unsigned(31496, LUT_AMPL_WIDTH - 1),
		19300 => to_unsigned(31495, LUT_AMPL_WIDTH - 1),
		19301 => to_unsigned(31494, LUT_AMPL_WIDTH - 1),
		19302 => to_unsigned(31493, LUT_AMPL_WIDTH - 1),
		19303 => to_unsigned(31492, LUT_AMPL_WIDTH - 1),
		19304 => to_unsigned(31491, LUT_AMPL_WIDTH - 1),
		19305 => to_unsigned(31490, LUT_AMPL_WIDTH - 1),
		19306 => to_unsigned(31490, LUT_AMPL_WIDTH - 1),
		19307 => to_unsigned(31489, LUT_AMPL_WIDTH - 1),
		19308 => to_unsigned(31488, LUT_AMPL_WIDTH - 1),
		19309 => to_unsigned(31487, LUT_AMPL_WIDTH - 1),
		19310 => to_unsigned(31486, LUT_AMPL_WIDTH - 1),
		19311 => to_unsigned(31485, LUT_AMPL_WIDTH - 1),
		19312 => to_unsigned(31484, LUT_AMPL_WIDTH - 1),
		19313 => to_unsigned(31484, LUT_AMPL_WIDTH - 1),
		19314 => to_unsigned(31483, LUT_AMPL_WIDTH - 1),
		19315 => to_unsigned(31482, LUT_AMPL_WIDTH - 1),
		19316 => to_unsigned(31481, LUT_AMPL_WIDTH - 1),
		19317 => to_unsigned(31480, LUT_AMPL_WIDTH - 1),
		19318 => to_unsigned(31479, LUT_AMPL_WIDTH - 1),
		19319 => to_unsigned(31478, LUT_AMPL_WIDTH - 1),
		19320 => to_unsigned(31477, LUT_AMPL_WIDTH - 1),
		19321 => to_unsigned(31477, LUT_AMPL_WIDTH - 1),
		19322 => to_unsigned(31476, LUT_AMPL_WIDTH - 1),
		19323 => to_unsigned(31475, LUT_AMPL_WIDTH - 1),
		19324 => to_unsigned(31474, LUT_AMPL_WIDTH - 1),
		19325 => to_unsigned(31473, LUT_AMPL_WIDTH - 1),
		19326 => to_unsigned(31472, LUT_AMPL_WIDTH - 1),
		19327 => to_unsigned(31471, LUT_AMPL_WIDTH - 1),
		19328 => to_unsigned(31470, LUT_AMPL_WIDTH - 1),
		19329 => to_unsigned(31470, LUT_AMPL_WIDTH - 1),
		19330 => to_unsigned(31469, LUT_AMPL_WIDTH - 1),
		19331 => to_unsigned(31468, LUT_AMPL_WIDTH - 1),
		19332 => to_unsigned(31467, LUT_AMPL_WIDTH - 1),
		19333 => to_unsigned(31466, LUT_AMPL_WIDTH - 1),
		19334 => to_unsigned(31465, LUT_AMPL_WIDTH - 1),
		19335 => to_unsigned(31464, LUT_AMPL_WIDTH - 1),
		19336 => to_unsigned(31463, LUT_AMPL_WIDTH - 1),
		19337 => to_unsigned(31463, LUT_AMPL_WIDTH - 1),
		19338 => to_unsigned(31462, LUT_AMPL_WIDTH - 1),
		19339 => to_unsigned(31461, LUT_AMPL_WIDTH - 1),
		19340 => to_unsigned(31460, LUT_AMPL_WIDTH - 1),
		19341 => to_unsigned(31459, LUT_AMPL_WIDTH - 1),
		19342 => to_unsigned(31458, LUT_AMPL_WIDTH - 1),
		19343 => to_unsigned(31457, LUT_AMPL_WIDTH - 1),
		19344 => to_unsigned(31456, LUT_AMPL_WIDTH - 1),
		19345 => to_unsigned(31456, LUT_AMPL_WIDTH - 1),
		19346 => to_unsigned(31455, LUT_AMPL_WIDTH - 1),
		19347 => to_unsigned(31454, LUT_AMPL_WIDTH - 1),
		19348 => to_unsigned(31453, LUT_AMPL_WIDTH - 1),
		19349 => to_unsigned(31452, LUT_AMPL_WIDTH - 1),
		19350 => to_unsigned(31451, LUT_AMPL_WIDTH - 1),
		19351 => to_unsigned(31450, LUT_AMPL_WIDTH - 1),
		19352 => to_unsigned(31449, LUT_AMPL_WIDTH - 1),
		19353 => to_unsigned(31448, LUT_AMPL_WIDTH - 1),
		19354 => to_unsigned(31448, LUT_AMPL_WIDTH - 1),
		19355 => to_unsigned(31447, LUT_AMPL_WIDTH - 1),
		19356 => to_unsigned(31446, LUT_AMPL_WIDTH - 1),
		19357 => to_unsigned(31445, LUT_AMPL_WIDTH - 1),
		19358 => to_unsigned(31444, LUT_AMPL_WIDTH - 1),
		19359 => to_unsigned(31443, LUT_AMPL_WIDTH - 1),
		19360 => to_unsigned(31442, LUT_AMPL_WIDTH - 1),
		19361 => to_unsigned(31441, LUT_AMPL_WIDTH - 1),
		19362 => to_unsigned(31441, LUT_AMPL_WIDTH - 1),
		19363 => to_unsigned(31440, LUT_AMPL_WIDTH - 1),
		19364 => to_unsigned(31439, LUT_AMPL_WIDTH - 1),
		19365 => to_unsigned(31438, LUT_AMPL_WIDTH - 1),
		19366 => to_unsigned(31437, LUT_AMPL_WIDTH - 1),
		19367 => to_unsigned(31436, LUT_AMPL_WIDTH - 1),
		19368 => to_unsigned(31435, LUT_AMPL_WIDTH - 1),
		19369 => to_unsigned(31434, LUT_AMPL_WIDTH - 1),
		19370 => to_unsigned(31433, LUT_AMPL_WIDTH - 1),
		19371 => to_unsigned(31433, LUT_AMPL_WIDTH - 1),
		19372 => to_unsigned(31432, LUT_AMPL_WIDTH - 1),
		19373 => to_unsigned(31431, LUT_AMPL_WIDTH - 1),
		19374 => to_unsigned(31430, LUT_AMPL_WIDTH - 1),
		19375 => to_unsigned(31429, LUT_AMPL_WIDTH - 1),
		19376 => to_unsigned(31428, LUT_AMPL_WIDTH - 1),
		19377 => to_unsigned(31427, LUT_AMPL_WIDTH - 1),
		19378 => to_unsigned(31426, LUT_AMPL_WIDTH - 1),
		19379 => to_unsigned(31425, LUT_AMPL_WIDTH - 1),
		19380 => to_unsigned(31425, LUT_AMPL_WIDTH - 1),
		19381 => to_unsigned(31424, LUT_AMPL_WIDTH - 1),
		19382 => to_unsigned(31423, LUT_AMPL_WIDTH - 1),
		19383 => to_unsigned(31422, LUT_AMPL_WIDTH - 1),
		19384 => to_unsigned(31421, LUT_AMPL_WIDTH - 1),
		19385 => to_unsigned(31420, LUT_AMPL_WIDTH - 1),
		19386 => to_unsigned(31419, LUT_AMPL_WIDTH - 1),
		19387 => to_unsigned(31418, LUT_AMPL_WIDTH - 1),
		19388 => to_unsigned(31417, LUT_AMPL_WIDTH - 1),
		19389 => to_unsigned(31417, LUT_AMPL_WIDTH - 1),
		19390 => to_unsigned(31416, LUT_AMPL_WIDTH - 1),
		19391 => to_unsigned(31415, LUT_AMPL_WIDTH - 1),
		19392 => to_unsigned(31414, LUT_AMPL_WIDTH - 1),
		19393 => to_unsigned(31413, LUT_AMPL_WIDTH - 1),
		19394 => to_unsigned(31412, LUT_AMPL_WIDTH - 1),
		19395 => to_unsigned(31411, LUT_AMPL_WIDTH - 1),
		19396 => to_unsigned(31410, LUT_AMPL_WIDTH - 1),
		19397 => to_unsigned(31409, LUT_AMPL_WIDTH - 1),
		19398 => to_unsigned(31408, LUT_AMPL_WIDTH - 1),
		19399 => to_unsigned(31408, LUT_AMPL_WIDTH - 1),
		19400 => to_unsigned(31407, LUT_AMPL_WIDTH - 1),
		19401 => to_unsigned(31406, LUT_AMPL_WIDTH - 1),
		19402 => to_unsigned(31405, LUT_AMPL_WIDTH - 1),
		19403 => to_unsigned(31404, LUT_AMPL_WIDTH - 1),
		19404 => to_unsigned(31403, LUT_AMPL_WIDTH - 1),
		19405 => to_unsigned(31402, LUT_AMPL_WIDTH - 1),
		19406 => to_unsigned(31401, LUT_AMPL_WIDTH - 1),
		19407 => to_unsigned(31400, LUT_AMPL_WIDTH - 1),
		19408 => to_unsigned(31400, LUT_AMPL_WIDTH - 1),
		19409 => to_unsigned(31399, LUT_AMPL_WIDTH - 1),
		19410 => to_unsigned(31398, LUT_AMPL_WIDTH - 1),
		19411 => to_unsigned(31397, LUT_AMPL_WIDTH - 1),
		19412 => to_unsigned(31396, LUT_AMPL_WIDTH - 1),
		19413 => to_unsigned(31395, LUT_AMPL_WIDTH - 1),
		19414 => to_unsigned(31394, LUT_AMPL_WIDTH - 1),
		19415 => to_unsigned(31393, LUT_AMPL_WIDTH - 1),
		19416 => to_unsigned(31392, LUT_AMPL_WIDTH - 1),
		19417 => to_unsigned(31391, LUT_AMPL_WIDTH - 1),
		19418 => to_unsigned(31391, LUT_AMPL_WIDTH - 1),
		19419 => to_unsigned(31390, LUT_AMPL_WIDTH - 1),
		19420 => to_unsigned(31389, LUT_AMPL_WIDTH - 1),
		19421 => to_unsigned(31388, LUT_AMPL_WIDTH - 1),
		19422 => to_unsigned(31387, LUT_AMPL_WIDTH - 1),
		19423 => to_unsigned(31386, LUT_AMPL_WIDTH - 1),
		19424 => to_unsigned(31385, LUT_AMPL_WIDTH - 1),
		19425 => to_unsigned(31384, LUT_AMPL_WIDTH - 1),
		19426 => to_unsigned(31383, LUT_AMPL_WIDTH - 1),
		19427 => to_unsigned(31382, LUT_AMPL_WIDTH - 1),
		19428 => to_unsigned(31381, LUT_AMPL_WIDTH - 1),
		19429 => to_unsigned(31381, LUT_AMPL_WIDTH - 1),
		19430 => to_unsigned(31380, LUT_AMPL_WIDTH - 1),
		19431 => to_unsigned(31379, LUT_AMPL_WIDTH - 1),
		19432 => to_unsigned(31378, LUT_AMPL_WIDTH - 1),
		19433 => to_unsigned(31377, LUT_AMPL_WIDTH - 1),
		19434 => to_unsigned(31376, LUT_AMPL_WIDTH - 1),
		19435 => to_unsigned(31375, LUT_AMPL_WIDTH - 1),
		19436 => to_unsigned(31374, LUT_AMPL_WIDTH - 1),
		19437 => to_unsigned(31373, LUT_AMPL_WIDTH - 1),
		19438 => to_unsigned(31372, LUT_AMPL_WIDTH - 1),
		19439 => to_unsigned(31372, LUT_AMPL_WIDTH - 1),
		19440 => to_unsigned(31371, LUT_AMPL_WIDTH - 1),
		19441 => to_unsigned(31370, LUT_AMPL_WIDTH - 1),
		19442 => to_unsigned(31369, LUT_AMPL_WIDTH - 1),
		19443 => to_unsigned(31368, LUT_AMPL_WIDTH - 1),
		19444 => to_unsigned(31367, LUT_AMPL_WIDTH - 1),
		19445 => to_unsigned(31366, LUT_AMPL_WIDTH - 1),
		19446 => to_unsigned(31365, LUT_AMPL_WIDTH - 1),
		19447 => to_unsigned(31364, LUT_AMPL_WIDTH - 1),
		19448 => to_unsigned(31363, LUT_AMPL_WIDTH - 1),
		19449 => to_unsigned(31362, LUT_AMPL_WIDTH - 1),
		19450 => to_unsigned(31362, LUT_AMPL_WIDTH - 1),
		19451 => to_unsigned(31361, LUT_AMPL_WIDTH - 1),
		19452 => to_unsigned(31360, LUT_AMPL_WIDTH - 1),
		19453 => to_unsigned(31359, LUT_AMPL_WIDTH - 1),
		19454 => to_unsigned(31358, LUT_AMPL_WIDTH - 1),
		19455 => to_unsigned(31357, LUT_AMPL_WIDTH - 1),
		19456 => to_unsigned(31356, LUT_AMPL_WIDTH - 1),
		19457 => to_unsigned(31355, LUT_AMPL_WIDTH - 1),
		19458 => to_unsigned(31354, LUT_AMPL_WIDTH - 1),
		19459 => to_unsigned(31353, LUT_AMPL_WIDTH - 1),
		19460 => to_unsigned(31352, LUT_AMPL_WIDTH - 1),
		19461 => to_unsigned(31352, LUT_AMPL_WIDTH - 1),
		19462 => to_unsigned(31351, LUT_AMPL_WIDTH - 1),
		19463 => to_unsigned(31350, LUT_AMPL_WIDTH - 1),
		19464 => to_unsigned(31349, LUT_AMPL_WIDTH - 1),
		19465 => to_unsigned(31348, LUT_AMPL_WIDTH - 1),
		19466 => to_unsigned(31347, LUT_AMPL_WIDTH - 1),
		19467 => to_unsigned(31346, LUT_AMPL_WIDTH - 1),
		19468 => to_unsigned(31345, LUT_AMPL_WIDTH - 1),
		19469 => to_unsigned(31344, LUT_AMPL_WIDTH - 1),
		19470 => to_unsigned(31343, LUT_AMPL_WIDTH - 1),
		19471 => to_unsigned(31342, LUT_AMPL_WIDTH - 1),
		19472 => to_unsigned(31341, LUT_AMPL_WIDTH - 1),
		19473 => to_unsigned(31341, LUT_AMPL_WIDTH - 1),
		19474 => to_unsigned(31340, LUT_AMPL_WIDTH - 1),
		19475 => to_unsigned(31339, LUT_AMPL_WIDTH - 1),
		19476 => to_unsigned(31338, LUT_AMPL_WIDTH - 1),
		19477 => to_unsigned(31337, LUT_AMPL_WIDTH - 1),
		19478 => to_unsigned(31336, LUT_AMPL_WIDTH - 1),
		19479 => to_unsigned(31335, LUT_AMPL_WIDTH - 1),
		19480 => to_unsigned(31334, LUT_AMPL_WIDTH - 1),
		19481 => to_unsigned(31333, LUT_AMPL_WIDTH - 1),
		19482 => to_unsigned(31332, LUT_AMPL_WIDTH - 1),
		19483 => to_unsigned(31331, LUT_AMPL_WIDTH - 1),
		19484 => to_unsigned(31330, LUT_AMPL_WIDTH - 1),
		19485 => to_unsigned(31329, LUT_AMPL_WIDTH - 1),
		19486 => to_unsigned(31329, LUT_AMPL_WIDTH - 1),
		19487 => to_unsigned(31328, LUT_AMPL_WIDTH - 1),
		19488 => to_unsigned(31327, LUT_AMPL_WIDTH - 1),
		19489 => to_unsigned(31326, LUT_AMPL_WIDTH - 1),
		19490 => to_unsigned(31325, LUT_AMPL_WIDTH - 1),
		19491 => to_unsigned(31324, LUT_AMPL_WIDTH - 1),
		19492 => to_unsigned(31323, LUT_AMPL_WIDTH - 1),
		19493 => to_unsigned(31322, LUT_AMPL_WIDTH - 1),
		19494 => to_unsigned(31321, LUT_AMPL_WIDTH - 1),
		19495 => to_unsigned(31320, LUT_AMPL_WIDTH - 1),
		19496 => to_unsigned(31319, LUT_AMPL_WIDTH - 1),
		19497 => to_unsigned(31318, LUT_AMPL_WIDTH - 1),
		19498 => to_unsigned(31318, LUT_AMPL_WIDTH - 1),
		19499 => to_unsigned(31317, LUT_AMPL_WIDTH - 1),
		19500 => to_unsigned(31316, LUT_AMPL_WIDTH - 1),
		19501 => to_unsigned(31315, LUT_AMPL_WIDTH - 1),
		19502 => to_unsigned(31314, LUT_AMPL_WIDTH - 1),
		19503 => to_unsigned(31313, LUT_AMPL_WIDTH - 1),
		19504 => to_unsigned(31312, LUT_AMPL_WIDTH - 1),
		19505 => to_unsigned(31311, LUT_AMPL_WIDTH - 1),
		19506 => to_unsigned(31310, LUT_AMPL_WIDTH - 1),
		19507 => to_unsigned(31309, LUT_AMPL_WIDTH - 1),
		19508 => to_unsigned(31308, LUT_AMPL_WIDTH - 1),
		19509 => to_unsigned(31307, LUT_AMPL_WIDTH - 1),
		19510 => to_unsigned(31306, LUT_AMPL_WIDTH - 1),
		19511 => to_unsigned(31305, LUT_AMPL_WIDTH - 1),
		19512 => to_unsigned(31305, LUT_AMPL_WIDTH - 1),
		19513 => to_unsigned(31304, LUT_AMPL_WIDTH - 1),
		19514 => to_unsigned(31303, LUT_AMPL_WIDTH - 1),
		19515 => to_unsigned(31302, LUT_AMPL_WIDTH - 1),
		19516 => to_unsigned(31301, LUT_AMPL_WIDTH - 1),
		19517 => to_unsigned(31300, LUT_AMPL_WIDTH - 1),
		19518 => to_unsigned(31299, LUT_AMPL_WIDTH - 1),
		19519 => to_unsigned(31298, LUT_AMPL_WIDTH - 1),
		19520 => to_unsigned(31297, LUT_AMPL_WIDTH - 1),
		19521 => to_unsigned(31296, LUT_AMPL_WIDTH - 1),
		19522 => to_unsigned(31295, LUT_AMPL_WIDTH - 1),
		19523 => to_unsigned(31294, LUT_AMPL_WIDTH - 1),
		19524 => to_unsigned(31293, LUT_AMPL_WIDTH - 1),
		19525 => to_unsigned(31292, LUT_AMPL_WIDTH - 1),
		19526 => to_unsigned(31292, LUT_AMPL_WIDTH - 1),
		19527 => to_unsigned(31291, LUT_AMPL_WIDTH - 1),
		19528 => to_unsigned(31290, LUT_AMPL_WIDTH - 1),
		19529 => to_unsigned(31289, LUT_AMPL_WIDTH - 1),
		19530 => to_unsigned(31288, LUT_AMPL_WIDTH - 1),
		19531 => to_unsigned(31287, LUT_AMPL_WIDTH - 1),
		19532 => to_unsigned(31286, LUT_AMPL_WIDTH - 1),
		19533 => to_unsigned(31285, LUT_AMPL_WIDTH - 1),
		19534 => to_unsigned(31284, LUT_AMPL_WIDTH - 1),
		19535 => to_unsigned(31283, LUT_AMPL_WIDTH - 1),
		19536 => to_unsigned(31282, LUT_AMPL_WIDTH - 1),
		19537 => to_unsigned(31281, LUT_AMPL_WIDTH - 1),
		19538 => to_unsigned(31280, LUT_AMPL_WIDTH - 1),
		19539 => to_unsigned(31279, LUT_AMPL_WIDTH - 1),
		19540 => to_unsigned(31278, LUT_AMPL_WIDTH - 1),
		19541 => to_unsigned(31278, LUT_AMPL_WIDTH - 1),
		19542 => to_unsigned(31277, LUT_AMPL_WIDTH - 1),
		19543 => to_unsigned(31276, LUT_AMPL_WIDTH - 1),
		19544 => to_unsigned(31275, LUT_AMPL_WIDTH - 1),
		19545 => to_unsigned(31274, LUT_AMPL_WIDTH - 1),
		19546 => to_unsigned(31273, LUT_AMPL_WIDTH - 1),
		19547 => to_unsigned(31272, LUT_AMPL_WIDTH - 1),
		19548 => to_unsigned(31271, LUT_AMPL_WIDTH - 1),
		19549 => to_unsigned(31270, LUT_AMPL_WIDTH - 1),
		19550 => to_unsigned(31269, LUT_AMPL_WIDTH - 1),
		19551 => to_unsigned(31268, LUT_AMPL_WIDTH - 1),
		19552 => to_unsigned(31267, LUT_AMPL_WIDTH - 1),
		19553 => to_unsigned(31266, LUT_AMPL_WIDTH - 1),
		19554 => to_unsigned(31265, LUT_AMPL_WIDTH - 1),
		19555 => to_unsigned(31264, LUT_AMPL_WIDTH - 1),
		19556 => to_unsigned(31263, LUT_AMPL_WIDTH - 1),
		19557 => to_unsigned(31262, LUT_AMPL_WIDTH - 1),
		19558 => to_unsigned(31262, LUT_AMPL_WIDTH - 1),
		19559 => to_unsigned(31261, LUT_AMPL_WIDTH - 1),
		19560 => to_unsigned(31260, LUT_AMPL_WIDTH - 1),
		19561 => to_unsigned(31259, LUT_AMPL_WIDTH - 1),
		19562 => to_unsigned(31258, LUT_AMPL_WIDTH - 1),
		19563 => to_unsigned(31257, LUT_AMPL_WIDTH - 1),
		19564 => to_unsigned(31256, LUT_AMPL_WIDTH - 1),
		19565 => to_unsigned(31255, LUT_AMPL_WIDTH - 1),
		19566 => to_unsigned(31254, LUT_AMPL_WIDTH - 1),
		19567 => to_unsigned(31253, LUT_AMPL_WIDTH - 1),
		19568 => to_unsigned(31252, LUT_AMPL_WIDTH - 1),
		19569 => to_unsigned(31251, LUT_AMPL_WIDTH - 1),
		19570 => to_unsigned(31250, LUT_AMPL_WIDTH - 1),
		19571 => to_unsigned(31249, LUT_AMPL_WIDTH - 1),
		19572 => to_unsigned(31248, LUT_AMPL_WIDTH - 1),
		19573 => to_unsigned(31247, LUT_AMPL_WIDTH - 1),
		19574 => to_unsigned(31246, LUT_AMPL_WIDTH - 1),
		19575 => to_unsigned(31246, LUT_AMPL_WIDTH - 1),
		19576 => to_unsigned(31245, LUT_AMPL_WIDTH - 1),
		19577 => to_unsigned(31244, LUT_AMPL_WIDTH - 1),
		19578 => to_unsigned(31243, LUT_AMPL_WIDTH - 1),
		19579 => to_unsigned(31242, LUT_AMPL_WIDTH - 1),
		19580 => to_unsigned(31241, LUT_AMPL_WIDTH - 1),
		19581 => to_unsigned(31240, LUT_AMPL_WIDTH - 1),
		19582 => to_unsigned(31239, LUT_AMPL_WIDTH - 1),
		19583 => to_unsigned(31238, LUT_AMPL_WIDTH - 1),
		19584 => to_unsigned(31237, LUT_AMPL_WIDTH - 1),
		19585 => to_unsigned(31236, LUT_AMPL_WIDTH - 1),
		19586 => to_unsigned(31235, LUT_AMPL_WIDTH - 1),
		19587 => to_unsigned(31234, LUT_AMPL_WIDTH - 1),
		19588 => to_unsigned(31233, LUT_AMPL_WIDTH - 1),
		19589 => to_unsigned(31232, LUT_AMPL_WIDTH - 1),
		19590 => to_unsigned(31231, LUT_AMPL_WIDTH - 1),
		19591 => to_unsigned(31230, LUT_AMPL_WIDTH - 1),
		19592 => to_unsigned(31229, LUT_AMPL_WIDTH - 1),
		19593 => to_unsigned(31228, LUT_AMPL_WIDTH - 1),
		19594 => to_unsigned(31227, LUT_AMPL_WIDTH - 1),
		19595 => to_unsigned(31227, LUT_AMPL_WIDTH - 1),
		19596 => to_unsigned(31226, LUT_AMPL_WIDTH - 1),
		19597 => to_unsigned(31225, LUT_AMPL_WIDTH - 1),
		19598 => to_unsigned(31224, LUT_AMPL_WIDTH - 1),
		19599 => to_unsigned(31223, LUT_AMPL_WIDTH - 1),
		19600 => to_unsigned(31222, LUT_AMPL_WIDTH - 1),
		19601 => to_unsigned(31221, LUT_AMPL_WIDTH - 1),
		19602 => to_unsigned(31220, LUT_AMPL_WIDTH - 1),
		19603 => to_unsigned(31219, LUT_AMPL_WIDTH - 1),
		19604 => to_unsigned(31218, LUT_AMPL_WIDTH - 1),
		19605 => to_unsigned(31217, LUT_AMPL_WIDTH - 1),
		19606 => to_unsigned(31216, LUT_AMPL_WIDTH - 1),
		19607 => to_unsigned(31215, LUT_AMPL_WIDTH - 1),
		19608 => to_unsigned(31214, LUT_AMPL_WIDTH - 1),
		19609 => to_unsigned(31213, LUT_AMPL_WIDTH - 1),
		19610 => to_unsigned(31212, LUT_AMPL_WIDTH - 1),
		19611 => to_unsigned(31211, LUT_AMPL_WIDTH - 1),
		19612 => to_unsigned(31210, LUT_AMPL_WIDTH - 1),
		19613 => to_unsigned(31209, LUT_AMPL_WIDTH - 1),
		19614 => to_unsigned(31208, LUT_AMPL_WIDTH - 1),
		19615 => to_unsigned(31207, LUT_AMPL_WIDTH - 1),
		19616 => to_unsigned(31206, LUT_AMPL_WIDTH - 1),
		19617 => to_unsigned(31206, LUT_AMPL_WIDTH - 1),
		19618 => to_unsigned(31205, LUT_AMPL_WIDTH - 1),
		19619 => to_unsigned(31204, LUT_AMPL_WIDTH - 1),
		19620 => to_unsigned(31203, LUT_AMPL_WIDTH - 1),
		19621 => to_unsigned(31202, LUT_AMPL_WIDTH - 1),
		19622 => to_unsigned(31201, LUT_AMPL_WIDTH - 1),
		19623 => to_unsigned(31200, LUT_AMPL_WIDTH - 1),
		19624 => to_unsigned(31199, LUT_AMPL_WIDTH - 1),
		19625 => to_unsigned(31198, LUT_AMPL_WIDTH - 1),
		19626 => to_unsigned(31197, LUT_AMPL_WIDTH - 1),
		19627 => to_unsigned(31196, LUT_AMPL_WIDTH - 1),
		19628 => to_unsigned(31195, LUT_AMPL_WIDTH - 1),
		19629 => to_unsigned(31194, LUT_AMPL_WIDTH - 1),
		19630 => to_unsigned(31193, LUT_AMPL_WIDTH - 1),
		19631 => to_unsigned(31192, LUT_AMPL_WIDTH - 1),
		19632 => to_unsigned(31191, LUT_AMPL_WIDTH - 1),
		19633 => to_unsigned(31190, LUT_AMPL_WIDTH - 1),
		19634 => to_unsigned(31189, LUT_AMPL_WIDTH - 1),
		19635 => to_unsigned(31188, LUT_AMPL_WIDTH - 1),
		19636 => to_unsigned(31187, LUT_AMPL_WIDTH - 1),
		19637 => to_unsigned(31186, LUT_AMPL_WIDTH - 1),
		19638 => to_unsigned(31185, LUT_AMPL_WIDTH - 1),
		19639 => to_unsigned(31184, LUT_AMPL_WIDTH - 1),
		19640 => to_unsigned(31183, LUT_AMPL_WIDTH - 1),
		19641 => to_unsigned(31182, LUT_AMPL_WIDTH - 1),
		19642 => to_unsigned(31181, LUT_AMPL_WIDTH - 1),
		19643 => to_unsigned(31181, LUT_AMPL_WIDTH - 1),
		19644 => to_unsigned(31180, LUT_AMPL_WIDTH - 1),
		19645 => to_unsigned(31179, LUT_AMPL_WIDTH - 1),
		19646 => to_unsigned(31178, LUT_AMPL_WIDTH - 1),
		19647 => to_unsigned(31177, LUT_AMPL_WIDTH - 1),
		19648 => to_unsigned(31176, LUT_AMPL_WIDTH - 1),
		19649 => to_unsigned(31175, LUT_AMPL_WIDTH - 1),
		19650 => to_unsigned(31174, LUT_AMPL_WIDTH - 1),
		19651 => to_unsigned(31173, LUT_AMPL_WIDTH - 1),
		19652 => to_unsigned(31172, LUT_AMPL_WIDTH - 1),
		19653 => to_unsigned(31171, LUT_AMPL_WIDTH - 1),
		19654 => to_unsigned(31170, LUT_AMPL_WIDTH - 1),
		19655 => to_unsigned(31169, LUT_AMPL_WIDTH - 1),
		19656 => to_unsigned(31168, LUT_AMPL_WIDTH - 1),
		19657 => to_unsigned(31167, LUT_AMPL_WIDTH - 1),
		19658 => to_unsigned(31166, LUT_AMPL_WIDTH - 1),
		19659 => to_unsigned(31165, LUT_AMPL_WIDTH - 1),
		19660 => to_unsigned(31164, LUT_AMPL_WIDTH - 1),
		19661 => to_unsigned(31163, LUT_AMPL_WIDTH - 1),
		19662 => to_unsigned(31162, LUT_AMPL_WIDTH - 1),
		19663 => to_unsigned(31161, LUT_AMPL_WIDTH - 1),
		19664 => to_unsigned(31160, LUT_AMPL_WIDTH - 1),
		19665 => to_unsigned(31159, LUT_AMPL_WIDTH - 1),
		19666 => to_unsigned(31158, LUT_AMPL_WIDTH - 1),
		19667 => to_unsigned(31157, LUT_AMPL_WIDTH - 1),
		19668 => to_unsigned(31156, LUT_AMPL_WIDTH - 1),
		19669 => to_unsigned(31155, LUT_AMPL_WIDTH - 1),
		19670 => to_unsigned(31154, LUT_AMPL_WIDTH - 1),
		19671 => to_unsigned(31153, LUT_AMPL_WIDTH - 1),
		19672 => to_unsigned(31152, LUT_AMPL_WIDTH - 1),
		19673 => to_unsigned(31151, LUT_AMPL_WIDTH - 1),
		19674 => to_unsigned(31150, LUT_AMPL_WIDTH - 1),
		19675 => to_unsigned(31149, LUT_AMPL_WIDTH - 1),
		19676 => to_unsigned(31148, LUT_AMPL_WIDTH - 1),
		19677 => to_unsigned(31148, LUT_AMPL_WIDTH - 1),
		19678 => to_unsigned(31147, LUT_AMPL_WIDTH - 1),
		19679 => to_unsigned(31146, LUT_AMPL_WIDTH - 1),
		19680 => to_unsigned(31145, LUT_AMPL_WIDTH - 1),
		19681 => to_unsigned(31144, LUT_AMPL_WIDTH - 1),
		19682 => to_unsigned(31143, LUT_AMPL_WIDTH - 1),
		19683 => to_unsigned(31142, LUT_AMPL_WIDTH - 1),
		19684 => to_unsigned(31141, LUT_AMPL_WIDTH - 1),
		19685 => to_unsigned(31140, LUT_AMPL_WIDTH - 1),
		19686 => to_unsigned(31139, LUT_AMPL_WIDTH - 1),
		19687 => to_unsigned(31138, LUT_AMPL_WIDTH - 1),
		19688 => to_unsigned(31137, LUT_AMPL_WIDTH - 1),
		19689 => to_unsigned(31136, LUT_AMPL_WIDTH - 1),
		19690 => to_unsigned(31135, LUT_AMPL_WIDTH - 1),
		19691 => to_unsigned(31134, LUT_AMPL_WIDTH - 1),
		19692 => to_unsigned(31133, LUT_AMPL_WIDTH - 1),
		19693 => to_unsigned(31132, LUT_AMPL_WIDTH - 1),
		19694 => to_unsigned(31131, LUT_AMPL_WIDTH - 1),
		19695 => to_unsigned(31130, LUT_AMPL_WIDTH - 1),
		19696 => to_unsigned(31129, LUT_AMPL_WIDTH - 1),
		19697 => to_unsigned(31128, LUT_AMPL_WIDTH - 1),
		19698 => to_unsigned(31127, LUT_AMPL_WIDTH - 1),
		19699 => to_unsigned(31126, LUT_AMPL_WIDTH - 1),
		19700 => to_unsigned(31125, LUT_AMPL_WIDTH - 1),
		19701 => to_unsigned(31124, LUT_AMPL_WIDTH - 1),
		19702 => to_unsigned(31123, LUT_AMPL_WIDTH - 1),
		19703 => to_unsigned(31122, LUT_AMPL_WIDTH - 1),
		19704 => to_unsigned(31121, LUT_AMPL_WIDTH - 1),
		19705 => to_unsigned(31120, LUT_AMPL_WIDTH - 1),
		19706 => to_unsigned(31119, LUT_AMPL_WIDTH - 1),
		19707 => to_unsigned(31118, LUT_AMPL_WIDTH - 1),
		19708 => to_unsigned(31117, LUT_AMPL_WIDTH - 1),
		19709 => to_unsigned(31116, LUT_AMPL_WIDTH - 1),
		19710 => to_unsigned(31115, LUT_AMPL_WIDTH - 1),
		19711 => to_unsigned(31114, LUT_AMPL_WIDTH - 1),
		19712 => to_unsigned(31113, LUT_AMPL_WIDTH - 1),
		19713 => to_unsigned(31112, LUT_AMPL_WIDTH - 1),
		19714 => to_unsigned(31111, LUT_AMPL_WIDTH - 1),
		19715 => to_unsigned(31110, LUT_AMPL_WIDTH - 1),
		19716 => to_unsigned(31109, LUT_AMPL_WIDTH - 1),
		19717 => to_unsigned(31108, LUT_AMPL_WIDTH - 1),
		19718 => to_unsigned(31107, LUT_AMPL_WIDTH - 1),
		19719 => to_unsigned(31106, LUT_AMPL_WIDTH - 1),
		19720 => to_unsigned(31105, LUT_AMPL_WIDTH - 1),
		19721 => to_unsigned(31104, LUT_AMPL_WIDTH - 1),
		19722 => to_unsigned(31103, LUT_AMPL_WIDTH - 1),
		19723 => to_unsigned(31102, LUT_AMPL_WIDTH - 1),
		19724 => to_unsigned(31101, LUT_AMPL_WIDTH - 1),
		19725 => to_unsigned(31100, LUT_AMPL_WIDTH - 1),
		19726 => to_unsigned(31099, LUT_AMPL_WIDTH - 1),
		19727 => to_unsigned(31098, LUT_AMPL_WIDTH - 1),
		19728 => to_unsigned(31097, LUT_AMPL_WIDTH - 1),
		19729 => to_unsigned(31096, LUT_AMPL_WIDTH - 1),
		19730 => to_unsigned(31095, LUT_AMPL_WIDTH - 1),
		19731 => to_unsigned(31094, LUT_AMPL_WIDTH - 1),
		19732 => to_unsigned(31093, LUT_AMPL_WIDTH - 1),
		19733 => to_unsigned(31092, LUT_AMPL_WIDTH - 1),
		19734 => to_unsigned(31091, LUT_AMPL_WIDTH - 1),
		19735 => to_unsigned(31090, LUT_AMPL_WIDTH - 1),
		19736 => to_unsigned(31089, LUT_AMPL_WIDTH - 1),
		19737 => to_unsigned(31088, LUT_AMPL_WIDTH - 1),
		19738 => to_unsigned(31087, LUT_AMPL_WIDTH - 1),
		19739 => to_unsigned(31086, LUT_AMPL_WIDTH - 1),
		19740 => to_unsigned(31085, LUT_AMPL_WIDTH - 1),
		19741 => to_unsigned(31084, LUT_AMPL_WIDTH - 1),
		19742 => to_unsigned(31083, LUT_AMPL_WIDTH - 1),
		19743 => to_unsigned(31083, LUT_AMPL_WIDTH - 1),
		19744 => to_unsigned(31082, LUT_AMPL_WIDTH - 1),
		19745 => to_unsigned(31081, LUT_AMPL_WIDTH - 1),
		19746 => to_unsigned(31080, LUT_AMPL_WIDTH - 1),
		19747 => to_unsigned(31079, LUT_AMPL_WIDTH - 1),
		19748 => to_unsigned(31078, LUT_AMPL_WIDTH - 1),
		19749 => to_unsigned(31077, LUT_AMPL_WIDTH - 1),
		19750 => to_unsigned(31076, LUT_AMPL_WIDTH - 1),
		19751 => to_unsigned(31075, LUT_AMPL_WIDTH - 1),
		19752 => to_unsigned(31074, LUT_AMPL_WIDTH - 1),
		19753 => to_unsigned(31073, LUT_AMPL_WIDTH - 1),
		19754 => to_unsigned(31072, LUT_AMPL_WIDTH - 1),
		19755 => to_unsigned(31071, LUT_AMPL_WIDTH - 1),
		19756 => to_unsigned(31070, LUT_AMPL_WIDTH - 1),
		19757 => to_unsigned(31069, LUT_AMPL_WIDTH - 1),
		19758 => to_unsigned(31068, LUT_AMPL_WIDTH - 1),
		19759 => to_unsigned(31067, LUT_AMPL_WIDTH - 1),
		19760 => to_unsigned(31066, LUT_AMPL_WIDTH - 1),
		19761 => to_unsigned(31065, LUT_AMPL_WIDTH - 1),
		19762 => to_unsigned(31064, LUT_AMPL_WIDTH - 1),
		19763 => to_unsigned(31063, LUT_AMPL_WIDTH - 1),
		19764 => to_unsigned(31062, LUT_AMPL_WIDTH - 1),
		19765 => to_unsigned(31061, LUT_AMPL_WIDTH - 1),
		19766 => to_unsigned(31060, LUT_AMPL_WIDTH - 1),
		19767 => to_unsigned(31059, LUT_AMPL_WIDTH - 1),
		19768 => to_unsigned(31058, LUT_AMPL_WIDTH - 1),
		19769 => to_unsigned(31057, LUT_AMPL_WIDTH - 1),
		19770 => to_unsigned(31056, LUT_AMPL_WIDTH - 1),
		19771 => to_unsigned(31055, LUT_AMPL_WIDTH - 1),
		19772 => to_unsigned(31054, LUT_AMPL_WIDTH - 1),
		19773 => to_unsigned(31053, LUT_AMPL_WIDTH - 1),
		19774 => to_unsigned(31052, LUT_AMPL_WIDTH - 1),
		19775 => to_unsigned(31051, LUT_AMPL_WIDTH - 1),
		19776 => to_unsigned(31050, LUT_AMPL_WIDTH - 1),
		19777 => to_unsigned(31049, LUT_AMPL_WIDTH - 1),
		19778 => to_unsigned(31048, LUT_AMPL_WIDTH - 1),
		19779 => to_unsigned(31047, LUT_AMPL_WIDTH - 1),
		19780 => to_unsigned(31046, LUT_AMPL_WIDTH - 1),
		19781 => to_unsigned(31045, LUT_AMPL_WIDTH - 1),
		19782 => to_unsigned(31044, LUT_AMPL_WIDTH - 1),
		19783 => to_unsigned(31043, LUT_AMPL_WIDTH - 1),
		19784 => to_unsigned(31041, LUT_AMPL_WIDTH - 1),
		19785 => to_unsigned(31040, LUT_AMPL_WIDTH - 1),
		19786 => to_unsigned(31039, LUT_AMPL_WIDTH - 1),
		19787 => to_unsigned(31038, LUT_AMPL_WIDTH - 1),
		19788 => to_unsigned(31037, LUT_AMPL_WIDTH - 1),
		19789 => to_unsigned(31036, LUT_AMPL_WIDTH - 1),
		19790 => to_unsigned(31035, LUT_AMPL_WIDTH - 1),
		19791 => to_unsigned(31034, LUT_AMPL_WIDTH - 1),
		19792 => to_unsigned(31033, LUT_AMPL_WIDTH - 1),
		19793 => to_unsigned(31032, LUT_AMPL_WIDTH - 1),
		19794 => to_unsigned(31031, LUT_AMPL_WIDTH - 1),
		19795 => to_unsigned(31030, LUT_AMPL_WIDTH - 1),
		19796 => to_unsigned(31029, LUT_AMPL_WIDTH - 1),
		19797 => to_unsigned(31028, LUT_AMPL_WIDTH - 1),
		19798 => to_unsigned(31027, LUT_AMPL_WIDTH - 1),
		19799 => to_unsigned(31026, LUT_AMPL_WIDTH - 1),
		19800 => to_unsigned(31025, LUT_AMPL_WIDTH - 1),
		19801 => to_unsigned(31024, LUT_AMPL_WIDTH - 1),
		19802 => to_unsigned(31023, LUT_AMPL_WIDTH - 1),
		19803 => to_unsigned(31022, LUT_AMPL_WIDTH - 1),
		19804 => to_unsigned(31021, LUT_AMPL_WIDTH - 1),
		19805 => to_unsigned(31020, LUT_AMPL_WIDTH - 1),
		19806 => to_unsigned(31019, LUT_AMPL_WIDTH - 1),
		19807 => to_unsigned(31018, LUT_AMPL_WIDTH - 1),
		19808 => to_unsigned(31017, LUT_AMPL_WIDTH - 1),
		19809 => to_unsigned(31016, LUT_AMPL_WIDTH - 1),
		19810 => to_unsigned(31015, LUT_AMPL_WIDTH - 1),
		19811 => to_unsigned(31014, LUT_AMPL_WIDTH - 1),
		19812 => to_unsigned(31013, LUT_AMPL_WIDTH - 1),
		19813 => to_unsigned(31012, LUT_AMPL_WIDTH - 1),
		19814 => to_unsigned(31011, LUT_AMPL_WIDTH - 1),
		19815 => to_unsigned(31010, LUT_AMPL_WIDTH - 1),
		19816 => to_unsigned(31009, LUT_AMPL_WIDTH - 1),
		19817 => to_unsigned(31008, LUT_AMPL_WIDTH - 1),
		19818 => to_unsigned(31007, LUT_AMPL_WIDTH - 1),
		19819 => to_unsigned(31006, LUT_AMPL_WIDTH - 1),
		19820 => to_unsigned(31005, LUT_AMPL_WIDTH - 1),
		19821 => to_unsigned(31004, LUT_AMPL_WIDTH - 1),
		19822 => to_unsigned(31003, LUT_AMPL_WIDTH - 1),
		19823 => to_unsigned(31002, LUT_AMPL_WIDTH - 1),
		19824 => to_unsigned(31001, LUT_AMPL_WIDTH - 1),
		19825 => to_unsigned(31000, LUT_AMPL_WIDTH - 1),
		19826 => to_unsigned(30999, LUT_AMPL_WIDTH - 1),
		19827 => to_unsigned(30998, LUT_AMPL_WIDTH - 1),
		19828 => to_unsigned(30997, LUT_AMPL_WIDTH - 1),
		19829 => to_unsigned(30996, LUT_AMPL_WIDTH - 1),
		19830 => to_unsigned(30995, LUT_AMPL_WIDTH - 1),
		19831 => to_unsigned(30994, LUT_AMPL_WIDTH - 1),
		19832 => to_unsigned(30993, LUT_AMPL_WIDTH - 1),
		19833 => to_unsigned(30992, LUT_AMPL_WIDTH - 1),
		19834 => to_unsigned(30991, LUT_AMPL_WIDTH - 1),
		19835 => to_unsigned(30990, LUT_AMPL_WIDTH - 1),
		19836 => to_unsigned(30989, LUT_AMPL_WIDTH - 1),
		19837 => to_unsigned(30988, LUT_AMPL_WIDTH - 1),
		19838 => to_unsigned(30987, LUT_AMPL_WIDTH - 1),
		19839 => to_unsigned(30986, LUT_AMPL_WIDTH - 1),
		19840 => to_unsigned(30985, LUT_AMPL_WIDTH - 1),
		19841 => to_unsigned(30984, LUT_AMPL_WIDTH - 1),
		19842 => to_unsigned(30983, LUT_AMPL_WIDTH - 1),
		19843 => to_unsigned(30982, LUT_AMPL_WIDTH - 1),
		19844 => to_unsigned(30981, LUT_AMPL_WIDTH - 1),
		19845 => to_unsigned(30980, LUT_AMPL_WIDTH - 1),
		19846 => to_unsigned(30979, LUT_AMPL_WIDTH - 1),
		19847 => to_unsigned(30978, LUT_AMPL_WIDTH - 1),
		19848 => to_unsigned(30977, LUT_AMPL_WIDTH - 1),
		19849 => to_unsigned(30976, LUT_AMPL_WIDTH - 1),
		19850 => to_unsigned(30974, LUT_AMPL_WIDTH - 1),
		19851 => to_unsigned(30973, LUT_AMPL_WIDTH - 1),
		19852 => to_unsigned(30972, LUT_AMPL_WIDTH - 1),
		19853 => to_unsigned(30971, LUT_AMPL_WIDTH - 1),
		19854 => to_unsigned(30970, LUT_AMPL_WIDTH - 1),
		19855 => to_unsigned(30969, LUT_AMPL_WIDTH - 1),
		19856 => to_unsigned(30968, LUT_AMPL_WIDTH - 1),
		19857 => to_unsigned(30967, LUT_AMPL_WIDTH - 1),
		19858 => to_unsigned(30966, LUT_AMPL_WIDTH - 1),
		19859 => to_unsigned(30965, LUT_AMPL_WIDTH - 1),
		19860 => to_unsigned(30964, LUT_AMPL_WIDTH - 1),
		19861 => to_unsigned(30963, LUT_AMPL_WIDTH - 1),
		19862 => to_unsigned(30962, LUT_AMPL_WIDTH - 1),
		19863 => to_unsigned(30961, LUT_AMPL_WIDTH - 1),
		19864 => to_unsigned(30960, LUT_AMPL_WIDTH - 1),
		19865 => to_unsigned(30959, LUT_AMPL_WIDTH - 1),
		19866 => to_unsigned(30958, LUT_AMPL_WIDTH - 1),
		19867 => to_unsigned(30957, LUT_AMPL_WIDTH - 1),
		19868 => to_unsigned(30956, LUT_AMPL_WIDTH - 1),
		19869 => to_unsigned(30955, LUT_AMPL_WIDTH - 1),
		19870 => to_unsigned(30954, LUT_AMPL_WIDTH - 1),
		19871 => to_unsigned(30953, LUT_AMPL_WIDTH - 1),
		19872 => to_unsigned(30952, LUT_AMPL_WIDTH - 1),
		19873 => to_unsigned(30951, LUT_AMPL_WIDTH - 1),
		19874 => to_unsigned(30950, LUT_AMPL_WIDTH - 1),
		19875 => to_unsigned(30949, LUT_AMPL_WIDTH - 1),
		19876 => to_unsigned(30948, LUT_AMPL_WIDTH - 1),
		19877 => to_unsigned(30947, LUT_AMPL_WIDTH - 1),
		19878 => to_unsigned(30946, LUT_AMPL_WIDTH - 1),
		19879 => to_unsigned(30945, LUT_AMPL_WIDTH - 1),
		19880 => to_unsigned(30944, LUT_AMPL_WIDTH - 1),
		19881 => to_unsigned(30943, LUT_AMPL_WIDTH - 1),
		19882 => to_unsigned(30942, LUT_AMPL_WIDTH - 1),
		19883 => to_unsigned(30941, LUT_AMPL_WIDTH - 1),
		19884 => to_unsigned(30939, LUT_AMPL_WIDTH - 1),
		19885 => to_unsigned(30938, LUT_AMPL_WIDTH - 1),
		19886 => to_unsigned(30937, LUT_AMPL_WIDTH - 1),
		19887 => to_unsigned(30936, LUT_AMPL_WIDTH - 1),
		19888 => to_unsigned(30935, LUT_AMPL_WIDTH - 1),
		19889 => to_unsigned(30934, LUT_AMPL_WIDTH - 1),
		19890 => to_unsigned(30933, LUT_AMPL_WIDTH - 1),
		19891 => to_unsigned(30932, LUT_AMPL_WIDTH - 1),
		19892 => to_unsigned(30931, LUT_AMPL_WIDTH - 1),
		19893 => to_unsigned(30930, LUT_AMPL_WIDTH - 1),
		19894 => to_unsigned(30929, LUT_AMPL_WIDTH - 1),
		19895 => to_unsigned(30928, LUT_AMPL_WIDTH - 1),
		19896 => to_unsigned(30927, LUT_AMPL_WIDTH - 1),
		19897 => to_unsigned(30926, LUT_AMPL_WIDTH - 1),
		19898 => to_unsigned(30925, LUT_AMPL_WIDTH - 1),
		19899 => to_unsigned(30924, LUT_AMPL_WIDTH - 1),
		19900 => to_unsigned(30923, LUT_AMPL_WIDTH - 1),
		19901 => to_unsigned(30922, LUT_AMPL_WIDTH - 1),
		19902 => to_unsigned(30921, LUT_AMPL_WIDTH - 1),
		19903 => to_unsigned(30920, LUT_AMPL_WIDTH - 1),
		19904 => to_unsigned(30919, LUT_AMPL_WIDTH - 1),
		19905 => to_unsigned(30918, LUT_AMPL_WIDTH - 1),
		19906 => to_unsigned(30917, LUT_AMPL_WIDTH - 1),
		19907 => to_unsigned(30916, LUT_AMPL_WIDTH - 1),
		19908 => to_unsigned(30915, LUT_AMPL_WIDTH - 1),
		19909 => to_unsigned(30914, LUT_AMPL_WIDTH - 1),
		19910 => to_unsigned(30912, LUT_AMPL_WIDTH - 1),
		19911 => to_unsigned(30911, LUT_AMPL_WIDTH - 1),
		19912 => to_unsigned(30910, LUT_AMPL_WIDTH - 1),
		19913 => to_unsigned(30909, LUT_AMPL_WIDTH - 1),
		19914 => to_unsigned(30908, LUT_AMPL_WIDTH - 1),
		19915 => to_unsigned(30907, LUT_AMPL_WIDTH - 1),
		19916 => to_unsigned(30906, LUT_AMPL_WIDTH - 1),
		19917 => to_unsigned(30905, LUT_AMPL_WIDTH - 1),
		19918 => to_unsigned(30904, LUT_AMPL_WIDTH - 1),
		19919 => to_unsigned(30903, LUT_AMPL_WIDTH - 1),
		19920 => to_unsigned(30902, LUT_AMPL_WIDTH - 1),
		19921 => to_unsigned(30901, LUT_AMPL_WIDTH - 1),
		19922 => to_unsigned(30900, LUT_AMPL_WIDTH - 1),
		19923 => to_unsigned(30899, LUT_AMPL_WIDTH - 1),
		19924 => to_unsigned(30898, LUT_AMPL_WIDTH - 1),
		19925 => to_unsigned(30897, LUT_AMPL_WIDTH - 1),
		19926 => to_unsigned(30896, LUT_AMPL_WIDTH - 1),
		19927 => to_unsigned(30895, LUT_AMPL_WIDTH - 1),
		19928 => to_unsigned(30894, LUT_AMPL_WIDTH - 1),
		19929 => to_unsigned(30893, LUT_AMPL_WIDTH - 1),
		19930 => to_unsigned(30892, LUT_AMPL_WIDTH - 1),
		19931 => to_unsigned(30891, LUT_AMPL_WIDTH - 1),
		19932 => to_unsigned(30889, LUT_AMPL_WIDTH - 1),
		19933 => to_unsigned(30888, LUT_AMPL_WIDTH - 1),
		19934 => to_unsigned(30887, LUT_AMPL_WIDTH - 1),
		19935 => to_unsigned(30886, LUT_AMPL_WIDTH - 1),
		19936 => to_unsigned(30885, LUT_AMPL_WIDTH - 1),
		19937 => to_unsigned(30884, LUT_AMPL_WIDTH - 1),
		19938 => to_unsigned(30883, LUT_AMPL_WIDTH - 1),
		19939 => to_unsigned(30882, LUT_AMPL_WIDTH - 1),
		19940 => to_unsigned(30881, LUT_AMPL_WIDTH - 1),
		19941 => to_unsigned(30880, LUT_AMPL_WIDTH - 1),
		19942 => to_unsigned(30879, LUT_AMPL_WIDTH - 1),
		19943 => to_unsigned(30878, LUT_AMPL_WIDTH - 1),
		19944 => to_unsigned(30877, LUT_AMPL_WIDTH - 1),
		19945 => to_unsigned(30876, LUT_AMPL_WIDTH - 1),
		19946 => to_unsigned(30875, LUT_AMPL_WIDTH - 1),
		19947 => to_unsigned(30874, LUT_AMPL_WIDTH - 1),
		19948 => to_unsigned(30873, LUT_AMPL_WIDTH - 1),
		19949 => to_unsigned(30872, LUT_AMPL_WIDTH - 1),
		19950 => to_unsigned(30871, LUT_AMPL_WIDTH - 1),
		19951 => to_unsigned(30870, LUT_AMPL_WIDTH - 1),
		19952 => to_unsigned(30868, LUT_AMPL_WIDTH - 1),
		19953 => to_unsigned(30867, LUT_AMPL_WIDTH - 1),
		19954 => to_unsigned(30866, LUT_AMPL_WIDTH - 1),
		19955 => to_unsigned(30865, LUT_AMPL_WIDTH - 1),
		19956 => to_unsigned(30864, LUT_AMPL_WIDTH - 1),
		19957 => to_unsigned(30863, LUT_AMPL_WIDTH - 1),
		19958 => to_unsigned(30862, LUT_AMPL_WIDTH - 1),
		19959 => to_unsigned(30861, LUT_AMPL_WIDTH - 1),
		19960 => to_unsigned(30860, LUT_AMPL_WIDTH - 1),
		19961 => to_unsigned(30859, LUT_AMPL_WIDTH - 1),
		19962 => to_unsigned(30858, LUT_AMPL_WIDTH - 1),
		19963 => to_unsigned(30857, LUT_AMPL_WIDTH - 1),
		19964 => to_unsigned(30856, LUT_AMPL_WIDTH - 1),
		19965 => to_unsigned(30855, LUT_AMPL_WIDTH - 1),
		19966 => to_unsigned(30854, LUT_AMPL_WIDTH - 1),
		19967 => to_unsigned(30853, LUT_AMPL_WIDTH - 1),
		19968 => to_unsigned(30852, LUT_AMPL_WIDTH - 1),
		19969 => to_unsigned(30851, LUT_AMPL_WIDTH - 1),
		19970 => to_unsigned(30849, LUT_AMPL_WIDTH - 1),
		19971 => to_unsigned(30848, LUT_AMPL_WIDTH - 1),
		19972 => to_unsigned(30847, LUT_AMPL_WIDTH - 1),
		19973 => to_unsigned(30846, LUT_AMPL_WIDTH - 1),
		19974 => to_unsigned(30845, LUT_AMPL_WIDTH - 1),
		19975 => to_unsigned(30844, LUT_AMPL_WIDTH - 1),
		19976 => to_unsigned(30843, LUT_AMPL_WIDTH - 1),
		19977 => to_unsigned(30842, LUT_AMPL_WIDTH - 1),
		19978 => to_unsigned(30841, LUT_AMPL_WIDTH - 1),
		19979 => to_unsigned(30840, LUT_AMPL_WIDTH - 1),
		19980 => to_unsigned(30839, LUT_AMPL_WIDTH - 1),
		19981 => to_unsigned(30838, LUT_AMPL_WIDTH - 1),
		19982 => to_unsigned(30837, LUT_AMPL_WIDTH - 1),
		19983 => to_unsigned(30836, LUT_AMPL_WIDTH - 1),
		19984 => to_unsigned(30835, LUT_AMPL_WIDTH - 1),
		19985 => to_unsigned(30834, LUT_AMPL_WIDTH - 1),
		19986 => to_unsigned(30832, LUT_AMPL_WIDTH - 1),
		19987 => to_unsigned(30831, LUT_AMPL_WIDTH - 1),
		19988 => to_unsigned(30830, LUT_AMPL_WIDTH - 1),
		19989 => to_unsigned(30829, LUT_AMPL_WIDTH - 1),
		19990 => to_unsigned(30828, LUT_AMPL_WIDTH - 1),
		19991 => to_unsigned(30827, LUT_AMPL_WIDTH - 1),
		19992 => to_unsigned(30826, LUT_AMPL_WIDTH - 1),
		19993 => to_unsigned(30825, LUT_AMPL_WIDTH - 1),
		19994 => to_unsigned(30824, LUT_AMPL_WIDTH - 1),
		19995 => to_unsigned(30823, LUT_AMPL_WIDTH - 1),
		19996 => to_unsigned(30822, LUT_AMPL_WIDTH - 1),
		19997 => to_unsigned(30821, LUT_AMPL_WIDTH - 1),
		19998 => to_unsigned(30820, LUT_AMPL_WIDTH - 1),
		19999 => to_unsigned(30819, LUT_AMPL_WIDTH - 1),
		20000 => to_unsigned(30818, LUT_AMPL_WIDTH - 1),
		20001 => to_unsigned(30816, LUT_AMPL_WIDTH - 1),
		20002 => to_unsigned(30815, LUT_AMPL_WIDTH - 1),
		20003 => to_unsigned(30814, LUT_AMPL_WIDTH - 1),
		20004 => to_unsigned(30813, LUT_AMPL_WIDTH - 1),
		20005 => to_unsigned(30812, LUT_AMPL_WIDTH - 1),
		20006 => to_unsigned(30811, LUT_AMPL_WIDTH - 1),
		20007 => to_unsigned(30810, LUT_AMPL_WIDTH - 1),
		20008 => to_unsigned(30809, LUT_AMPL_WIDTH - 1),
		20009 => to_unsigned(30808, LUT_AMPL_WIDTH - 1),
		20010 => to_unsigned(30807, LUT_AMPL_WIDTH - 1),
		20011 => to_unsigned(30806, LUT_AMPL_WIDTH - 1),
		20012 => to_unsigned(30805, LUT_AMPL_WIDTH - 1),
		20013 => to_unsigned(30804, LUT_AMPL_WIDTH - 1),
		20014 => to_unsigned(30803, LUT_AMPL_WIDTH - 1),
		20015 => to_unsigned(30802, LUT_AMPL_WIDTH - 1),
		20016 => to_unsigned(30800, LUT_AMPL_WIDTH - 1),
		20017 => to_unsigned(30799, LUT_AMPL_WIDTH - 1),
		20018 => to_unsigned(30798, LUT_AMPL_WIDTH - 1),
		20019 => to_unsigned(30797, LUT_AMPL_WIDTH - 1),
		20020 => to_unsigned(30796, LUT_AMPL_WIDTH - 1),
		20021 => to_unsigned(30795, LUT_AMPL_WIDTH - 1),
		20022 => to_unsigned(30794, LUT_AMPL_WIDTH - 1),
		20023 => to_unsigned(30793, LUT_AMPL_WIDTH - 1),
		20024 => to_unsigned(30792, LUT_AMPL_WIDTH - 1),
		20025 => to_unsigned(30791, LUT_AMPL_WIDTH - 1),
		20026 => to_unsigned(30790, LUT_AMPL_WIDTH - 1),
		20027 => to_unsigned(30789, LUT_AMPL_WIDTH - 1),
		20028 => to_unsigned(30788, LUT_AMPL_WIDTH - 1),
		20029 => to_unsigned(30786, LUT_AMPL_WIDTH - 1),
		20030 => to_unsigned(30785, LUT_AMPL_WIDTH - 1),
		20031 => to_unsigned(30784, LUT_AMPL_WIDTH - 1),
		20032 => to_unsigned(30783, LUT_AMPL_WIDTH - 1),
		20033 => to_unsigned(30782, LUT_AMPL_WIDTH - 1),
		20034 => to_unsigned(30781, LUT_AMPL_WIDTH - 1),
		20035 => to_unsigned(30780, LUT_AMPL_WIDTH - 1),
		20036 => to_unsigned(30779, LUT_AMPL_WIDTH - 1),
		20037 => to_unsigned(30778, LUT_AMPL_WIDTH - 1),
		20038 => to_unsigned(30777, LUT_AMPL_WIDTH - 1),
		20039 => to_unsigned(30776, LUT_AMPL_WIDTH - 1),
		20040 => to_unsigned(30775, LUT_AMPL_WIDTH - 1),
		20041 => to_unsigned(30774, LUT_AMPL_WIDTH - 1),
		20042 => to_unsigned(30772, LUT_AMPL_WIDTH - 1),
		20043 => to_unsigned(30771, LUT_AMPL_WIDTH - 1),
		20044 => to_unsigned(30770, LUT_AMPL_WIDTH - 1),
		20045 => to_unsigned(30769, LUT_AMPL_WIDTH - 1),
		20046 => to_unsigned(30768, LUT_AMPL_WIDTH - 1),
		20047 => to_unsigned(30767, LUT_AMPL_WIDTH - 1),
		20048 => to_unsigned(30766, LUT_AMPL_WIDTH - 1),
		20049 => to_unsigned(30765, LUT_AMPL_WIDTH - 1),
		20050 => to_unsigned(30764, LUT_AMPL_WIDTH - 1),
		20051 => to_unsigned(30763, LUT_AMPL_WIDTH - 1),
		20052 => to_unsigned(30762, LUT_AMPL_WIDTH - 1),
		20053 => to_unsigned(30761, LUT_AMPL_WIDTH - 1),
		20054 => to_unsigned(30760, LUT_AMPL_WIDTH - 1),
		20055 => to_unsigned(30758, LUT_AMPL_WIDTH - 1),
		20056 => to_unsigned(30757, LUT_AMPL_WIDTH - 1),
		20057 => to_unsigned(30756, LUT_AMPL_WIDTH - 1),
		20058 => to_unsigned(30755, LUT_AMPL_WIDTH - 1),
		20059 => to_unsigned(30754, LUT_AMPL_WIDTH - 1),
		20060 => to_unsigned(30753, LUT_AMPL_WIDTH - 1),
		20061 => to_unsigned(30752, LUT_AMPL_WIDTH - 1),
		20062 => to_unsigned(30751, LUT_AMPL_WIDTH - 1),
		20063 => to_unsigned(30750, LUT_AMPL_WIDTH - 1),
		20064 => to_unsigned(30749, LUT_AMPL_WIDTH - 1),
		20065 => to_unsigned(30748, LUT_AMPL_WIDTH - 1),
		20066 => to_unsigned(30746, LUT_AMPL_WIDTH - 1),
		20067 => to_unsigned(30745, LUT_AMPL_WIDTH - 1),
		20068 => to_unsigned(30744, LUT_AMPL_WIDTH - 1),
		20069 => to_unsigned(30743, LUT_AMPL_WIDTH - 1),
		20070 => to_unsigned(30742, LUT_AMPL_WIDTH - 1),
		20071 => to_unsigned(30741, LUT_AMPL_WIDTH - 1),
		20072 => to_unsigned(30740, LUT_AMPL_WIDTH - 1),
		20073 => to_unsigned(30739, LUT_AMPL_WIDTH - 1),
		20074 => to_unsigned(30738, LUT_AMPL_WIDTH - 1),
		20075 => to_unsigned(30737, LUT_AMPL_WIDTH - 1),
		20076 => to_unsigned(30736, LUT_AMPL_WIDTH - 1),
		20077 => to_unsigned(30735, LUT_AMPL_WIDTH - 1),
		20078 => to_unsigned(30733, LUT_AMPL_WIDTH - 1),
		20079 => to_unsigned(30732, LUT_AMPL_WIDTH - 1),
		20080 => to_unsigned(30731, LUT_AMPL_WIDTH - 1),
		20081 => to_unsigned(30730, LUT_AMPL_WIDTH - 1),
		20082 => to_unsigned(30729, LUT_AMPL_WIDTH - 1),
		20083 => to_unsigned(30728, LUT_AMPL_WIDTH - 1),
		20084 => to_unsigned(30727, LUT_AMPL_WIDTH - 1),
		20085 => to_unsigned(30726, LUT_AMPL_WIDTH - 1),
		20086 => to_unsigned(30725, LUT_AMPL_WIDTH - 1),
		20087 => to_unsigned(30724, LUT_AMPL_WIDTH - 1),
		20088 => to_unsigned(30723, LUT_AMPL_WIDTH - 1),
		20089 => to_unsigned(30721, LUT_AMPL_WIDTH - 1),
		20090 => to_unsigned(30720, LUT_AMPL_WIDTH - 1),
		20091 => to_unsigned(30719, LUT_AMPL_WIDTH - 1),
		20092 => to_unsigned(30718, LUT_AMPL_WIDTH - 1),
		20093 => to_unsigned(30717, LUT_AMPL_WIDTH - 1),
		20094 => to_unsigned(30716, LUT_AMPL_WIDTH - 1),
		20095 => to_unsigned(30715, LUT_AMPL_WIDTH - 1),
		20096 => to_unsigned(30714, LUT_AMPL_WIDTH - 1),
		20097 => to_unsigned(30713, LUT_AMPL_WIDTH - 1),
		20098 => to_unsigned(30712, LUT_AMPL_WIDTH - 1),
		20099 => to_unsigned(30711, LUT_AMPL_WIDTH - 1),
		20100 => to_unsigned(30709, LUT_AMPL_WIDTH - 1),
		20101 => to_unsigned(30708, LUT_AMPL_WIDTH - 1),
		20102 => to_unsigned(30707, LUT_AMPL_WIDTH - 1),
		20103 => to_unsigned(30706, LUT_AMPL_WIDTH - 1),
		20104 => to_unsigned(30705, LUT_AMPL_WIDTH - 1),
		20105 => to_unsigned(30704, LUT_AMPL_WIDTH - 1),
		20106 => to_unsigned(30703, LUT_AMPL_WIDTH - 1),
		20107 => to_unsigned(30702, LUT_AMPL_WIDTH - 1),
		20108 => to_unsigned(30701, LUT_AMPL_WIDTH - 1),
		20109 => to_unsigned(30700, LUT_AMPL_WIDTH - 1),
		20110 => to_unsigned(30698, LUT_AMPL_WIDTH - 1),
		20111 => to_unsigned(30697, LUT_AMPL_WIDTH - 1),
		20112 => to_unsigned(30696, LUT_AMPL_WIDTH - 1),
		20113 => to_unsigned(30695, LUT_AMPL_WIDTH - 1),
		20114 => to_unsigned(30694, LUT_AMPL_WIDTH - 1),
		20115 => to_unsigned(30693, LUT_AMPL_WIDTH - 1),
		20116 => to_unsigned(30692, LUT_AMPL_WIDTH - 1),
		20117 => to_unsigned(30691, LUT_AMPL_WIDTH - 1),
		20118 => to_unsigned(30690, LUT_AMPL_WIDTH - 1),
		20119 => to_unsigned(30689, LUT_AMPL_WIDTH - 1),
		20120 => to_unsigned(30687, LUT_AMPL_WIDTH - 1),
		20121 => to_unsigned(30686, LUT_AMPL_WIDTH - 1),
		20122 => to_unsigned(30685, LUT_AMPL_WIDTH - 1),
		20123 => to_unsigned(30684, LUT_AMPL_WIDTH - 1),
		20124 => to_unsigned(30683, LUT_AMPL_WIDTH - 1),
		20125 => to_unsigned(30682, LUT_AMPL_WIDTH - 1),
		20126 => to_unsigned(30681, LUT_AMPL_WIDTH - 1),
		20127 => to_unsigned(30680, LUT_AMPL_WIDTH - 1),
		20128 => to_unsigned(30679, LUT_AMPL_WIDTH - 1),
		20129 => to_unsigned(30678, LUT_AMPL_WIDTH - 1),
		20130 => to_unsigned(30676, LUT_AMPL_WIDTH - 1),
		20131 => to_unsigned(30675, LUT_AMPL_WIDTH - 1),
		20132 => to_unsigned(30674, LUT_AMPL_WIDTH - 1),
		20133 => to_unsigned(30673, LUT_AMPL_WIDTH - 1),
		20134 => to_unsigned(30672, LUT_AMPL_WIDTH - 1),
		20135 => to_unsigned(30671, LUT_AMPL_WIDTH - 1),
		20136 => to_unsigned(30670, LUT_AMPL_WIDTH - 1),
		20137 => to_unsigned(30669, LUT_AMPL_WIDTH - 1),
		20138 => to_unsigned(30668, LUT_AMPL_WIDTH - 1),
		20139 => to_unsigned(30666, LUT_AMPL_WIDTH - 1),
		20140 => to_unsigned(30665, LUT_AMPL_WIDTH - 1),
		20141 => to_unsigned(30664, LUT_AMPL_WIDTH - 1),
		20142 => to_unsigned(30663, LUT_AMPL_WIDTH - 1),
		20143 => to_unsigned(30662, LUT_AMPL_WIDTH - 1),
		20144 => to_unsigned(30661, LUT_AMPL_WIDTH - 1),
		20145 => to_unsigned(30660, LUT_AMPL_WIDTH - 1),
		20146 => to_unsigned(30659, LUT_AMPL_WIDTH - 1),
		20147 => to_unsigned(30658, LUT_AMPL_WIDTH - 1),
		20148 => to_unsigned(30656, LUT_AMPL_WIDTH - 1),
		20149 => to_unsigned(30655, LUT_AMPL_WIDTH - 1),
		20150 => to_unsigned(30654, LUT_AMPL_WIDTH - 1),
		20151 => to_unsigned(30653, LUT_AMPL_WIDTH - 1),
		20152 => to_unsigned(30652, LUT_AMPL_WIDTH - 1),
		20153 => to_unsigned(30651, LUT_AMPL_WIDTH - 1),
		20154 => to_unsigned(30650, LUT_AMPL_WIDTH - 1),
		20155 => to_unsigned(30649, LUT_AMPL_WIDTH - 1),
		20156 => to_unsigned(30648, LUT_AMPL_WIDTH - 1),
		20157 => to_unsigned(30646, LUT_AMPL_WIDTH - 1),
		20158 => to_unsigned(30645, LUT_AMPL_WIDTH - 1),
		20159 => to_unsigned(30644, LUT_AMPL_WIDTH - 1),
		20160 => to_unsigned(30643, LUT_AMPL_WIDTH - 1),
		20161 => to_unsigned(30642, LUT_AMPL_WIDTH - 1),
		20162 => to_unsigned(30641, LUT_AMPL_WIDTH - 1),
		20163 => to_unsigned(30640, LUT_AMPL_WIDTH - 1),
		20164 => to_unsigned(30639, LUT_AMPL_WIDTH - 1),
		20165 => to_unsigned(30638, LUT_AMPL_WIDTH - 1),
		20166 => to_unsigned(30636, LUT_AMPL_WIDTH - 1),
		20167 => to_unsigned(30635, LUT_AMPL_WIDTH - 1),
		20168 => to_unsigned(30634, LUT_AMPL_WIDTH - 1),
		20169 => to_unsigned(30633, LUT_AMPL_WIDTH - 1),
		20170 => to_unsigned(30632, LUT_AMPL_WIDTH - 1),
		20171 => to_unsigned(30631, LUT_AMPL_WIDTH - 1),
		20172 => to_unsigned(30630, LUT_AMPL_WIDTH - 1),
		20173 => to_unsigned(30629, LUT_AMPL_WIDTH - 1),
		20174 => to_unsigned(30628, LUT_AMPL_WIDTH - 1),
		20175 => to_unsigned(30626, LUT_AMPL_WIDTH - 1),
		20176 => to_unsigned(30625, LUT_AMPL_WIDTH - 1),
		20177 => to_unsigned(30624, LUT_AMPL_WIDTH - 1),
		20178 => to_unsigned(30623, LUT_AMPL_WIDTH - 1),
		20179 => to_unsigned(30622, LUT_AMPL_WIDTH - 1),
		20180 => to_unsigned(30621, LUT_AMPL_WIDTH - 1),
		20181 => to_unsigned(30620, LUT_AMPL_WIDTH - 1),
		20182 => to_unsigned(30619, LUT_AMPL_WIDTH - 1),
		20183 => to_unsigned(30617, LUT_AMPL_WIDTH - 1),
		20184 => to_unsigned(30616, LUT_AMPL_WIDTH - 1),
		20185 => to_unsigned(30615, LUT_AMPL_WIDTH - 1),
		20186 => to_unsigned(30614, LUT_AMPL_WIDTH - 1),
		20187 => to_unsigned(30613, LUT_AMPL_WIDTH - 1),
		20188 => to_unsigned(30612, LUT_AMPL_WIDTH - 1),
		20189 => to_unsigned(30611, LUT_AMPL_WIDTH - 1),
		20190 => to_unsigned(30610, LUT_AMPL_WIDTH - 1),
		20191 => to_unsigned(30609, LUT_AMPL_WIDTH - 1),
		20192 => to_unsigned(30607, LUT_AMPL_WIDTH - 1),
		20193 => to_unsigned(30606, LUT_AMPL_WIDTH - 1),
		20194 => to_unsigned(30605, LUT_AMPL_WIDTH - 1),
		20195 => to_unsigned(30604, LUT_AMPL_WIDTH - 1),
		20196 => to_unsigned(30603, LUT_AMPL_WIDTH - 1),
		20197 => to_unsigned(30602, LUT_AMPL_WIDTH - 1),
		20198 => to_unsigned(30601, LUT_AMPL_WIDTH - 1),
		20199 => to_unsigned(30600, LUT_AMPL_WIDTH - 1),
		20200 => to_unsigned(30598, LUT_AMPL_WIDTH - 1),
		20201 => to_unsigned(30597, LUT_AMPL_WIDTH - 1),
		20202 => to_unsigned(30596, LUT_AMPL_WIDTH - 1),
		20203 => to_unsigned(30595, LUT_AMPL_WIDTH - 1),
		20204 => to_unsigned(30594, LUT_AMPL_WIDTH - 1),
		20205 => to_unsigned(30593, LUT_AMPL_WIDTH - 1),
		20206 => to_unsigned(30592, LUT_AMPL_WIDTH - 1),
		20207 => to_unsigned(30591, LUT_AMPL_WIDTH - 1),
		20208 => to_unsigned(30589, LUT_AMPL_WIDTH - 1),
		20209 => to_unsigned(30588, LUT_AMPL_WIDTH - 1),
		20210 => to_unsigned(30587, LUT_AMPL_WIDTH - 1),
		20211 => to_unsigned(30586, LUT_AMPL_WIDTH - 1),
		20212 => to_unsigned(30585, LUT_AMPL_WIDTH - 1),
		20213 => to_unsigned(30584, LUT_AMPL_WIDTH - 1),
		20214 => to_unsigned(30583, LUT_AMPL_WIDTH - 1),
		20215 => to_unsigned(30582, LUT_AMPL_WIDTH - 1),
		20216 => to_unsigned(30580, LUT_AMPL_WIDTH - 1),
		20217 => to_unsigned(30579, LUT_AMPL_WIDTH - 1),
		20218 => to_unsigned(30578, LUT_AMPL_WIDTH - 1),
		20219 => to_unsigned(30577, LUT_AMPL_WIDTH - 1),
		20220 => to_unsigned(30576, LUT_AMPL_WIDTH - 1),
		20221 => to_unsigned(30575, LUT_AMPL_WIDTH - 1),
		20222 => to_unsigned(30574, LUT_AMPL_WIDTH - 1),
		20223 => to_unsigned(30573, LUT_AMPL_WIDTH - 1),
		20224 => to_unsigned(30571, LUT_AMPL_WIDTH - 1),
		20225 => to_unsigned(30570, LUT_AMPL_WIDTH - 1),
		20226 => to_unsigned(30569, LUT_AMPL_WIDTH - 1),
		20227 => to_unsigned(30568, LUT_AMPL_WIDTH - 1),
		20228 => to_unsigned(30567, LUT_AMPL_WIDTH - 1),
		20229 => to_unsigned(30566, LUT_AMPL_WIDTH - 1),
		20230 => to_unsigned(30565, LUT_AMPL_WIDTH - 1),
		20231 => to_unsigned(30563, LUT_AMPL_WIDTH - 1),
		20232 => to_unsigned(30562, LUT_AMPL_WIDTH - 1),
		20233 => to_unsigned(30561, LUT_AMPL_WIDTH - 1),
		20234 => to_unsigned(30560, LUT_AMPL_WIDTH - 1),
		20235 => to_unsigned(30559, LUT_AMPL_WIDTH - 1),
		20236 => to_unsigned(30558, LUT_AMPL_WIDTH - 1),
		20237 => to_unsigned(30557, LUT_AMPL_WIDTH - 1),
		20238 => to_unsigned(30556, LUT_AMPL_WIDTH - 1),
		20239 => to_unsigned(30554, LUT_AMPL_WIDTH - 1),
		20240 => to_unsigned(30553, LUT_AMPL_WIDTH - 1),
		20241 => to_unsigned(30552, LUT_AMPL_WIDTH - 1),
		20242 => to_unsigned(30551, LUT_AMPL_WIDTH - 1),
		20243 => to_unsigned(30550, LUT_AMPL_WIDTH - 1),
		20244 => to_unsigned(30549, LUT_AMPL_WIDTH - 1),
		20245 => to_unsigned(30548, LUT_AMPL_WIDTH - 1),
		20246 => to_unsigned(30546, LUT_AMPL_WIDTH - 1),
		20247 => to_unsigned(30545, LUT_AMPL_WIDTH - 1),
		20248 => to_unsigned(30544, LUT_AMPL_WIDTH - 1),
		20249 => to_unsigned(30543, LUT_AMPL_WIDTH - 1),
		20250 => to_unsigned(30542, LUT_AMPL_WIDTH - 1),
		20251 => to_unsigned(30541, LUT_AMPL_WIDTH - 1),
		20252 => to_unsigned(30540, LUT_AMPL_WIDTH - 1),
		20253 => to_unsigned(30538, LUT_AMPL_WIDTH - 1),
		20254 => to_unsigned(30537, LUT_AMPL_WIDTH - 1),
		20255 => to_unsigned(30536, LUT_AMPL_WIDTH - 1),
		20256 => to_unsigned(30535, LUT_AMPL_WIDTH - 1),
		20257 => to_unsigned(30534, LUT_AMPL_WIDTH - 1),
		20258 => to_unsigned(30533, LUT_AMPL_WIDTH - 1),
		20259 => to_unsigned(30532, LUT_AMPL_WIDTH - 1),
		20260 => to_unsigned(30530, LUT_AMPL_WIDTH - 1),
		20261 => to_unsigned(30529, LUT_AMPL_WIDTH - 1),
		20262 => to_unsigned(30528, LUT_AMPL_WIDTH - 1),
		20263 => to_unsigned(30527, LUT_AMPL_WIDTH - 1),
		20264 => to_unsigned(30526, LUT_AMPL_WIDTH - 1),
		20265 => to_unsigned(30525, LUT_AMPL_WIDTH - 1),
		20266 => to_unsigned(30524, LUT_AMPL_WIDTH - 1),
		20267 => to_unsigned(30522, LUT_AMPL_WIDTH - 1),
		20268 => to_unsigned(30521, LUT_AMPL_WIDTH - 1),
		20269 => to_unsigned(30520, LUT_AMPL_WIDTH - 1),
		20270 => to_unsigned(30519, LUT_AMPL_WIDTH - 1),
		20271 => to_unsigned(30518, LUT_AMPL_WIDTH - 1),
		20272 => to_unsigned(30517, LUT_AMPL_WIDTH - 1),
		20273 => to_unsigned(30516, LUT_AMPL_WIDTH - 1),
		20274 => to_unsigned(30514, LUT_AMPL_WIDTH - 1),
		20275 => to_unsigned(30513, LUT_AMPL_WIDTH - 1),
		20276 => to_unsigned(30512, LUT_AMPL_WIDTH - 1),
		20277 => to_unsigned(30511, LUT_AMPL_WIDTH - 1),
		20278 => to_unsigned(30510, LUT_AMPL_WIDTH - 1),
		20279 => to_unsigned(30509, LUT_AMPL_WIDTH - 1),
		20280 => to_unsigned(30508, LUT_AMPL_WIDTH - 1),
		20281 => to_unsigned(30506, LUT_AMPL_WIDTH - 1),
		20282 => to_unsigned(30505, LUT_AMPL_WIDTH - 1),
		20283 => to_unsigned(30504, LUT_AMPL_WIDTH - 1),
		20284 => to_unsigned(30503, LUT_AMPL_WIDTH - 1),
		20285 => to_unsigned(30502, LUT_AMPL_WIDTH - 1),
		20286 => to_unsigned(30501, LUT_AMPL_WIDTH - 1),
		20287 => to_unsigned(30500, LUT_AMPL_WIDTH - 1),
		20288 => to_unsigned(30498, LUT_AMPL_WIDTH - 1),
		20289 => to_unsigned(30497, LUT_AMPL_WIDTH - 1),
		20290 => to_unsigned(30496, LUT_AMPL_WIDTH - 1),
		20291 => to_unsigned(30495, LUT_AMPL_WIDTH - 1),
		20292 => to_unsigned(30494, LUT_AMPL_WIDTH - 1),
		20293 => to_unsigned(30493, LUT_AMPL_WIDTH - 1),
		20294 => to_unsigned(30492, LUT_AMPL_WIDTH - 1),
		20295 => to_unsigned(30490, LUT_AMPL_WIDTH - 1),
		20296 => to_unsigned(30489, LUT_AMPL_WIDTH - 1),
		20297 => to_unsigned(30488, LUT_AMPL_WIDTH - 1),
		20298 => to_unsigned(30487, LUT_AMPL_WIDTH - 1),
		20299 => to_unsigned(30486, LUT_AMPL_WIDTH - 1),
		20300 => to_unsigned(30485, LUT_AMPL_WIDTH - 1),
		20301 => to_unsigned(30483, LUT_AMPL_WIDTH - 1),
		20302 => to_unsigned(30482, LUT_AMPL_WIDTH - 1),
		20303 => to_unsigned(30481, LUT_AMPL_WIDTH - 1),
		20304 => to_unsigned(30480, LUT_AMPL_WIDTH - 1),
		20305 => to_unsigned(30479, LUT_AMPL_WIDTH - 1),
		20306 => to_unsigned(30478, LUT_AMPL_WIDTH - 1),
		20307 => to_unsigned(30477, LUT_AMPL_WIDTH - 1),
		20308 => to_unsigned(30475, LUT_AMPL_WIDTH - 1),
		20309 => to_unsigned(30474, LUT_AMPL_WIDTH - 1),
		20310 => to_unsigned(30473, LUT_AMPL_WIDTH - 1),
		20311 => to_unsigned(30472, LUT_AMPL_WIDTH - 1),
		20312 => to_unsigned(30471, LUT_AMPL_WIDTH - 1),
		20313 => to_unsigned(30470, LUT_AMPL_WIDTH - 1),
		20314 => to_unsigned(30468, LUT_AMPL_WIDTH - 1),
		20315 => to_unsigned(30467, LUT_AMPL_WIDTH - 1),
		20316 => to_unsigned(30466, LUT_AMPL_WIDTH - 1),
		20317 => to_unsigned(30465, LUT_AMPL_WIDTH - 1),
		20318 => to_unsigned(30464, LUT_AMPL_WIDTH - 1),
		20319 => to_unsigned(30463, LUT_AMPL_WIDTH - 1),
		20320 => to_unsigned(30462, LUT_AMPL_WIDTH - 1),
		20321 => to_unsigned(30460, LUT_AMPL_WIDTH - 1),
		20322 => to_unsigned(30459, LUT_AMPL_WIDTH - 1),
		20323 => to_unsigned(30458, LUT_AMPL_WIDTH - 1),
		20324 => to_unsigned(30457, LUT_AMPL_WIDTH - 1),
		20325 => to_unsigned(30456, LUT_AMPL_WIDTH - 1),
		20326 => to_unsigned(30455, LUT_AMPL_WIDTH - 1),
		20327 => to_unsigned(30453, LUT_AMPL_WIDTH - 1),
		20328 => to_unsigned(30452, LUT_AMPL_WIDTH - 1),
		20329 => to_unsigned(30451, LUT_AMPL_WIDTH - 1),
		20330 => to_unsigned(30450, LUT_AMPL_WIDTH - 1),
		20331 => to_unsigned(30449, LUT_AMPL_WIDTH - 1),
		20332 => to_unsigned(30448, LUT_AMPL_WIDTH - 1),
		20333 => to_unsigned(30446, LUT_AMPL_WIDTH - 1),
		20334 => to_unsigned(30445, LUT_AMPL_WIDTH - 1),
		20335 => to_unsigned(30444, LUT_AMPL_WIDTH - 1),
		20336 => to_unsigned(30443, LUT_AMPL_WIDTH - 1),
		20337 => to_unsigned(30442, LUT_AMPL_WIDTH - 1),
		20338 => to_unsigned(30441, LUT_AMPL_WIDTH - 1),
		20339 => to_unsigned(30439, LUT_AMPL_WIDTH - 1),
		20340 => to_unsigned(30438, LUT_AMPL_WIDTH - 1),
		20341 => to_unsigned(30437, LUT_AMPL_WIDTH - 1),
		20342 => to_unsigned(30436, LUT_AMPL_WIDTH - 1),
		20343 => to_unsigned(30435, LUT_AMPL_WIDTH - 1),
		20344 => to_unsigned(30434, LUT_AMPL_WIDTH - 1),
		20345 => to_unsigned(30433, LUT_AMPL_WIDTH - 1),
		20346 => to_unsigned(30431, LUT_AMPL_WIDTH - 1),
		20347 => to_unsigned(30430, LUT_AMPL_WIDTH - 1),
		20348 => to_unsigned(30429, LUT_AMPL_WIDTH - 1),
		20349 => to_unsigned(30428, LUT_AMPL_WIDTH - 1),
		20350 => to_unsigned(30427, LUT_AMPL_WIDTH - 1),
		20351 => to_unsigned(30426, LUT_AMPL_WIDTH - 1),
		20352 => to_unsigned(30424, LUT_AMPL_WIDTH - 1),
		20353 => to_unsigned(30423, LUT_AMPL_WIDTH - 1),
		20354 => to_unsigned(30422, LUT_AMPL_WIDTH - 1),
		20355 => to_unsigned(30421, LUT_AMPL_WIDTH - 1),
		20356 => to_unsigned(30420, LUT_AMPL_WIDTH - 1),
		20357 => to_unsigned(30419, LUT_AMPL_WIDTH - 1),
		20358 => to_unsigned(30417, LUT_AMPL_WIDTH - 1),
		20359 => to_unsigned(30416, LUT_AMPL_WIDTH - 1),
		20360 => to_unsigned(30415, LUT_AMPL_WIDTH - 1),
		20361 => to_unsigned(30414, LUT_AMPL_WIDTH - 1),
		20362 => to_unsigned(30413, LUT_AMPL_WIDTH - 1),
		20363 => to_unsigned(30412, LUT_AMPL_WIDTH - 1),
		20364 => to_unsigned(30410, LUT_AMPL_WIDTH - 1),
		20365 => to_unsigned(30409, LUT_AMPL_WIDTH - 1),
		20366 => to_unsigned(30408, LUT_AMPL_WIDTH - 1),
		20367 => to_unsigned(30407, LUT_AMPL_WIDTH - 1),
		20368 => to_unsigned(30406, LUT_AMPL_WIDTH - 1),
		20369 => to_unsigned(30404, LUT_AMPL_WIDTH - 1),
		20370 => to_unsigned(30403, LUT_AMPL_WIDTH - 1),
		20371 => to_unsigned(30402, LUT_AMPL_WIDTH - 1),
		20372 => to_unsigned(30401, LUT_AMPL_WIDTH - 1),
		20373 => to_unsigned(30400, LUT_AMPL_WIDTH - 1),
		20374 => to_unsigned(30399, LUT_AMPL_WIDTH - 1),
		20375 => to_unsigned(30397, LUT_AMPL_WIDTH - 1),
		20376 => to_unsigned(30396, LUT_AMPL_WIDTH - 1),
		20377 => to_unsigned(30395, LUT_AMPL_WIDTH - 1),
		20378 => to_unsigned(30394, LUT_AMPL_WIDTH - 1),
		20379 => to_unsigned(30393, LUT_AMPL_WIDTH - 1),
		20380 => to_unsigned(30392, LUT_AMPL_WIDTH - 1),
		20381 => to_unsigned(30390, LUT_AMPL_WIDTH - 1),
		20382 => to_unsigned(30389, LUT_AMPL_WIDTH - 1),
		20383 => to_unsigned(30388, LUT_AMPL_WIDTH - 1),
		20384 => to_unsigned(30387, LUT_AMPL_WIDTH - 1),
		20385 => to_unsigned(30386, LUT_AMPL_WIDTH - 1),
		20386 => to_unsigned(30385, LUT_AMPL_WIDTH - 1),
		20387 => to_unsigned(30383, LUT_AMPL_WIDTH - 1),
		20388 => to_unsigned(30382, LUT_AMPL_WIDTH - 1),
		20389 => to_unsigned(30381, LUT_AMPL_WIDTH - 1),
		20390 => to_unsigned(30380, LUT_AMPL_WIDTH - 1),
		20391 => to_unsigned(30379, LUT_AMPL_WIDTH - 1),
		20392 => to_unsigned(30377, LUT_AMPL_WIDTH - 1),
		20393 => to_unsigned(30376, LUT_AMPL_WIDTH - 1),
		20394 => to_unsigned(30375, LUT_AMPL_WIDTH - 1),
		20395 => to_unsigned(30374, LUT_AMPL_WIDTH - 1),
		20396 => to_unsigned(30373, LUT_AMPL_WIDTH - 1),
		20397 => to_unsigned(30372, LUT_AMPL_WIDTH - 1),
		20398 => to_unsigned(30370, LUT_AMPL_WIDTH - 1),
		20399 => to_unsigned(30369, LUT_AMPL_WIDTH - 1),
		20400 => to_unsigned(30368, LUT_AMPL_WIDTH - 1),
		20401 => to_unsigned(30367, LUT_AMPL_WIDTH - 1),
		20402 => to_unsigned(30366, LUT_AMPL_WIDTH - 1),
		20403 => to_unsigned(30365, LUT_AMPL_WIDTH - 1),
		20404 => to_unsigned(30363, LUT_AMPL_WIDTH - 1),
		20405 => to_unsigned(30362, LUT_AMPL_WIDTH - 1),
		20406 => to_unsigned(30361, LUT_AMPL_WIDTH - 1),
		20407 => to_unsigned(30360, LUT_AMPL_WIDTH - 1),
		20408 => to_unsigned(30359, LUT_AMPL_WIDTH - 1),
		20409 => to_unsigned(30357, LUT_AMPL_WIDTH - 1),
		20410 => to_unsigned(30356, LUT_AMPL_WIDTH - 1),
		20411 => to_unsigned(30355, LUT_AMPL_WIDTH - 1),
		20412 => to_unsigned(30354, LUT_AMPL_WIDTH - 1),
		20413 => to_unsigned(30353, LUT_AMPL_WIDTH - 1),
		20414 => to_unsigned(30351, LUT_AMPL_WIDTH - 1),
		20415 => to_unsigned(30350, LUT_AMPL_WIDTH - 1),
		20416 => to_unsigned(30349, LUT_AMPL_WIDTH - 1),
		20417 => to_unsigned(30348, LUT_AMPL_WIDTH - 1),
		20418 => to_unsigned(30347, LUT_AMPL_WIDTH - 1),
		20419 => to_unsigned(30346, LUT_AMPL_WIDTH - 1),
		20420 => to_unsigned(30344, LUT_AMPL_WIDTH - 1),
		20421 => to_unsigned(30343, LUT_AMPL_WIDTH - 1),
		20422 => to_unsigned(30342, LUT_AMPL_WIDTH - 1),
		20423 => to_unsigned(30341, LUT_AMPL_WIDTH - 1),
		20424 => to_unsigned(30340, LUT_AMPL_WIDTH - 1),
		20425 => to_unsigned(30338, LUT_AMPL_WIDTH - 1),
		20426 => to_unsigned(30337, LUT_AMPL_WIDTH - 1),
		20427 => to_unsigned(30336, LUT_AMPL_WIDTH - 1),
		20428 => to_unsigned(30335, LUT_AMPL_WIDTH - 1),
		20429 => to_unsigned(30334, LUT_AMPL_WIDTH - 1),
		20430 => to_unsigned(30333, LUT_AMPL_WIDTH - 1),
		20431 => to_unsigned(30331, LUT_AMPL_WIDTH - 1),
		20432 => to_unsigned(30330, LUT_AMPL_WIDTH - 1),
		20433 => to_unsigned(30329, LUT_AMPL_WIDTH - 1),
		20434 => to_unsigned(30328, LUT_AMPL_WIDTH - 1),
		20435 => to_unsigned(30327, LUT_AMPL_WIDTH - 1),
		20436 => to_unsigned(30325, LUT_AMPL_WIDTH - 1),
		20437 => to_unsigned(30324, LUT_AMPL_WIDTH - 1),
		20438 => to_unsigned(30323, LUT_AMPL_WIDTH - 1),
		20439 => to_unsigned(30322, LUT_AMPL_WIDTH - 1),
		20440 => to_unsigned(30321, LUT_AMPL_WIDTH - 1),
		20441 => to_unsigned(30319, LUT_AMPL_WIDTH - 1),
		20442 => to_unsigned(30318, LUT_AMPL_WIDTH - 1),
		20443 => to_unsigned(30317, LUT_AMPL_WIDTH - 1),
		20444 => to_unsigned(30316, LUT_AMPL_WIDTH - 1),
		20445 => to_unsigned(30315, LUT_AMPL_WIDTH - 1),
		20446 => to_unsigned(30313, LUT_AMPL_WIDTH - 1),
		20447 => to_unsigned(30312, LUT_AMPL_WIDTH - 1),
		20448 => to_unsigned(30311, LUT_AMPL_WIDTH - 1),
		20449 => to_unsigned(30310, LUT_AMPL_WIDTH - 1),
		20450 => to_unsigned(30309, LUT_AMPL_WIDTH - 1),
		20451 => to_unsigned(30308, LUT_AMPL_WIDTH - 1),
		20452 => to_unsigned(30306, LUT_AMPL_WIDTH - 1),
		20453 => to_unsigned(30305, LUT_AMPL_WIDTH - 1),
		20454 => to_unsigned(30304, LUT_AMPL_WIDTH - 1),
		20455 => to_unsigned(30303, LUT_AMPL_WIDTH - 1),
		20456 => to_unsigned(30302, LUT_AMPL_WIDTH - 1),
		20457 => to_unsigned(30300, LUT_AMPL_WIDTH - 1),
		20458 => to_unsigned(30299, LUT_AMPL_WIDTH - 1),
		20459 => to_unsigned(30298, LUT_AMPL_WIDTH - 1),
		20460 => to_unsigned(30297, LUT_AMPL_WIDTH - 1),
		20461 => to_unsigned(30296, LUT_AMPL_WIDTH - 1),
		20462 => to_unsigned(30294, LUT_AMPL_WIDTH - 1),
		20463 => to_unsigned(30293, LUT_AMPL_WIDTH - 1),
		20464 => to_unsigned(30292, LUT_AMPL_WIDTH - 1),
		20465 => to_unsigned(30291, LUT_AMPL_WIDTH - 1),
		20466 => to_unsigned(30290, LUT_AMPL_WIDTH - 1),
		20467 => to_unsigned(30288, LUT_AMPL_WIDTH - 1),
		20468 => to_unsigned(30287, LUT_AMPL_WIDTH - 1),
		20469 => to_unsigned(30286, LUT_AMPL_WIDTH - 1),
		20470 => to_unsigned(30285, LUT_AMPL_WIDTH - 1),
		20471 => to_unsigned(30284, LUT_AMPL_WIDTH - 1),
		20472 => to_unsigned(30282, LUT_AMPL_WIDTH - 1),
		20473 => to_unsigned(30281, LUT_AMPL_WIDTH - 1),
		20474 => to_unsigned(30280, LUT_AMPL_WIDTH - 1),
		20475 => to_unsigned(30279, LUT_AMPL_WIDTH - 1),
		20476 => to_unsigned(30278, LUT_AMPL_WIDTH - 1),
		20477 => to_unsigned(30276, LUT_AMPL_WIDTH - 1),
		20478 => to_unsigned(30275, LUT_AMPL_WIDTH - 1),
		20479 => to_unsigned(30274, LUT_AMPL_WIDTH - 1),
		20480 => to_unsigned(30273, LUT_AMPL_WIDTH - 1),
		20481 => to_unsigned(30272, LUT_AMPL_WIDTH - 1),
		20482 => to_unsigned(30270, LUT_AMPL_WIDTH - 1),
		20483 => to_unsigned(30269, LUT_AMPL_WIDTH - 1),
		20484 => to_unsigned(30268, LUT_AMPL_WIDTH - 1),
		20485 => to_unsigned(30267, LUT_AMPL_WIDTH - 1),
		20486 => to_unsigned(30266, LUT_AMPL_WIDTH - 1),
		20487 => to_unsigned(30264, LUT_AMPL_WIDTH - 1),
		20488 => to_unsigned(30263, LUT_AMPL_WIDTH - 1),
		20489 => to_unsigned(30262, LUT_AMPL_WIDTH - 1),
		20490 => to_unsigned(30261, LUT_AMPL_WIDTH - 1),
		20491 => to_unsigned(30260, LUT_AMPL_WIDTH - 1),
		20492 => to_unsigned(30258, LUT_AMPL_WIDTH - 1),
		20493 => to_unsigned(30257, LUT_AMPL_WIDTH - 1),
		20494 => to_unsigned(30256, LUT_AMPL_WIDTH - 1),
		20495 => to_unsigned(30255, LUT_AMPL_WIDTH - 1),
		20496 => to_unsigned(30253, LUT_AMPL_WIDTH - 1),
		20497 => to_unsigned(30252, LUT_AMPL_WIDTH - 1),
		20498 => to_unsigned(30251, LUT_AMPL_WIDTH - 1),
		20499 => to_unsigned(30250, LUT_AMPL_WIDTH - 1),
		20500 => to_unsigned(30249, LUT_AMPL_WIDTH - 1),
		20501 => to_unsigned(30247, LUT_AMPL_WIDTH - 1),
		20502 => to_unsigned(30246, LUT_AMPL_WIDTH - 1),
		20503 => to_unsigned(30245, LUT_AMPL_WIDTH - 1),
		20504 => to_unsigned(30244, LUT_AMPL_WIDTH - 1),
		20505 => to_unsigned(30243, LUT_AMPL_WIDTH - 1),
		20506 => to_unsigned(30241, LUT_AMPL_WIDTH - 1),
		20507 => to_unsigned(30240, LUT_AMPL_WIDTH - 1),
		20508 => to_unsigned(30239, LUT_AMPL_WIDTH - 1),
		20509 => to_unsigned(30238, LUT_AMPL_WIDTH - 1),
		20510 => to_unsigned(30237, LUT_AMPL_WIDTH - 1),
		20511 => to_unsigned(30235, LUT_AMPL_WIDTH - 1),
		20512 => to_unsigned(30234, LUT_AMPL_WIDTH - 1),
		20513 => to_unsigned(30233, LUT_AMPL_WIDTH - 1),
		20514 => to_unsigned(30232, LUT_AMPL_WIDTH - 1),
		20515 => to_unsigned(30231, LUT_AMPL_WIDTH - 1),
		20516 => to_unsigned(30229, LUT_AMPL_WIDTH - 1),
		20517 => to_unsigned(30228, LUT_AMPL_WIDTH - 1),
		20518 => to_unsigned(30227, LUT_AMPL_WIDTH - 1),
		20519 => to_unsigned(30226, LUT_AMPL_WIDTH - 1),
		20520 => to_unsigned(30224, LUT_AMPL_WIDTH - 1),
		20521 => to_unsigned(30223, LUT_AMPL_WIDTH - 1),
		20522 => to_unsigned(30222, LUT_AMPL_WIDTH - 1),
		20523 => to_unsigned(30221, LUT_AMPL_WIDTH - 1),
		20524 => to_unsigned(30220, LUT_AMPL_WIDTH - 1),
		20525 => to_unsigned(30218, LUT_AMPL_WIDTH - 1),
		20526 => to_unsigned(30217, LUT_AMPL_WIDTH - 1),
		20527 => to_unsigned(30216, LUT_AMPL_WIDTH - 1),
		20528 => to_unsigned(30215, LUT_AMPL_WIDTH - 1),
		20529 => to_unsigned(30214, LUT_AMPL_WIDTH - 1),
		20530 => to_unsigned(30212, LUT_AMPL_WIDTH - 1),
		20531 => to_unsigned(30211, LUT_AMPL_WIDTH - 1),
		20532 => to_unsigned(30210, LUT_AMPL_WIDTH - 1),
		20533 => to_unsigned(30209, LUT_AMPL_WIDTH - 1),
		20534 => to_unsigned(30207, LUT_AMPL_WIDTH - 1),
		20535 => to_unsigned(30206, LUT_AMPL_WIDTH - 1),
		20536 => to_unsigned(30205, LUT_AMPL_WIDTH - 1),
		20537 => to_unsigned(30204, LUT_AMPL_WIDTH - 1),
		20538 => to_unsigned(30203, LUT_AMPL_WIDTH - 1),
		20539 => to_unsigned(30201, LUT_AMPL_WIDTH - 1),
		20540 => to_unsigned(30200, LUT_AMPL_WIDTH - 1),
		20541 => to_unsigned(30199, LUT_AMPL_WIDTH - 1),
		20542 => to_unsigned(30198, LUT_AMPL_WIDTH - 1),
		20543 => to_unsigned(30196, LUT_AMPL_WIDTH - 1),
		20544 => to_unsigned(30195, LUT_AMPL_WIDTH - 1),
		20545 => to_unsigned(30194, LUT_AMPL_WIDTH - 1),
		20546 => to_unsigned(30193, LUT_AMPL_WIDTH - 1),
		20547 => to_unsigned(30192, LUT_AMPL_WIDTH - 1),
		20548 => to_unsigned(30190, LUT_AMPL_WIDTH - 1),
		20549 => to_unsigned(30189, LUT_AMPL_WIDTH - 1),
		20550 => to_unsigned(30188, LUT_AMPL_WIDTH - 1),
		20551 => to_unsigned(30187, LUT_AMPL_WIDTH - 1),
		20552 => to_unsigned(30185, LUT_AMPL_WIDTH - 1),
		20553 => to_unsigned(30184, LUT_AMPL_WIDTH - 1),
		20554 => to_unsigned(30183, LUT_AMPL_WIDTH - 1),
		20555 => to_unsigned(30182, LUT_AMPL_WIDTH - 1),
		20556 => to_unsigned(30181, LUT_AMPL_WIDTH - 1),
		20557 => to_unsigned(30179, LUT_AMPL_WIDTH - 1),
		20558 => to_unsigned(30178, LUT_AMPL_WIDTH - 1),
		20559 => to_unsigned(30177, LUT_AMPL_WIDTH - 1),
		20560 => to_unsigned(30176, LUT_AMPL_WIDTH - 1),
		20561 => to_unsigned(30174, LUT_AMPL_WIDTH - 1),
		20562 => to_unsigned(30173, LUT_AMPL_WIDTH - 1),
		20563 => to_unsigned(30172, LUT_AMPL_WIDTH - 1),
		20564 => to_unsigned(30171, LUT_AMPL_WIDTH - 1),
		20565 => to_unsigned(30170, LUT_AMPL_WIDTH - 1),
		20566 => to_unsigned(30168, LUT_AMPL_WIDTH - 1),
		20567 => to_unsigned(30167, LUT_AMPL_WIDTH - 1),
		20568 => to_unsigned(30166, LUT_AMPL_WIDTH - 1),
		20569 => to_unsigned(30165, LUT_AMPL_WIDTH - 1),
		20570 => to_unsigned(30163, LUT_AMPL_WIDTH - 1),
		20571 => to_unsigned(30162, LUT_AMPL_WIDTH - 1),
		20572 => to_unsigned(30161, LUT_AMPL_WIDTH - 1),
		20573 => to_unsigned(30160, LUT_AMPL_WIDTH - 1),
		20574 => to_unsigned(30159, LUT_AMPL_WIDTH - 1),
		20575 => to_unsigned(30157, LUT_AMPL_WIDTH - 1),
		20576 => to_unsigned(30156, LUT_AMPL_WIDTH - 1),
		20577 => to_unsigned(30155, LUT_AMPL_WIDTH - 1),
		20578 => to_unsigned(30154, LUT_AMPL_WIDTH - 1),
		20579 => to_unsigned(30152, LUT_AMPL_WIDTH - 1),
		20580 => to_unsigned(30151, LUT_AMPL_WIDTH - 1),
		20581 => to_unsigned(30150, LUT_AMPL_WIDTH - 1),
		20582 => to_unsigned(30149, LUT_AMPL_WIDTH - 1),
		20583 => to_unsigned(30147, LUT_AMPL_WIDTH - 1),
		20584 => to_unsigned(30146, LUT_AMPL_WIDTH - 1),
		20585 => to_unsigned(30145, LUT_AMPL_WIDTH - 1),
		20586 => to_unsigned(30144, LUT_AMPL_WIDTH - 1),
		20587 => to_unsigned(30143, LUT_AMPL_WIDTH - 1),
		20588 => to_unsigned(30141, LUT_AMPL_WIDTH - 1),
		20589 => to_unsigned(30140, LUT_AMPL_WIDTH - 1),
		20590 => to_unsigned(30139, LUT_AMPL_WIDTH - 1),
		20591 => to_unsigned(30138, LUT_AMPL_WIDTH - 1),
		20592 => to_unsigned(30136, LUT_AMPL_WIDTH - 1),
		20593 => to_unsigned(30135, LUT_AMPL_WIDTH - 1),
		20594 => to_unsigned(30134, LUT_AMPL_WIDTH - 1),
		20595 => to_unsigned(30133, LUT_AMPL_WIDTH - 1),
		20596 => to_unsigned(30131, LUT_AMPL_WIDTH - 1),
		20597 => to_unsigned(30130, LUT_AMPL_WIDTH - 1),
		20598 => to_unsigned(30129, LUT_AMPL_WIDTH - 1),
		20599 => to_unsigned(30128, LUT_AMPL_WIDTH - 1),
		20600 => to_unsigned(30126, LUT_AMPL_WIDTH - 1),
		20601 => to_unsigned(30125, LUT_AMPL_WIDTH - 1),
		20602 => to_unsigned(30124, LUT_AMPL_WIDTH - 1),
		20603 => to_unsigned(30123, LUT_AMPL_WIDTH - 1),
		20604 => to_unsigned(30122, LUT_AMPL_WIDTH - 1),
		20605 => to_unsigned(30120, LUT_AMPL_WIDTH - 1),
		20606 => to_unsigned(30119, LUT_AMPL_WIDTH - 1),
		20607 => to_unsigned(30118, LUT_AMPL_WIDTH - 1),
		20608 => to_unsigned(30117, LUT_AMPL_WIDTH - 1),
		20609 => to_unsigned(30115, LUT_AMPL_WIDTH - 1),
		20610 => to_unsigned(30114, LUT_AMPL_WIDTH - 1),
		20611 => to_unsigned(30113, LUT_AMPL_WIDTH - 1),
		20612 => to_unsigned(30112, LUT_AMPL_WIDTH - 1),
		20613 => to_unsigned(30110, LUT_AMPL_WIDTH - 1),
		20614 => to_unsigned(30109, LUT_AMPL_WIDTH - 1),
		20615 => to_unsigned(30108, LUT_AMPL_WIDTH - 1),
		20616 => to_unsigned(30107, LUT_AMPL_WIDTH - 1),
		20617 => to_unsigned(30105, LUT_AMPL_WIDTH - 1),
		20618 => to_unsigned(30104, LUT_AMPL_WIDTH - 1),
		20619 => to_unsigned(30103, LUT_AMPL_WIDTH - 1),
		20620 => to_unsigned(30102, LUT_AMPL_WIDTH - 1),
		20621 => to_unsigned(30100, LUT_AMPL_WIDTH - 1),
		20622 => to_unsigned(30099, LUT_AMPL_WIDTH - 1),
		20623 => to_unsigned(30098, LUT_AMPL_WIDTH - 1),
		20624 => to_unsigned(30097, LUT_AMPL_WIDTH - 1),
		20625 => to_unsigned(30096, LUT_AMPL_WIDTH - 1),
		20626 => to_unsigned(30094, LUT_AMPL_WIDTH - 1),
		20627 => to_unsigned(30093, LUT_AMPL_WIDTH - 1),
		20628 => to_unsigned(30092, LUT_AMPL_WIDTH - 1),
		20629 => to_unsigned(30091, LUT_AMPL_WIDTH - 1),
		20630 => to_unsigned(30089, LUT_AMPL_WIDTH - 1),
		20631 => to_unsigned(30088, LUT_AMPL_WIDTH - 1),
		20632 => to_unsigned(30087, LUT_AMPL_WIDTH - 1),
		20633 => to_unsigned(30086, LUT_AMPL_WIDTH - 1),
		20634 => to_unsigned(30084, LUT_AMPL_WIDTH - 1),
		20635 => to_unsigned(30083, LUT_AMPL_WIDTH - 1),
		20636 => to_unsigned(30082, LUT_AMPL_WIDTH - 1),
		20637 => to_unsigned(30081, LUT_AMPL_WIDTH - 1),
		20638 => to_unsigned(30079, LUT_AMPL_WIDTH - 1),
		20639 => to_unsigned(30078, LUT_AMPL_WIDTH - 1),
		20640 => to_unsigned(30077, LUT_AMPL_WIDTH - 1),
		20641 => to_unsigned(30076, LUT_AMPL_WIDTH - 1),
		20642 => to_unsigned(30074, LUT_AMPL_WIDTH - 1),
		20643 => to_unsigned(30073, LUT_AMPL_WIDTH - 1),
		20644 => to_unsigned(30072, LUT_AMPL_WIDTH - 1),
		20645 => to_unsigned(30071, LUT_AMPL_WIDTH - 1),
		20646 => to_unsigned(30069, LUT_AMPL_WIDTH - 1),
		20647 => to_unsigned(30068, LUT_AMPL_WIDTH - 1),
		20648 => to_unsigned(30067, LUT_AMPL_WIDTH - 1),
		20649 => to_unsigned(30066, LUT_AMPL_WIDTH - 1),
		20650 => to_unsigned(30064, LUT_AMPL_WIDTH - 1),
		20651 => to_unsigned(30063, LUT_AMPL_WIDTH - 1),
		20652 => to_unsigned(30062, LUT_AMPL_WIDTH - 1),
		20653 => to_unsigned(30061, LUT_AMPL_WIDTH - 1),
		20654 => to_unsigned(30059, LUT_AMPL_WIDTH - 1),
		20655 => to_unsigned(30058, LUT_AMPL_WIDTH - 1),
		20656 => to_unsigned(30057, LUT_AMPL_WIDTH - 1),
		20657 => to_unsigned(30056, LUT_AMPL_WIDTH - 1),
		20658 => to_unsigned(30054, LUT_AMPL_WIDTH - 1),
		20659 => to_unsigned(30053, LUT_AMPL_WIDTH - 1),
		20660 => to_unsigned(30052, LUT_AMPL_WIDTH - 1),
		20661 => to_unsigned(30051, LUT_AMPL_WIDTH - 1),
		20662 => to_unsigned(30049, LUT_AMPL_WIDTH - 1),
		20663 => to_unsigned(30048, LUT_AMPL_WIDTH - 1),
		20664 => to_unsigned(30047, LUT_AMPL_WIDTH - 1),
		20665 => to_unsigned(30046, LUT_AMPL_WIDTH - 1),
		20666 => to_unsigned(30044, LUT_AMPL_WIDTH - 1),
		20667 => to_unsigned(30043, LUT_AMPL_WIDTH - 1),
		20668 => to_unsigned(30042, LUT_AMPL_WIDTH - 1),
		20669 => to_unsigned(30041, LUT_AMPL_WIDTH - 1),
		20670 => to_unsigned(30039, LUT_AMPL_WIDTH - 1),
		20671 => to_unsigned(30038, LUT_AMPL_WIDTH - 1),
		20672 => to_unsigned(30037, LUT_AMPL_WIDTH - 1),
		20673 => to_unsigned(30036, LUT_AMPL_WIDTH - 1),
		20674 => to_unsigned(30034, LUT_AMPL_WIDTH - 1),
		20675 => to_unsigned(30033, LUT_AMPL_WIDTH - 1),
		20676 => to_unsigned(30032, LUT_AMPL_WIDTH - 1),
		20677 => to_unsigned(30031, LUT_AMPL_WIDTH - 1),
		20678 => to_unsigned(30029, LUT_AMPL_WIDTH - 1),
		20679 => to_unsigned(30028, LUT_AMPL_WIDTH - 1),
		20680 => to_unsigned(30027, LUT_AMPL_WIDTH - 1),
		20681 => to_unsigned(30026, LUT_AMPL_WIDTH - 1),
		20682 => to_unsigned(30024, LUT_AMPL_WIDTH - 1),
		20683 => to_unsigned(30023, LUT_AMPL_WIDTH - 1),
		20684 => to_unsigned(30022, LUT_AMPL_WIDTH - 1),
		20685 => to_unsigned(30020, LUT_AMPL_WIDTH - 1),
		20686 => to_unsigned(30019, LUT_AMPL_WIDTH - 1),
		20687 => to_unsigned(30018, LUT_AMPL_WIDTH - 1),
		20688 => to_unsigned(30017, LUT_AMPL_WIDTH - 1),
		20689 => to_unsigned(30015, LUT_AMPL_WIDTH - 1),
		20690 => to_unsigned(30014, LUT_AMPL_WIDTH - 1),
		20691 => to_unsigned(30013, LUT_AMPL_WIDTH - 1),
		20692 => to_unsigned(30012, LUT_AMPL_WIDTH - 1),
		20693 => to_unsigned(30010, LUT_AMPL_WIDTH - 1),
		20694 => to_unsigned(30009, LUT_AMPL_WIDTH - 1),
		20695 => to_unsigned(30008, LUT_AMPL_WIDTH - 1),
		20696 => to_unsigned(30007, LUT_AMPL_WIDTH - 1),
		20697 => to_unsigned(30005, LUT_AMPL_WIDTH - 1),
		20698 => to_unsigned(30004, LUT_AMPL_WIDTH - 1),
		20699 => to_unsigned(30003, LUT_AMPL_WIDTH - 1),
		20700 => to_unsigned(30002, LUT_AMPL_WIDTH - 1),
		20701 => to_unsigned(30000, LUT_AMPL_WIDTH - 1),
		20702 => to_unsigned(29999, LUT_AMPL_WIDTH - 1),
		20703 => to_unsigned(29998, LUT_AMPL_WIDTH - 1),
		20704 => to_unsigned(29997, LUT_AMPL_WIDTH - 1),
		20705 => to_unsigned(29995, LUT_AMPL_WIDTH - 1),
		20706 => to_unsigned(29994, LUT_AMPL_WIDTH - 1),
		20707 => to_unsigned(29993, LUT_AMPL_WIDTH - 1),
		20708 => to_unsigned(29991, LUT_AMPL_WIDTH - 1),
		20709 => to_unsigned(29990, LUT_AMPL_WIDTH - 1),
		20710 => to_unsigned(29989, LUT_AMPL_WIDTH - 1),
		20711 => to_unsigned(29988, LUT_AMPL_WIDTH - 1),
		20712 => to_unsigned(29986, LUT_AMPL_WIDTH - 1),
		20713 => to_unsigned(29985, LUT_AMPL_WIDTH - 1),
		20714 => to_unsigned(29984, LUT_AMPL_WIDTH - 1),
		20715 => to_unsigned(29983, LUT_AMPL_WIDTH - 1),
		20716 => to_unsigned(29981, LUT_AMPL_WIDTH - 1),
		20717 => to_unsigned(29980, LUT_AMPL_WIDTH - 1),
		20718 => to_unsigned(29979, LUT_AMPL_WIDTH - 1),
		20719 => to_unsigned(29978, LUT_AMPL_WIDTH - 1),
		20720 => to_unsigned(29976, LUT_AMPL_WIDTH - 1),
		20721 => to_unsigned(29975, LUT_AMPL_WIDTH - 1),
		20722 => to_unsigned(29974, LUT_AMPL_WIDTH - 1),
		20723 => to_unsigned(29972, LUT_AMPL_WIDTH - 1),
		20724 => to_unsigned(29971, LUT_AMPL_WIDTH - 1),
		20725 => to_unsigned(29970, LUT_AMPL_WIDTH - 1),
		20726 => to_unsigned(29969, LUT_AMPL_WIDTH - 1),
		20727 => to_unsigned(29967, LUT_AMPL_WIDTH - 1),
		20728 => to_unsigned(29966, LUT_AMPL_WIDTH - 1),
		20729 => to_unsigned(29965, LUT_AMPL_WIDTH - 1),
		20730 => to_unsigned(29964, LUT_AMPL_WIDTH - 1),
		20731 => to_unsigned(29962, LUT_AMPL_WIDTH - 1),
		20732 => to_unsigned(29961, LUT_AMPL_WIDTH - 1),
		20733 => to_unsigned(29960, LUT_AMPL_WIDTH - 1),
		20734 => to_unsigned(29958, LUT_AMPL_WIDTH - 1),
		20735 => to_unsigned(29957, LUT_AMPL_WIDTH - 1),
		20736 => to_unsigned(29956, LUT_AMPL_WIDTH - 1),
		20737 => to_unsigned(29955, LUT_AMPL_WIDTH - 1),
		20738 => to_unsigned(29953, LUT_AMPL_WIDTH - 1),
		20739 => to_unsigned(29952, LUT_AMPL_WIDTH - 1),
		20740 => to_unsigned(29951, LUT_AMPL_WIDTH - 1),
		20741 => to_unsigned(29950, LUT_AMPL_WIDTH - 1),
		20742 => to_unsigned(29948, LUT_AMPL_WIDTH - 1),
		20743 => to_unsigned(29947, LUT_AMPL_WIDTH - 1),
		20744 => to_unsigned(29946, LUT_AMPL_WIDTH - 1),
		20745 => to_unsigned(29944, LUT_AMPL_WIDTH - 1),
		20746 => to_unsigned(29943, LUT_AMPL_WIDTH - 1),
		20747 => to_unsigned(29942, LUT_AMPL_WIDTH - 1),
		20748 => to_unsigned(29941, LUT_AMPL_WIDTH - 1),
		20749 => to_unsigned(29939, LUT_AMPL_WIDTH - 1),
		20750 => to_unsigned(29938, LUT_AMPL_WIDTH - 1),
		20751 => to_unsigned(29937, LUT_AMPL_WIDTH - 1),
		20752 => to_unsigned(29936, LUT_AMPL_WIDTH - 1),
		20753 => to_unsigned(29934, LUT_AMPL_WIDTH - 1),
		20754 => to_unsigned(29933, LUT_AMPL_WIDTH - 1),
		20755 => to_unsigned(29932, LUT_AMPL_WIDTH - 1),
		20756 => to_unsigned(29930, LUT_AMPL_WIDTH - 1),
		20757 => to_unsigned(29929, LUT_AMPL_WIDTH - 1),
		20758 => to_unsigned(29928, LUT_AMPL_WIDTH - 1),
		20759 => to_unsigned(29927, LUT_AMPL_WIDTH - 1),
		20760 => to_unsigned(29925, LUT_AMPL_WIDTH - 1),
		20761 => to_unsigned(29924, LUT_AMPL_WIDTH - 1),
		20762 => to_unsigned(29923, LUT_AMPL_WIDTH - 1),
		20763 => to_unsigned(29921, LUT_AMPL_WIDTH - 1),
		20764 => to_unsigned(29920, LUT_AMPL_WIDTH - 1),
		20765 => to_unsigned(29919, LUT_AMPL_WIDTH - 1),
		20766 => to_unsigned(29918, LUT_AMPL_WIDTH - 1),
		20767 => to_unsigned(29916, LUT_AMPL_WIDTH - 1),
		20768 => to_unsigned(29915, LUT_AMPL_WIDTH - 1),
		20769 => to_unsigned(29914, LUT_AMPL_WIDTH - 1),
		20770 => to_unsigned(29912, LUT_AMPL_WIDTH - 1),
		20771 => to_unsigned(29911, LUT_AMPL_WIDTH - 1),
		20772 => to_unsigned(29910, LUT_AMPL_WIDTH - 1),
		20773 => to_unsigned(29909, LUT_AMPL_WIDTH - 1),
		20774 => to_unsigned(29907, LUT_AMPL_WIDTH - 1),
		20775 => to_unsigned(29906, LUT_AMPL_WIDTH - 1),
		20776 => to_unsigned(29905, LUT_AMPL_WIDTH - 1),
		20777 => to_unsigned(29903, LUT_AMPL_WIDTH - 1),
		20778 => to_unsigned(29902, LUT_AMPL_WIDTH - 1),
		20779 => to_unsigned(29901, LUT_AMPL_WIDTH - 1),
		20780 => to_unsigned(29900, LUT_AMPL_WIDTH - 1),
		20781 => to_unsigned(29898, LUT_AMPL_WIDTH - 1),
		20782 => to_unsigned(29897, LUT_AMPL_WIDTH - 1),
		20783 => to_unsigned(29896, LUT_AMPL_WIDTH - 1),
		20784 => to_unsigned(29894, LUT_AMPL_WIDTH - 1),
		20785 => to_unsigned(29893, LUT_AMPL_WIDTH - 1),
		20786 => to_unsigned(29892, LUT_AMPL_WIDTH - 1),
		20787 => to_unsigned(29891, LUT_AMPL_WIDTH - 1),
		20788 => to_unsigned(29889, LUT_AMPL_WIDTH - 1),
		20789 => to_unsigned(29888, LUT_AMPL_WIDTH - 1),
		20790 => to_unsigned(29887, LUT_AMPL_WIDTH - 1),
		20791 => to_unsigned(29885, LUT_AMPL_WIDTH - 1),
		20792 => to_unsigned(29884, LUT_AMPL_WIDTH - 1),
		20793 => to_unsigned(29883, LUT_AMPL_WIDTH - 1),
		20794 => to_unsigned(29882, LUT_AMPL_WIDTH - 1),
		20795 => to_unsigned(29880, LUT_AMPL_WIDTH - 1),
		20796 => to_unsigned(29879, LUT_AMPL_WIDTH - 1),
		20797 => to_unsigned(29878, LUT_AMPL_WIDTH - 1),
		20798 => to_unsigned(29876, LUT_AMPL_WIDTH - 1),
		20799 => to_unsigned(29875, LUT_AMPL_WIDTH - 1),
		20800 => to_unsigned(29874, LUT_AMPL_WIDTH - 1),
		20801 => to_unsigned(29873, LUT_AMPL_WIDTH - 1),
		20802 => to_unsigned(29871, LUT_AMPL_WIDTH - 1),
		20803 => to_unsigned(29870, LUT_AMPL_WIDTH - 1),
		20804 => to_unsigned(29869, LUT_AMPL_WIDTH - 1),
		20805 => to_unsigned(29867, LUT_AMPL_WIDTH - 1),
		20806 => to_unsigned(29866, LUT_AMPL_WIDTH - 1),
		20807 => to_unsigned(29865, LUT_AMPL_WIDTH - 1),
		20808 => to_unsigned(29864, LUT_AMPL_WIDTH - 1),
		20809 => to_unsigned(29862, LUT_AMPL_WIDTH - 1),
		20810 => to_unsigned(29861, LUT_AMPL_WIDTH - 1),
		20811 => to_unsigned(29860, LUT_AMPL_WIDTH - 1),
		20812 => to_unsigned(29858, LUT_AMPL_WIDTH - 1),
		20813 => to_unsigned(29857, LUT_AMPL_WIDTH - 1),
		20814 => to_unsigned(29856, LUT_AMPL_WIDTH - 1),
		20815 => to_unsigned(29854, LUT_AMPL_WIDTH - 1),
		20816 => to_unsigned(29853, LUT_AMPL_WIDTH - 1),
		20817 => to_unsigned(29852, LUT_AMPL_WIDTH - 1),
		20818 => to_unsigned(29851, LUT_AMPL_WIDTH - 1),
		20819 => to_unsigned(29849, LUT_AMPL_WIDTH - 1),
		20820 => to_unsigned(29848, LUT_AMPL_WIDTH - 1),
		20821 => to_unsigned(29847, LUT_AMPL_WIDTH - 1),
		20822 => to_unsigned(29845, LUT_AMPL_WIDTH - 1),
		20823 => to_unsigned(29844, LUT_AMPL_WIDTH - 1),
		20824 => to_unsigned(29843, LUT_AMPL_WIDTH - 1),
		20825 => to_unsigned(29842, LUT_AMPL_WIDTH - 1),
		20826 => to_unsigned(29840, LUT_AMPL_WIDTH - 1),
		20827 => to_unsigned(29839, LUT_AMPL_WIDTH - 1),
		20828 => to_unsigned(29838, LUT_AMPL_WIDTH - 1),
		20829 => to_unsigned(29836, LUT_AMPL_WIDTH - 1),
		20830 => to_unsigned(29835, LUT_AMPL_WIDTH - 1),
		20831 => to_unsigned(29834, LUT_AMPL_WIDTH - 1),
		20832 => to_unsigned(29832, LUT_AMPL_WIDTH - 1),
		20833 => to_unsigned(29831, LUT_AMPL_WIDTH - 1),
		20834 => to_unsigned(29830, LUT_AMPL_WIDTH - 1),
		20835 => to_unsigned(29829, LUT_AMPL_WIDTH - 1),
		20836 => to_unsigned(29827, LUT_AMPL_WIDTH - 1),
		20837 => to_unsigned(29826, LUT_AMPL_WIDTH - 1),
		20838 => to_unsigned(29825, LUT_AMPL_WIDTH - 1),
		20839 => to_unsigned(29823, LUT_AMPL_WIDTH - 1),
		20840 => to_unsigned(29822, LUT_AMPL_WIDTH - 1),
		20841 => to_unsigned(29821, LUT_AMPL_WIDTH - 1),
		20842 => to_unsigned(29819, LUT_AMPL_WIDTH - 1),
		20843 => to_unsigned(29818, LUT_AMPL_WIDTH - 1),
		20844 => to_unsigned(29817, LUT_AMPL_WIDTH - 1),
		20845 => to_unsigned(29816, LUT_AMPL_WIDTH - 1),
		20846 => to_unsigned(29814, LUT_AMPL_WIDTH - 1),
		20847 => to_unsigned(29813, LUT_AMPL_WIDTH - 1),
		20848 => to_unsigned(29812, LUT_AMPL_WIDTH - 1),
		20849 => to_unsigned(29810, LUT_AMPL_WIDTH - 1),
		20850 => to_unsigned(29809, LUT_AMPL_WIDTH - 1),
		20851 => to_unsigned(29808, LUT_AMPL_WIDTH - 1),
		20852 => to_unsigned(29806, LUT_AMPL_WIDTH - 1),
		20853 => to_unsigned(29805, LUT_AMPL_WIDTH - 1),
		20854 => to_unsigned(29804, LUT_AMPL_WIDTH - 1),
		20855 => to_unsigned(29802, LUT_AMPL_WIDTH - 1),
		20856 => to_unsigned(29801, LUT_AMPL_WIDTH - 1),
		20857 => to_unsigned(29800, LUT_AMPL_WIDTH - 1),
		20858 => to_unsigned(29799, LUT_AMPL_WIDTH - 1),
		20859 => to_unsigned(29797, LUT_AMPL_WIDTH - 1),
		20860 => to_unsigned(29796, LUT_AMPL_WIDTH - 1),
		20861 => to_unsigned(29795, LUT_AMPL_WIDTH - 1),
		20862 => to_unsigned(29793, LUT_AMPL_WIDTH - 1),
		20863 => to_unsigned(29792, LUT_AMPL_WIDTH - 1),
		20864 => to_unsigned(29791, LUT_AMPL_WIDTH - 1),
		20865 => to_unsigned(29789, LUT_AMPL_WIDTH - 1),
		20866 => to_unsigned(29788, LUT_AMPL_WIDTH - 1),
		20867 => to_unsigned(29787, LUT_AMPL_WIDTH - 1),
		20868 => to_unsigned(29785, LUT_AMPL_WIDTH - 1),
		20869 => to_unsigned(29784, LUT_AMPL_WIDTH - 1),
		20870 => to_unsigned(29783, LUT_AMPL_WIDTH - 1),
		20871 => to_unsigned(29782, LUT_AMPL_WIDTH - 1),
		20872 => to_unsigned(29780, LUT_AMPL_WIDTH - 1),
		20873 => to_unsigned(29779, LUT_AMPL_WIDTH - 1),
		20874 => to_unsigned(29778, LUT_AMPL_WIDTH - 1),
		20875 => to_unsigned(29776, LUT_AMPL_WIDTH - 1),
		20876 => to_unsigned(29775, LUT_AMPL_WIDTH - 1),
		20877 => to_unsigned(29774, LUT_AMPL_WIDTH - 1),
		20878 => to_unsigned(29772, LUT_AMPL_WIDTH - 1),
		20879 => to_unsigned(29771, LUT_AMPL_WIDTH - 1),
		20880 => to_unsigned(29770, LUT_AMPL_WIDTH - 1),
		20881 => to_unsigned(29768, LUT_AMPL_WIDTH - 1),
		20882 => to_unsigned(29767, LUT_AMPL_WIDTH - 1),
		20883 => to_unsigned(29766, LUT_AMPL_WIDTH - 1),
		20884 => to_unsigned(29764, LUT_AMPL_WIDTH - 1),
		20885 => to_unsigned(29763, LUT_AMPL_WIDTH - 1),
		20886 => to_unsigned(29762, LUT_AMPL_WIDTH - 1),
		20887 => to_unsigned(29761, LUT_AMPL_WIDTH - 1),
		20888 => to_unsigned(29759, LUT_AMPL_WIDTH - 1),
		20889 => to_unsigned(29758, LUT_AMPL_WIDTH - 1),
		20890 => to_unsigned(29757, LUT_AMPL_WIDTH - 1),
		20891 => to_unsigned(29755, LUT_AMPL_WIDTH - 1),
		20892 => to_unsigned(29754, LUT_AMPL_WIDTH - 1),
		20893 => to_unsigned(29753, LUT_AMPL_WIDTH - 1),
		20894 => to_unsigned(29751, LUT_AMPL_WIDTH - 1),
		20895 => to_unsigned(29750, LUT_AMPL_WIDTH - 1),
		20896 => to_unsigned(29749, LUT_AMPL_WIDTH - 1),
		20897 => to_unsigned(29747, LUT_AMPL_WIDTH - 1),
		20898 => to_unsigned(29746, LUT_AMPL_WIDTH - 1),
		20899 => to_unsigned(29745, LUT_AMPL_WIDTH - 1),
		20900 => to_unsigned(29743, LUT_AMPL_WIDTH - 1),
		20901 => to_unsigned(29742, LUT_AMPL_WIDTH - 1),
		20902 => to_unsigned(29741, LUT_AMPL_WIDTH - 1),
		20903 => to_unsigned(29739, LUT_AMPL_WIDTH - 1),
		20904 => to_unsigned(29738, LUT_AMPL_WIDTH - 1),
		20905 => to_unsigned(29737, LUT_AMPL_WIDTH - 1),
		20906 => to_unsigned(29736, LUT_AMPL_WIDTH - 1),
		20907 => to_unsigned(29734, LUT_AMPL_WIDTH - 1),
		20908 => to_unsigned(29733, LUT_AMPL_WIDTH - 1),
		20909 => to_unsigned(29732, LUT_AMPL_WIDTH - 1),
		20910 => to_unsigned(29730, LUT_AMPL_WIDTH - 1),
		20911 => to_unsigned(29729, LUT_AMPL_WIDTH - 1),
		20912 => to_unsigned(29728, LUT_AMPL_WIDTH - 1),
		20913 => to_unsigned(29726, LUT_AMPL_WIDTH - 1),
		20914 => to_unsigned(29725, LUT_AMPL_WIDTH - 1),
		20915 => to_unsigned(29724, LUT_AMPL_WIDTH - 1),
		20916 => to_unsigned(29722, LUT_AMPL_WIDTH - 1),
		20917 => to_unsigned(29721, LUT_AMPL_WIDTH - 1),
		20918 => to_unsigned(29720, LUT_AMPL_WIDTH - 1),
		20919 => to_unsigned(29718, LUT_AMPL_WIDTH - 1),
		20920 => to_unsigned(29717, LUT_AMPL_WIDTH - 1),
		20921 => to_unsigned(29716, LUT_AMPL_WIDTH - 1),
		20922 => to_unsigned(29714, LUT_AMPL_WIDTH - 1),
		20923 => to_unsigned(29713, LUT_AMPL_WIDTH - 1),
		20924 => to_unsigned(29712, LUT_AMPL_WIDTH - 1),
		20925 => to_unsigned(29710, LUT_AMPL_WIDTH - 1),
		20926 => to_unsigned(29709, LUT_AMPL_WIDTH - 1),
		20927 => to_unsigned(29708, LUT_AMPL_WIDTH - 1),
		20928 => to_unsigned(29706, LUT_AMPL_WIDTH - 1),
		20929 => to_unsigned(29705, LUT_AMPL_WIDTH - 1),
		20930 => to_unsigned(29704, LUT_AMPL_WIDTH - 1),
		20931 => to_unsigned(29702, LUT_AMPL_WIDTH - 1),
		20932 => to_unsigned(29701, LUT_AMPL_WIDTH - 1),
		20933 => to_unsigned(29700, LUT_AMPL_WIDTH - 1),
		20934 => to_unsigned(29698, LUT_AMPL_WIDTH - 1),
		20935 => to_unsigned(29697, LUT_AMPL_WIDTH - 1),
		20936 => to_unsigned(29696, LUT_AMPL_WIDTH - 1),
		20937 => to_unsigned(29694, LUT_AMPL_WIDTH - 1),
		20938 => to_unsigned(29693, LUT_AMPL_WIDTH - 1),
		20939 => to_unsigned(29692, LUT_AMPL_WIDTH - 1),
		20940 => to_unsigned(29690, LUT_AMPL_WIDTH - 1),
		20941 => to_unsigned(29689, LUT_AMPL_WIDTH - 1),
		20942 => to_unsigned(29688, LUT_AMPL_WIDTH - 1),
		20943 => to_unsigned(29687, LUT_AMPL_WIDTH - 1),
		20944 => to_unsigned(29685, LUT_AMPL_WIDTH - 1),
		20945 => to_unsigned(29684, LUT_AMPL_WIDTH - 1),
		20946 => to_unsigned(29683, LUT_AMPL_WIDTH - 1),
		20947 => to_unsigned(29681, LUT_AMPL_WIDTH - 1),
		20948 => to_unsigned(29680, LUT_AMPL_WIDTH - 1),
		20949 => to_unsigned(29679, LUT_AMPL_WIDTH - 1),
		20950 => to_unsigned(29677, LUT_AMPL_WIDTH - 1),
		20951 => to_unsigned(29676, LUT_AMPL_WIDTH - 1),
		20952 => to_unsigned(29675, LUT_AMPL_WIDTH - 1),
		20953 => to_unsigned(29673, LUT_AMPL_WIDTH - 1),
		20954 => to_unsigned(29672, LUT_AMPL_WIDTH - 1),
		20955 => to_unsigned(29671, LUT_AMPL_WIDTH - 1),
		20956 => to_unsigned(29669, LUT_AMPL_WIDTH - 1),
		20957 => to_unsigned(29668, LUT_AMPL_WIDTH - 1),
		20958 => to_unsigned(29667, LUT_AMPL_WIDTH - 1),
		20959 => to_unsigned(29665, LUT_AMPL_WIDTH - 1),
		20960 => to_unsigned(29664, LUT_AMPL_WIDTH - 1),
		20961 => to_unsigned(29663, LUT_AMPL_WIDTH - 1),
		20962 => to_unsigned(29661, LUT_AMPL_WIDTH - 1),
		20963 => to_unsigned(29660, LUT_AMPL_WIDTH - 1),
		20964 => to_unsigned(29659, LUT_AMPL_WIDTH - 1),
		20965 => to_unsigned(29657, LUT_AMPL_WIDTH - 1),
		20966 => to_unsigned(29656, LUT_AMPL_WIDTH - 1),
		20967 => to_unsigned(29655, LUT_AMPL_WIDTH - 1),
		20968 => to_unsigned(29653, LUT_AMPL_WIDTH - 1),
		20969 => to_unsigned(29652, LUT_AMPL_WIDTH - 1),
		20970 => to_unsigned(29651, LUT_AMPL_WIDTH - 1),
		20971 => to_unsigned(29649, LUT_AMPL_WIDTH - 1),
		20972 => to_unsigned(29648, LUT_AMPL_WIDTH - 1),
		20973 => to_unsigned(29646, LUT_AMPL_WIDTH - 1),
		20974 => to_unsigned(29645, LUT_AMPL_WIDTH - 1),
		20975 => to_unsigned(29644, LUT_AMPL_WIDTH - 1),
		20976 => to_unsigned(29642, LUT_AMPL_WIDTH - 1),
		20977 => to_unsigned(29641, LUT_AMPL_WIDTH - 1),
		20978 => to_unsigned(29640, LUT_AMPL_WIDTH - 1),
		20979 => to_unsigned(29638, LUT_AMPL_WIDTH - 1),
		20980 => to_unsigned(29637, LUT_AMPL_WIDTH - 1),
		20981 => to_unsigned(29636, LUT_AMPL_WIDTH - 1),
		20982 => to_unsigned(29634, LUT_AMPL_WIDTH - 1),
		20983 => to_unsigned(29633, LUT_AMPL_WIDTH - 1),
		20984 => to_unsigned(29632, LUT_AMPL_WIDTH - 1),
		20985 => to_unsigned(29630, LUT_AMPL_WIDTH - 1),
		20986 => to_unsigned(29629, LUT_AMPL_WIDTH - 1),
		20987 => to_unsigned(29628, LUT_AMPL_WIDTH - 1),
		20988 => to_unsigned(29626, LUT_AMPL_WIDTH - 1),
		20989 => to_unsigned(29625, LUT_AMPL_WIDTH - 1),
		20990 => to_unsigned(29624, LUT_AMPL_WIDTH - 1),
		20991 => to_unsigned(29622, LUT_AMPL_WIDTH - 1),
		20992 => to_unsigned(29621, LUT_AMPL_WIDTH - 1),
		20993 => to_unsigned(29620, LUT_AMPL_WIDTH - 1),
		20994 => to_unsigned(29618, LUT_AMPL_WIDTH - 1),
		20995 => to_unsigned(29617, LUT_AMPL_WIDTH - 1),
		20996 => to_unsigned(29616, LUT_AMPL_WIDTH - 1),
		20997 => to_unsigned(29614, LUT_AMPL_WIDTH - 1),
		20998 => to_unsigned(29613, LUT_AMPL_WIDTH - 1),
		20999 => to_unsigned(29612, LUT_AMPL_WIDTH - 1),
		21000 => to_unsigned(29610, LUT_AMPL_WIDTH - 1),
		21001 => to_unsigned(29609, LUT_AMPL_WIDTH - 1),
		21002 => to_unsigned(29608, LUT_AMPL_WIDTH - 1),
		21003 => to_unsigned(29606, LUT_AMPL_WIDTH - 1),
		21004 => to_unsigned(29605, LUT_AMPL_WIDTH - 1),
		21005 => to_unsigned(29604, LUT_AMPL_WIDTH - 1),
		21006 => to_unsigned(29602, LUT_AMPL_WIDTH - 1),
		21007 => to_unsigned(29601, LUT_AMPL_WIDTH - 1),
		21008 => to_unsigned(29599, LUT_AMPL_WIDTH - 1),
		21009 => to_unsigned(29598, LUT_AMPL_WIDTH - 1),
		21010 => to_unsigned(29597, LUT_AMPL_WIDTH - 1),
		21011 => to_unsigned(29595, LUT_AMPL_WIDTH - 1),
		21012 => to_unsigned(29594, LUT_AMPL_WIDTH - 1),
		21013 => to_unsigned(29593, LUT_AMPL_WIDTH - 1),
		21014 => to_unsigned(29591, LUT_AMPL_WIDTH - 1),
		21015 => to_unsigned(29590, LUT_AMPL_WIDTH - 1),
		21016 => to_unsigned(29589, LUT_AMPL_WIDTH - 1),
		21017 => to_unsigned(29587, LUT_AMPL_WIDTH - 1),
		21018 => to_unsigned(29586, LUT_AMPL_WIDTH - 1),
		21019 => to_unsigned(29585, LUT_AMPL_WIDTH - 1),
		21020 => to_unsigned(29583, LUT_AMPL_WIDTH - 1),
		21021 => to_unsigned(29582, LUT_AMPL_WIDTH - 1),
		21022 => to_unsigned(29581, LUT_AMPL_WIDTH - 1),
		21023 => to_unsigned(29579, LUT_AMPL_WIDTH - 1),
		21024 => to_unsigned(29578, LUT_AMPL_WIDTH - 1),
		21025 => to_unsigned(29577, LUT_AMPL_WIDTH - 1),
		21026 => to_unsigned(29575, LUT_AMPL_WIDTH - 1),
		21027 => to_unsigned(29574, LUT_AMPL_WIDTH - 1),
		21028 => to_unsigned(29572, LUT_AMPL_WIDTH - 1),
		21029 => to_unsigned(29571, LUT_AMPL_WIDTH - 1),
		21030 => to_unsigned(29570, LUT_AMPL_WIDTH - 1),
		21031 => to_unsigned(29568, LUT_AMPL_WIDTH - 1),
		21032 => to_unsigned(29567, LUT_AMPL_WIDTH - 1),
		21033 => to_unsigned(29566, LUT_AMPL_WIDTH - 1),
		21034 => to_unsigned(29564, LUT_AMPL_WIDTH - 1),
		21035 => to_unsigned(29563, LUT_AMPL_WIDTH - 1),
		21036 => to_unsigned(29562, LUT_AMPL_WIDTH - 1),
		21037 => to_unsigned(29560, LUT_AMPL_WIDTH - 1),
		21038 => to_unsigned(29559, LUT_AMPL_WIDTH - 1),
		21039 => to_unsigned(29558, LUT_AMPL_WIDTH - 1),
		21040 => to_unsigned(29556, LUT_AMPL_WIDTH - 1),
		21041 => to_unsigned(29555, LUT_AMPL_WIDTH - 1),
		21042 => to_unsigned(29554, LUT_AMPL_WIDTH - 1),
		21043 => to_unsigned(29552, LUT_AMPL_WIDTH - 1),
		21044 => to_unsigned(29551, LUT_AMPL_WIDTH - 1),
		21045 => to_unsigned(29549, LUT_AMPL_WIDTH - 1),
		21046 => to_unsigned(29548, LUT_AMPL_WIDTH - 1),
		21047 => to_unsigned(29547, LUT_AMPL_WIDTH - 1),
		21048 => to_unsigned(29545, LUT_AMPL_WIDTH - 1),
		21049 => to_unsigned(29544, LUT_AMPL_WIDTH - 1),
		21050 => to_unsigned(29543, LUT_AMPL_WIDTH - 1),
		21051 => to_unsigned(29541, LUT_AMPL_WIDTH - 1),
		21052 => to_unsigned(29540, LUT_AMPL_WIDTH - 1),
		21053 => to_unsigned(29539, LUT_AMPL_WIDTH - 1),
		21054 => to_unsigned(29537, LUT_AMPL_WIDTH - 1),
		21055 => to_unsigned(29536, LUT_AMPL_WIDTH - 1),
		21056 => to_unsigned(29534, LUT_AMPL_WIDTH - 1),
		21057 => to_unsigned(29533, LUT_AMPL_WIDTH - 1),
		21058 => to_unsigned(29532, LUT_AMPL_WIDTH - 1),
		21059 => to_unsigned(29530, LUT_AMPL_WIDTH - 1),
		21060 => to_unsigned(29529, LUT_AMPL_WIDTH - 1),
		21061 => to_unsigned(29528, LUT_AMPL_WIDTH - 1),
		21062 => to_unsigned(29526, LUT_AMPL_WIDTH - 1),
		21063 => to_unsigned(29525, LUT_AMPL_WIDTH - 1),
		21064 => to_unsigned(29524, LUT_AMPL_WIDTH - 1),
		21065 => to_unsigned(29522, LUT_AMPL_WIDTH - 1),
		21066 => to_unsigned(29521, LUT_AMPL_WIDTH - 1),
		21067 => to_unsigned(29520, LUT_AMPL_WIDTH - 1),
		21068 => to_unsigned(29518, LUT_AMPL_WIDTH - 1),
		21069 => to_unsigned(29517, LUT_AMPL_WIDTH - 1),
		21070 => to_unsigned(29515, LUT_AMPL_WIDTH - 1),
		21071 => to_unsigned(29514, LUT_AMPL_WIDTH - 1),
		21072 => to_unsigned(29513, LUT_AMPL_WIDTH - 1),
		21073 => to_unsigned(29511, LUT_AMPL_WIDTH - 1),
		21074 => to_unsigned(29510, LUT_AMPL_WIDTH - 1),
		21075 => to_unsigned(29509, LUT_AMPL_WIDTH - 1),
		21076 => to_unsigned(29507, LUT_AMPL_WIDTH - 1),
		21077 => to_unsigned(29506, LUT_AMPL_WIDTH - 1),
		21078 => to_unsigned(29504, LUT_AMPL_WIDTH - 1),
		21079 => to_unsigned(29503, LUT_AMPL_WIDTH - 1),
		21080 => to_unsigned(29502, LUT_AMPL_WIDTH - 1),
		21081 => to_unsigned(29500, LUT_AMPL_WIDTH - 1),
		21082 => to_unsigned(29499, LUT_AMPL_WIDTH - 1),
		21083 => to_unsigned(29498, LUT_AMPL_WIDTH - 1),
		21084 => to_unsigned(29496, LUT_AMPL_WIDTH - 1),
		21085 => to_unsigned(29495, LUT_AMPL_WIDTH - 1),
		21086 => to_unsigned(29494, LUT_AMPL_WIDTH - 1),
		21087 => to_unsigned(29492, LUT_AMPL_WIDTH - 1),
		21088 => to_unsigned(29491, LUT_AMPL_WIDTH - 1),
		21089 => to_unsigned(29489, LUT_AMPL_WIDTH - 1),
		21090 => to_unsigned(29488, LUT_AMPL_WIDTH - 1),
		21091 => to_unsigned(29487, LUT_AMPL_WIDTH - 1),
		21092 => to_unsigned(29485, LUT_AMPL_WIDTH - 1),
		21093 => to_unsigned(29484, LUT_AMPL_WIDTH - 1),
		21094 => to_unsigned(29483, LUT_AMPL_WIDTH - 1),
		21095 => to_unsigned(29481, LUT_AMPL_WIDTH - 1),
		21096 => to_unsigned(29480, LUT_AMPL_WIDTH - 1),
		21097 => to_unsigned(29478, LUT_AMPL_WIDTH - 1),
		21098 => to_unsigned(29477, LUT_AMPL_WIDTH - 1),
		21099 => to_unsigned(29476, LUT_AMPL_WIDTH - 1),
		21100 => to_unsigned(29474, LUT_AMPL_WIDTH - 1),
		21101 => to_unsigned(29473, LUT_AMPL_WIDTH - 1),
		21102 => to_unsigned(29472, LUT_AMPL_WIDTH - 1),
		21103 => to_unsigned(29470, LUT_AMPL_WIDTH - 1),
		21104 => to_unsigned(29469, LUT_AMPL_WIDTH - 1),
		21105 => to_unsigned(29468, LUT_AMPL_WIDTH - 1),
		21106 => to_unsigned(29466, LUT_AMPL_WIDTH - 1),
		21107 => to_unsigned(29465, LUT_AMPL_WIDTH - 1),
		21108 => to_unsigned(29463, LUT_AMPL_WIDTH - 1),
		21109 => to_unsigned(29462, LUT_AMPL_WIDTH - 1),
		21110 => to_unsigned(29461, LUT_AMPL_WIDTH - 1),
		21111 => to_unsigned(29459, LUT_AMPL_WIDTH - 1),
		21112 => to_unsigned(29458, LUT_AMPL_WIDTH - 1),
		21113 => to_unsigned(29457, LUT_AMPL_WIDTH - 1),
		21114 => to_unsigned(29455, LUT_AMPL_WIDTH - 1),
		21115 => to_unsigned(29454, LUT_AMPL_WIDTH - 1),
		21116 => to_unsigned(29452, LUT_AMPL_WIDTH - 1),
		21117 => to_unsigned(29451, LUT_AMPL_WIDTH - 1),
		21118 => to_unsigned(29450, LUT_AMPL_WIDTH - 1),
		21119 => to_unsigned(29448, LUT_AMPL_WIDTH - 1),
		21120 => to_unsigned(29447, LUT_AMPL_WIDTH - 1),
		21121 => to_unsigned(29445, LUT_AMPL_WIDTH - 1),
		21122 => to_unsigned(29444, LUT_AMPL_WIDTH - 1),
		21123 => to_unsigned(29443, LUT_AMPL_WIDTH - 1),
		21124 => to_unsigned(29441, LUT_AMPL_WIDTH - 1),
		21125 => to_unsigned(29440, LUT_AMPL_WIDTH - 1),
		21126 => to_unsigned(29439, LUT_AMPL_WIDTH - 1),
		21127 => to_unsigned(29437, LUT_AMPL_WIDTH - 1),
		21128 => to_unsigned(29436, LUT_AMPL_WIDTH - 1),
		21129 => to_unsigned(29434, LUT_AMPL_WIDTH - 1),
		21130 => to_unsigned(29433, LUT_AMPL_WIDTH - 1),
		21131 => to_unsigned(29432, LUT_AMPL_WIDTH - 1),
		21132 => to_unsigned(29430, LUT_AMPL_WIDTH - 1),
		21133 => to_unsigned(29429, LUT_AMPL_WIDTH - 1),
		21134 => to_unsigned(29428, LUT_AMPL_WIDTH - 1),
		21135 => to_unsigned(29426, LUT_AMPL_WIDTH - 1),
		21136 => to_unsigned(29425, LUT_AMPL_WIDTH - 1),
		21137 => to_unsigned(29423, LUT_AMPL_WIDTH - 1),
		21138 => to_unsigned(29422, LUT_AMPL_WIDTH - 1),
		21139 => to_unsigned(29421, LUT_AMPL_WIDTH - 1),
		21140 => to_unsigned(29419, LUT_AMPL_WIDTH - 1),
		21141 => to_unsigned(29418, LUT_AMPL_WIDTH - 1),
		21142 => to_unsigned(29416, LUT_AMPL_WIDTH - 1),
		21143 => to_unsigned(29415, LUT_AMPL_WIDTH - 1),
		21144 => to_unsigned(29414, LUT_AMPL_WIDTH - 1),
		21145 => to_unsigned(29412, LUT_AMPL_WIDTH - 1),
		21146 => to_unsigned(29411, LUT_AMPL_WIDTH - 1),
		21147 => to_unsigned(29410, LUT_AMPL_WIDTH - 1),
		21148 => to_unsigned(29408, LUT_AMPL_WIDTH - 1),
		21149 => to_unsigned(29407, LUT_AMPL_WIDTH - 1),
		21150 => to_unsigned(29405, LUT_AMPL_WIDTH - 1),
		21151 => to_unsigned(29404, LUT_AMPL_WIDTH - 1),
		21152 => to_unsigned(29403, LUT_AMPL_WIDTH - 1),
		21153 => to_unsigned(29401, LUT_AMPL_WIDTH - 1),
		21154 => to_unsigned(29400, LUT_AMPL_WIDTH - 1),
		21155 => to_unsigned(29398, LUT_AMPL_WIDTH - 1),
		21156 => to_unsigned(29397, LUT_AMPL_WIDTH - 1),
		21157 => to_unsigned(29396, LUT_AMPL_WIDTH - 1),
		21158 => to_unsigned(29394, LUT_AMPL_WIDTH - 1),
		21159 => to_unsigned(29393, LUT_AMPL_WIDTH - 1),
		21160 => to_unsigned(29392, LUT_AMPL_WIDTH - 1),
		21161 => to_unsigned(29390, LUT_AMPL_WIDTH - 1),
		21162 => to_unsigned(29389, LUT_AMPL_WIDTH - 1),
		21163 => to_unsigned(29387, LUT_AMPL_WIDTH - 1),
		21164 => to_unsigned(29386, LUT_AMPL_WIDTH - 1),
		21165 => to_unsigned(29385, LUT_AMPL_WIDTH - 1),
		21166 => to_unsigned(29383, LUT_AMPL_WIDTH - 1),
		21167 => to_unsigned(29382, LUT_AMPL_WIDTH - 1),
		21168 => to_unsigned(29380, LUT_AMPL_WIDTH - 1),
		21169 => to_unsigned(29379, LUT_AMPL_WIDTH - 1),
		21170 => to_unsigned(29378, LUT_AMPL_WIDTH - 1),
		21171 => to_unsigned(29376, LUT_AMPL_WIDTH - 1),
		21172 => to_unsigned(29375, LUT_AMPL_WIDTH - 1),
		21173 => to_unsigned(29373, LUT_AMPL_WIDTH - 1),
		21174 => to_unsigned(29372, LUT_AMPL_WIDTH - 1),
		21175 => to_unsigned(29371, LUT_AMPL_WIDTH - 1),
		21176 => to_unsigned(29369, LUT_AMPL_WIDTH - 1),
		21177 => to_unsigned(29368, LUT_AMPL_WIDTH - 1),
		21178 => to_unsigned(29366, LUT_AMPL_WIDTH - 1),
		21179 => to_unsigned(29365, LUT_AMPL_WIDTH - 1),
		21180 => to_unsigned(29364, LUT_AMPL_WIDTH - 1),
		21181 => to_unsigned(29362, LUT_AMPL_WIDTH - 1),
		21182 => to_unsigned(29361, LUT_AMPL_WIDTH - 1),
		21183 => to_unsigned(29360, LUT_AMPL_WIDTH - 1),
		21184 => to_unsigned(29358, LUT_AMPL_WIDTH - 1),
		21185 => to_unsigned(29357, LUT_AMPL_WIDTH - 1),
		21186 => to_unsigned(29355, LUT_AMPL_WIDTH - 1),
		21187 => to_unsigned(29354, LUT_AMPL_WIDTH - 1),
		21188 => to_unsigned(29353, LUT_AMPL_WIDTH - 1),
		21189 => to_unsigned(29351, LUT_AMPL_WIDTH - 1),
		21190 => to_unsigned(29350, LUT_AMPL_WIDTH - 1),
		21191 => to_unsigned(29348, LUT_AMPL_WIDTH - 1),
		21192 => to_unsigned(29347, LUT_AMPL_WIDTH - 1),
		21193 => to_unsigned(29346, LUT_AMPL_WIDTH - 1),
		21194 => to_unsigned(29344, LUT_AMPL_WIDTH - 1),
		21195 => to_unsigned(29343, LUT_AMPL_WIDTH - 1),
		21196 => to_unsigned(29341, LUT_AMPL_WIDTH - 1),
		21197 => to_unsigned(29340, LUT_AMPL_WIDTH - 1),
		21198 => to_unsigned(29339, LUT_AMPL_WIDTH - 1),
		21199 => to_unsigned(29337, LUT_AMPL_WIDTH - 1),
		21200 => to_unsigned(29336, LUT_AMPL_WIDTH - 1),
		21201 => to_unsigned(29334, LUT_AMPL_WIDTH - 1),
		21202 => to_unsigned(29333, LUT_AMPL_WIDTH - 1),
		21203 => to_unsigned(29332, LUT_AMPL_WIDTH - 1),
		21204 => to_unsigned(29330, LUT_AMPL_WIDTH - 1),
		21205 => to_unsigned(29329, LUT_AMPL_WIDTH - 1),
		21206 => to_unsigned(29327, LUT_AMPL_WIDTH - 1),
		21207 => to_unsigned(29326, LUT_AMPL_WIDTH - 1),
		21208 => to_unsigned(29325, LUT_AMPL_WIDTH - 1),
		21209 => to_unsigned(29323, LUT_AMPL_WIDTH - 1),
		21210 => to_unsigned(29322, LUT_AMPL_WIDTH - 1),
		21211 => to_unsigned(29320, LUT_AMPL_WIDTH - 1),
		21212 => to_unsigned(29319, LUT_AMPL_WIDTH - 1),
		21213 => to_unsigned(29318, LUT_AMPL_WIDTH - 1),
		21214 => to_unsigned(29316, LUT_AMPL_WIDTH - 1),
		21215 => to_unsigned(29315, LUT_AMPL_WIDTH - 1),
		21216 => to_unsigned(29313, LUT_AMPL_WIDTH - 1),
		21217 => to_unsigned(29312, LUT_AMPL_WIDTH - 1),
		21218 => to_unsigned(29311, LUT_AMPL_WIDTH - 1),
		21219 => to_unsigned(29309, LUT_AMPL_WIDTH - 1),
		21220 => to_unsigned(29308, LUT_AMPL_WIDTH - 1),
		21221 => to_unsigned(29306, LUT_AMPL_WIDTH - 1),
		21222 => to_unsigned(29305, LUT_AMPL_WIDTH - 1),
		21223 => to_unsigned(29304, LUT_AMPL_WIDTH - 1),
		21224 => to_unsigned(29302, LUT_AMPL_WIDTH - 1),
		21225 => to_unsigned(29301, LUT_AMPL_WIDTH - 1),
		21226 => to_unsigned(29299, LUT_AMPL_WIDTH - 1),
		21227 => to_unsigned(29298, LUT_AMPL_WIDTH - 1),
		21228 => to_unsigned(29296, LUT_AMPL_WIDTH - 1),
		21229 => to_unsigned(29295, LUT_AMPL_WIDTH - 1),
		21230 => to_unsigned(29294, LUT_AMPL_WIDTH - 1),
		21231 => to_unsigned(29292, LUT_AMPL_WIDTH - 1),
		21232 => to_unsigned(29291, LUT_AMPL_WIDTH - 1),
		21233 => to_unsigned(29289, LUT_AMPL_WIDTH - 1),
		21234 => to_unsigned(29288, LUT_AMPL_WIDTH - 1),
		21235 => to_unsigned(29287, LUT_AMPL_WIDTH - 1),
		21236 => to_unsigned(29285, LUT_AMPL_WIDTH - 1),
		21237 => to_unsigned(29284, LUT_AMPL_WIDTH - 1),
		21238 => to_unsigned(29282, LUT_AMPL_WIDTH - 1),
		21239 => to_unsigned(29281, LUT_AMPL_WIDTH - 1),
		21240 => to_unsigned(29280, LUT_AMPL_WIDTH - 1),
		21241 => to_unsigned(29278, LUT_AMPL_WIDTH - 1),
		21242 => to_unsigned(29277, LUT_AMPL_WIDTH - 1),
		21243 => to_unsigned(29275, LUT_AMPL_WIDTH - 1),
		21244 => to_unsigned(29274, LUT_AMPL_WIDTH - 1),
		21245 => to_unsigned(29273, LUT_AMPL_WIDTH - 1),
		21246 => to_unsigned(29271, LUT_AMPL_WIDTH - 1),
		21247 => to_unsigned(29270, LUT_AMPL_WIDTH - 1),
		21248 => to_unsigned(29268, LUT_AMPL_WIDTH - 1),
		21249 => to_unsigned(29267, LUT_AMPL_WIDTH - 1),
		21250 => to_unsigned(29265, LUT_AMPL_WIDTH - 1),
		21251 => to_unsigned(29264, LUT_AMPL_WIDTH - 1),
		21252 => to_unsigned(29263, LUT_AMPL_WIDTH - 1),
		21253 => to_unsigned(29261, LUT_AMPL_WIDTH - 1),
		21254 => to_unsigned(29260, LUT_AMPL_WIDTH - 1),
		21255 => to_unsigned(29258, LUT_AMPL_WIDTH - 1),
		21256 => to_unsigned(29257, LUT_AMPL_WIDTH - 1),
		21257 => to_unsigned(29256, LUT_AMPL_WIDTH - 1),
		21258 => to_unsigned(29254, LUT_AMPL_WIDTH - 1),
		21259 => to_unsigned(29253, LUT_AMPL_WIDTH - 1),
		21260 => to_unsigned(29251, LUT_AMPL_WIDTH - 1),
		21261 => to_unsigned(29250, LUT_AMPL_WIDTH - 1),
		21262 => to_unsigned(29248, LUT_AMPL_WIDTH - 1),
		21263 => to_unsigned(29247, LUT_AMPL_WIDTH - 1),
		21264 => to_unsigned(29246, LUT_AMPL_WIDTH - 1),
		21265 => to_unsigned(29244, LUT_AMPL_WIDTH - 1),
		21266 => to_unsigned(29243, LUT_AMPL_WIDTH - 1),
		21267 => to_unsigned(29241, LUT_AMPL_WIDTH - 1),
		21268 => to_unsigned(29240, LUT_AMPL_WIDTH - 1),
		21269 => to_unsigned(29239, LUT_AMPL_WIDTH - 1),
		21270 => to_unsigned(29237, LUT_AMPL_WIDTH - 1),
		21271 => to_unsigned(29236, LUT_AMPL_WIDTH - 1),
		21272 => to_unsigned(29234, LUT_AMPL_WIDTH - 1),
		21273 => to_unsigned(29233, LUT_AMPL_WIDTH - 1),
		21274 => to_unsigned(29231, LUT_AMPL_WIDTH - 1),
		21275 => to_unsigned(29230, LUT_AMPL_WIDTH - 1),
		21276 => to_unsigned(29229, LUT_AMPL_WIDTH - 1),
		21277 => to_unsigned(29227, LUT_AMPL_WIDTH - 1),
		21278 => to_unsigned(29226, LUT_AMPL_WIDTH - 1),
		21279 => to_unsigned(29224, LUT_AMPL_WIDTH - 1),
		21280 => to_unsigned(29223, LUT_AMPL_WIDTH - 1),
		21281 => to_unsigned(29222, LUT_AMPL_WIDTH - 1),
		21282 => to_unsigned(29220, LUT_AMPL_WIDTH - 1),
		21283 => to_unsigned(29219, LUT_AMPL_WIDTH - 1),
		21284 => to_unsigned(29217, LUT_AMPL_WIDTH - 1),
		21285 => to_unsigned(29216, LUT_AMPL_WIDTH - 1),
		21286 => to_unsigned(29214, LUT_AMPL_WIDTH - 1),
		21287 => to_unsigned(29213, LUT_AMPL_WIDTH - 1),
		21288 => to_unsigned(29212, LUT_AMPL_WIDTH - 1),
		21289 => to_unsigned(29210, LUT_AMPL_WIDTH - 1),
		21290 => to_unsigned(29209, LUT_AMPL_WIDTH - 1),
		21291 => to_unsigned(29207, LUT_AMPL_WIDTH - 1),
		21292 => to_unsigned(29206, LUT_AMPL_WIDTH - 1),
		21293 => to_unsigned(29204, LUT_AMPL_WIDTH - 1),
		21294 => to_unsigned(29203, LUT_AMPL_WIDTH - 1),
		21295 => to_unsigned(29202, LUT_AMPL_WIDTH - 1),
		21296 => to_unsigned(29200, LUT_AMPL_WIDTH - 1),
		21297 => to_unsigned(29199, LUT_AMPL_WIDTH - 1),
		21298 => to_unsigned(29197, LUT_AMPL_WIDTH - 1),
		21299 => to_unsigned(29196, LUT_AMPL_WIDTH - 1),
		21300 => to_unsigned(29194, LUT_AMPL_WIDTH - 1),
		21301 => to_unsigned(29193, LUT_AMPL_WIDTH - 1),
		21302 => to_unsigned(29192, LUT_AMPL_WIDTH - 1),
		21303 => to_unsigned(29190, LUT_AMPL_WIDTH - 1),
		21304 => to_unsigned(29189, LUT_AMPL_WIDTH - 1),
		21305 => to_unsigned(29187, LUT_AMPL_WIDTH - 1),
		21306 => to_unsigned(29186, LUT_AMPL_WIDTH - 1),
		21307 => to_unsigned(29184, LUT_AMPL_WIDTH - 1),
		21308 => to_unsigned(29183, LUT_AMPL_WIDTH - 1),
		21309 => to_unsigned(29182, LUT_AMPL_WIDTH - 1),
		21310 => to_unsigned(29180, LUT_AMPL_WIDTH - 1),
		21311 => to_unsigned(29179, LUT_AMPL_WIDTH - 1),
		21312 => to_unsigned(29177, LUT_AMPL_WIDTH - 1),
		21313 => to_unsigned(29176, LUT_AMPL_WIDTH - 1),
		21314 => to_unsigned(29174, LUT_AMPL_WIDTH - 1),
		21315 => to_unsigned(29173, LUT_AMPL_WIDTH - 1),
		21316 => to_unsigned(29172, LUT_AMPL_WIDTH - 1),
		21317 => to_unsigned(29170, LUT_AMPL_WIDTH - 1),
		21318 => to_unsigned(29169, LUT_AMPL_WIDTH - 1),
		21319 => to_unsigned(29167, LUT_AMPL_WIDTH - 1),
		21320 => to_unsigned(29166, LUT_AMPL_WIDTH - 1),
		21321 => to_unsigned(29164, LUT_AMPL_WIDTH - 1),
		21322 => to_unsigned(29163, LUT_AMPL_WIDTH - 1),
		21323 => to_unsigned(29162, LUT_AMPL_WIDTH - 1),
		21324 => to_unsigned(29160, LUT_AMPL_WIDTH - 1),
		21325 => to_unsigned(29159, LUT_AMPL_WIDTH - 1),
		21326 => to_unsigned(29157, LUT_AMPL_WIDTH - 1),
		21327 => to_unsigned(29156, LUT_AMPL_WIDTH - 1),
		21328 => to_unsigned(29154, LUT_AMPL_WIDTH - 1),
		21329 => to_unsigned(29153, LUT_AMPL_WIDTH - 1),
		21330 => to_unsigned(29152, LUT_AMPL_WIDTH - 1),
		21331 => to_unsigned(29150, LUT_AMPL_WIDTH - 1),
		21332 => to_unsigned(29149, LUT_AMPL_WIDTH - 1),
		21333 => to_unsigned(29147, LUT_AMPL_WIDTH - 1),
		21334 => to_unsigned(29146, LUT_AMPL_WIDTH - 1),
		21335 => to_unsigned(29144, LUT_AMPL_WIDTH - 1),
		21336 => to_unsigned(29143, LUT_AMPL_WIDTH - 1),
		21337 => to_unsigned(29142, LUT_AMPL_WIDTH - 1),
		21338 => to_unsigned(29140, LUT_AMPL_WIDTH - 1),
		21339 => to_unsigned(29139, LUT_AMPL_WIDTH - 1),
		21340 => to_unsigned(29137, LUT_AMPL_WIDTH - 1),
		21341 => to_unsigned(29136, LUT_AMPL_WIDTH - 1),
		21342 => to_unsigned(29134, LUT_AMPL_WIDTH - 1),
		21343 => to_unsigned(29133, LUT_AMPL_WIDTH - 1),
		21344 => to_unsigned(29131, LUT_AMPL_WIDTH - 1),
		21345 => to_unsigned(29130, LUT_AMPL_WIDTH - 1),
		21346 => to_unsigned(29129, LUT_AMPL_WIDTH - 1),
		21347 => to_unsigned(29127, LUT_AMPL_WIDTH - 1),
		21348 => to_unsigned(29126, LUT_AMPL_WIDTH - 1),
		21349 => to_unsigned(29124, LUT_AMPL_WIDTH - 1),
		21350 => to_unsigned(29123, LUT_AMPL_WIDTH - 1),
		21351 => to_unsigned(29121, LUT_AMPL_WIDTH - 1),
		21352 => to_unsigned(29120, LUT_AMPL_WIDTH - 1),
		21353 => to_unsigned(29118, LUT_AMPL_WIDTH - 1),
		21354 => to_unsigned(29117, LUT_AMPL_WIDTH - 1),
		21355 => to_unsigned(29116, LUT_AMPL_WIDTH - 1),
		21356 => to_unsigned(29114, LUT_AMPL_WIDTH - 1),
		21357 => to_unsigned(29113, LUT_AMPL_WIDTH - 1),
		21358 => to_unsigned(29111, LUT_AMPL_WIDTH - 1),
		21359 => to_unsigned(29110, LUT_AMPL_WIDTH - 1),
		21360 => to_unsigned(29108, LUT_AMPL_WIDTH - 1),
		21361 => to_unsigned(29107, LUT_AMPL_WIDTH - 1),
		21362 => to_unsigned(29106, LUT_AMPL_WIDTH - 1),
		21363 => to_unsigned(29104, LUT_AMPL_WIDTH - 1),
		21364 => to_unsigned(29103, LUT_AMPL_WIDTH - 1),
		21365 => to_unsigned(29101, LUT_AMPL_WIDTH - 1),
		21366 => to_unsigned(29100, LUT_AMPL_WIDTH - 1),
		21367 => to_unsigned(29098, LUT_AMPL_WIDTH - 1),
		21368 => to_unsigned(29097, LUT_AMPL_WIDTH - 1),
		21369 => to_unsigned(29095, LUT_AMPL_WIDTH - 1),
		21370 => to_unsigned(29094, LUT_AMPL_WIDTH - 1),
		21371 => to_unsigned(29093, LUT_AMPL_WIDTH - 1),
		21372 => to_unsigned(29091, LUT_AMPL_WIDTH - 1),
		21373 => to_unsigned(29090, LUT_AMPL_WIDTH - 1),
		21374 => to_unsigned(29088, LUT_AMPL_WIDTH - 1),
		21375 => to_unsigned(29087, LUT_AMPL_WIDTH - 1),
		21376 => to_unsigned(29085, LUT_AMPL_WIDTH - 1),
		21377 => to_unsigned(29084, LUT_AMPL_WIDTH - 1),
		21378 => to_unsigned(29082, LUT_AMPL_WIDTH - 1),
		21379 => to_unsigned(29081, LUT_AMPL_WIDTH - 1),
		21380 => to_unsigned(29079, LUT_AMPL_WIDTH - 1),
		21381 => to_unsigned(29078, LUT_AMPL_WIDTH - 1),
		21382 => to_unsigned(29077, LUT_AMPL_WIDTH - 1),
		21383 => to_unsigned(29075, LUT_AMPL_WIDTH - 1),
		21384 => to_unsigned(29074, LUT_AMPL_WIDTH - 1),
		21385 => to_unsigned(29072, LUT_AMPL_WIDTH - 1),
		21386 => to_unsigned(29071, LUT_AMPL_WIDTH - 1),
		21387 => to_unsigned(29069, LUT_AMPL_WIDTH - 1),
		21388 => to_unsigned(29068, LUT_AMPL_WIDTH - 1),
		21389 => to_unsigned(29066, LUT_AMPL_WIDTH - 1),
		21390 => to_unsigned(29065, LUT_AMPL_WIDTH - 1),
		21391 => to_unsigned(29064, LUT_AMPL_WIDTH - 1),
		21392 => to_unsigned(29062, LUT_AMPL_WIDTH - 1),
		21393 => to_unsigned(29061, LUT_AMPL_WIDTH - 1),
		21394 => to_unsigned(29059, LUT_AMPL_WIDTH - 1),
		21395 => to_unsigned(29058, LUT_AMPL_WIDTH - 1),
		21396 => to_unsigned(29056, LUT_AMPL_WIDTH - 1),
		21397 => to_unsigned(29055, LUT_AMPL_WIDTH - 1),
		21398 => to_unsigned(29053, LUT_AMPL_WIDTH - 1),
		21399 => to_unsigned(29052, LUT_AMPL_WIDTH - 1),
		21400 => to_unsigned(29050, LUT_AMPL_WIDTH - 1),
		21401 => to_unsigned(29049, LUT_AMPL_WIDTH - 1),
		21402 => to_unsigned(29048, LUT_AMPL_WIDTH - 1),
		21403 => to_unsigned(29046, LUT_AMPL_WIDTH - 1),
		21404 => to_unsigned(29045, LUT_AMPL_WIDTH - 1),
		21405 => to_unsigned(29043, LUT_AMPL_WIDTH - 1),
		21406 => to_unsigned(29042, LUT_AMPL_WIDTH - 1),
		21407 => to_unsigned(29040, LUT_AMPL_WIDTH - 1),
		21408 => to_unsigned(29039, LUT_AMPL_WIDTH - 1),
		21409 => to_unsigned(29037, LUT_AMPL_WIDTH - 1),
		21410 => to_unsigned(29036, LUT_AMPL_WIDTH - 1),
		21411 => to_unsigned(29034, LUT_AMPL_WIDTH - 1),
		21412 => to_unsigned(29033, LUT_AMPL_WIDTH - 1),
		21413 => to_unsigned(29032, LUT_AMPL_WIDTH - 1),
		21414 => to_unsigned(29030, LUT_AMPL_WIDTH - 1),
		21415 => to_unsigned(29029, LUT_AMPL_WIDTH - 1),
		21416 => to_unsigned(29027, LUT_AMPL_WIDTH - 1),
		21417 => to_unsigned(29026, LUT_AMPL_WIDTH - 1),
		21418 => to_unsigned(29024, LUT_AMPL_WIDTH - 1),
		21419 => to_unsigned(29023, LUT_AMPL_WIDTH - 1),
		21420 => to_unsigned(29021, LUT_AMPL_WIDTH - 1),
		21421 => to_unsigned(29020, LUT_AMPL_WIDTH - 1),
		21422 => to_unsigned(29018, LUT_AMPL_WIDTH - 1),
		21423 => to_unsigned(29017, LUT_AMPL_WIDTH - 1),
		21424 => to_unsigned(29016, LUT_AMPL_WIDTH - 1),
		21425 => to_unsigned(29014, LUT_AMPL_WIDTH - 1),
		21426 => to_unsigned(29013, LUT_AMPL_WIDTH - 1),
		21427 => to_unsigned(29011, LUT_AMPL_WIDTH - 1),
		21428 => to_unsigned(29010, LUT_AMPL_WIDTH - 1),
		21429 => to_unsigned(29008, LUT_AMPL_WIDTH - 1),
		21430 => to_unsigned(29007, LUT_AMPL_WIDTH - 1),
		21431 => to_unsigned(29005, LUT_AMPL_WIDTH - 1),
		21432 => to_unsigned(29004, LUT_AMPL_WIDTH - 1),
		21433 => to_unsigned(29002, LUT_AMPL_WIDTH - 1),
		21434 => to_unsigned(29001, LUT_AMPL_WIDTH - 1),
		21435 => to_unsigned(28999, LUT_AMPL_WIDTH - 1),
		21436 => to_unsigned(28998, LUT_AMPL_WIDTH - 1),
		21437 => to_unsigned(28997, LUT_AMPL_WIDTH - 1),
		21438 => to_unsigned(28995, LUT_AMPL_WIDTH - 1),
		21439 => to_unsigned(28994, LUT_AMPL_WIDTH - 1),
		21440 => to_unsigned(28992, LUT_AMPL_WIDTH - 1),
		21441 => to_unsigned(28991, LUT_AMPL_WIDTH - 1),
		21442 => to_unsigned(28989, LUT_AMPL_WIDTH - 1),
		21443 => to_unsigned(28988, LUT_AMPL_WIDTH - 1),
		21444 => to_unsigned(28986, LUT_AMPL_WIDTH - 1),
		21445 => to_unsigned(28985, LUT_AMPL_WIDTH - 1),
		21446 => to_unsigned(28983, LUT_AMPL_WIDTH - 1),
		21447 => to_unsigned(28982, LUT_AMPL_WIDTH - 1),
		21448 => to_unsigned(28980, LUT_AMPL_WIDTH - 1),
		21449 => to_unsigned(28979, LUT_AMPL_WIDTH - 1),
		21450 => to_unsigned(28977, LUT_AMPL_WIDTH - 1),
		21451 => to_unsigned(28976, LUT_AMPL_WIDTH - 1),
		21452 => to_unsigned(28975, LUT_AMPL_WIDTH - 1),
		21453 => to_unsigned(28973, LUT_AMPL_WIDTH - 1),
		21454 => to_unsigned(28972, LUT_AMPL_WIDTH - 1),
		21455 => to_unsigned(28970, LUT_AMPL_WIDTH - 1),
		21456 => to_unsigned(28969, LUT_AMPL_WIDTH - 1),
		21457 => to_unsigned(28967, LUT_AMPL_WIDTH - 1),
		21458 => to_unsigned(28966, LUT_AMPL_WIDTH - 1),
		21459 => to_unsigned(28964, LUT_AMPL_WIDTH - 1),
		21460 => to_unsigned(28963, LUT_AMPL_WIDTH - 1),
		21461 => to_unsigned(28961, LUT_AMPL_WIDTH - 1),
		21462 => to_unsigned(28960, LUT_AMPL_WIDTH - 1),
		21463 => to_unsigned(28958, LUT_AMPL_WIDTH - 1),
		21464 => to_unsigned(28957, LUT_AMPL_WIDTH - 1),
		21465 => to_unsigned(28955, LUT_AMPL_WIDTH - 1),
		21466 => to_unsigned(28954, LUT_AMPL_WIDTH - 1),
		21467 => to_unsigned(28953, LUT_AMPL_WIDTH - 1),
		21468 => to_unsigned(28951, LUT_AMPL_WIDTH - 1),
		21469 => to_unsigned(28950, LUT_AMPL_WIDTH - 1),
		21470 => to_unsigned(28948, LUT_AMPL_WIDTH - 1),
		21471 => to_unsigned(28947, LUT_AMPL_WIDTH - 1),
		21472 => to_unsigned(28945, LUT_AMPL_WIDTH - 1),
		21473 => to_unsigned(28944, LUT_AMPL_WIDTH - 1),
		21474 => to_unsigned(28942, LUT_AMPL_WIDTH - 1),
		21475 => to_unsigned(28941, LUT_AMPL_WIDTH - 1),
		21476 => to_unsigned(28939, LUT_AMPL_WIDTH - 1),
		21477 => to_unsigned(28938, LUT_AMPL_WIDTH - 1),
		21478 => to_unsigned(28936, LUT_AMPL_WIDTH - 1),
		21479 => to_unsigned(28935, LUT_AMPL_WIDTH - 1),
		21480 => to_unsigned(28933, LUT_AMPL_WIDTH - 1),
		21481 => to_unsigned(28932, LUT_AMPL_WIDTH - 1),
		21482 => to_unsigned(28930, LUT_AMPL_WIDTH - 1),
		21483 => to_unsigned(28929, LUT_AMPL_WIDTH - 1),
		21484 => to_unsigned(28927, LUT_AMPL_WIDTH - 1),
		21485 => to_unsigned(28926, LUT_AMPL_WIDTH - 1),
		21486 => to_unsigned(28925, LUT_AMPL_WIDTH - 1),
		21487 => to_unsigned(28923, LUT_AMPL_WIDTH - 1),
		21488 => to_unsigned(28922, LUT_AMPL_WIDTH - 1),
		21489 => to_unsigned(28920, LUT_AMPL_WIDTH - 1),
		21490 => to_unsigned(28919, LUT_AMPL_WIDTH - 1),
		21491 => to_unsigned(28917, LUT_AMPL_WIDTH - 1),
		21492 => to_unsigned(28916, LUT_AMPL_WIDTH - 1),
		21493 => to_unsigned(28914, LUT_AMPL_WIDTH - 1),
		21494 => to_unsigned(28913, LUT_AMPL_WIDTH - 1),
		21495 => to_unsigned(28911, LUT_AMPL_WIDTH - 1),
		21496 => to_unsigned(28910, LUT_AMPL_WIDTH - 1),
		21497 => to_unsigned(28908, LUT_AMPL_WIDTH - 1),
		21498 => to_unsigned(28907, LUT_AMPL_WIDTH - 1),
		21499 => to_unsigned(28905, LUT_AMPL_WIDTH - 1),
		21500 => to_unsigned(28904, LUT_AMPL_WIDTH - 1),
		21501 => to_unsigned(28902, LUT_AMPL_WIDTH - 1),
		21502 => to_unsigned(28901, LUT_AMPL_WIDTH - 1),
		21503 => to_unsigned(28899, LUT_AMPL_WIDTH - 1),
		21504 => to_unsigned(28898, LUT_AMPL_WIDTH - 1),
		21505 => to_unsigned(28896, LUT_AMPL_WIDTH - 1),
		21506 => to_unsigned(28895, LUT_AMPL_WIDTH - 1),
		21507 => to_unsigned(28893, LUT_AMPL_WIDTH - 1),
		21508 => to_unsigned(28892, LUT_AMPL_WIDTH - 1),
		21509 => to_unsigned(28891, LUT_AMPL_WIDTH - 1),
		21510 => to_unsigned(28889, LUT_AMPL_WIDTH - 1),
		21511 => to_unsigned(28888, LUT_AMPL_WIDTH - 1),
		21512 => to_unsigned(28886, LUT_AMPL_WIDTH - 1),
		21513 => to_unsigned(28885, LUT_AMPL_WIDTH - 1),
		21514 => to_unsigned(28883, LUT_AMPL_WIDTH - 1),
		21515 => to_unsigned(28882, LUT_AMPL_WIDTH - 1),
		21516 => to_unsigned(28880, LUT_AMPL_WIDTH - 1),
		21517 => to_unsigned(28879, LUT_AMPL_WIDTH - 1),
		21518 => to_unsigned(28877, LUT_AMPL_WIDTH - 1),
		21519 => to_unsigned(28876, LUT_AMPL_WIDTH - 1),
		21520 => to_unsigned(28874, LUT_AMPL_WIDTH - 1),
		21521 => to_unsigned(28873, LUT_AMPL_WIDTH - 1),
		21522 => to_unsigned(28871, LUT_AMPL_WIDTH - 1),
		21523 => to_unsigned(28870, LUT_AMPL_WIDTH - 1),
		21524 => to_unsigned(28868, LUT_AMPL_WIDTH - 1),
		21525 => to_unsigned(28867, LUT_AMPL_WIDTH - 1),
		21526 => to_unsigned(28865, LUT_AMPL_WIDTH - 1),
		21527 => to_unsigned(28864, LUT_AMPL_WIDTH - 1),
		21528 => to_unsigned(28862, LUT_AMPL_WIDTH - 1),
		21529 => to_unsigned(28861, LUT_AMPL_WIDTH - 1),
		21530 => to_unsigned(28859, LUT_AMPL_WIDTH - 1),
		21531 => to_unsigned(28858, LUT_AMPL_WIDTH - 1),
		21532 => to_unsigned(28856, LUT_AMPL_WIDTH - 1),
		21533 => to_unsigned(28855, LUT_AMPL_WIDTH - 1),
		21534 => to_unsigned(28853, LUT_AMPL_WIDTH - 1),
		21535 => to_unsigned(28852, LUT_AMPL_WIDTH - 1),
		21536 => to_unsigned(28850, LUT_AMPL_WIDTH - 1),
		21537 => to_unsigned(28849, LUT_AMPL_WIDTH - 1),
		21538 => to_unsigned(28847, LUT_AMPL_WIDTH - 1),
		21539 => to_unsigned(28846, LUT_AMPL_WIDTH - 1),
		21540 => to_unsigned(28844, LUT_AMPL_WIDTH - 1),
		21541 => to_unsigned(28843, LUT_AMPL_WIDTH - 1),
		21542 => to_unsigned(28841, LUT_AMPL_WIDTH - 1),
		21543 => to_unsigned(28840, LUT_AMPL_WIDTH - 1),
		21544 => to_unsigned(28838, LUT_AMPL_WIDTH - 1),
		21545 => to_unsigned(28837, LUT_AMPL_WIDTH - 1),
		21546 => to_unsigned(28835, LUT_AMPL_WIDTH - 1),
		21547 => to_unsigned(28834, LUT_AMPL_WIDTH - 1),
		21548 => to_unsigned(28832, LUT_AMPL_WIDTH - 1),
		21549 => to_unsigned(28831, LUT_AMPL_WIDTH - 1),
		21550 => to_unsigned(28830, LUT_AMPL_WIDTH - 1),
		21551 => to_unsigned(28828, LUT_AMPL_WIDTH - 1),
		21552 => to_unsigned(28827, LUT_AMPL_WIDTH - 1),
		21553 => to_unsigned(28825, LUT_AMPL_WIDTH - 1),
		21554 => to_unsigned(28824, LUT_AMPL_WIDTH - 1),
		21555 => to_unsigned(28822, LUT_AMPL_WIDTH - 1),
		21556 => to_unsigned(28821, LUT_AMPL_WIDTH - 1),
		21557 => to_unsigned(28819, LUT_AMPL_WIDTH - 1),
		21558 => to_unsigned(28818, LUT_AMPL_WIDTH - 1),
		21559 => to_unsigned(28816, LUT_AMPL_WIDTH - 1),
		21560 => to_unsigned(28815, LUT_AMPL_WIDTH - 1),
		21561 => to_unsigned(28813, LUT_AMPL_WIDTH - 1),
		21562 => to_unsigned(28812, LUT_AMPL_WIDTH - 1),
		21563 => to_unsigned(28810, LUT_AMPL_WIDTH - 1),
		21564 => to_unsigned(28809, LUT_AMPL_WIDTH - 1),
		21565 => to_unsigned(28807, LUT_AMPL_WIDTH - 1),
		21566 => to_unsigned(28806, LUT_AMPL_WIDTH - 1),
		21567 => to_unsigned(28804, LUT_AMPL_WIDTH - 1),
		21568 => to_unsigned(28803, LUT_AMPL_WIDTH - 1),
		21569 => to_unsigned(28801, LUT_AMPL_WIDTH - 1),
		21570 => to_unsigned(28800, LUT_AMPL_WIDTH - 1),
		21571 => to_unsigned(28798, LUT_AMPL_WIDTH - 1),
		21572 => to_unsigned(28797, LUT_AMPL_WIDTH - 1),
		21573 => to_unsigned(28795, LUT_AMPL_WIDTH - 1),
		21574 => to_unsigned(28794, LUT_AMPL_WIDTH - 1),
		21575 => to_unsigned(28792, LUT_AMPL_WIDTH - 1),
		21576 => to_unsigned(28791, LUT_AMPL_WIDTH - 1),
		21577 => to_unsigned(28789, LUT_AMPL_WIDTH - 1),
		21578 => to_unsigned(28788, LUT_AMPL_WIDTH - 1),
		21579 => to_unsigned(28786, LUT_AMPL_WIDTH - 1),
		21580 => to_unsigned(28785, LUT_AMPL_WIDTH - 1),
		21581 => to_unsigned(28783, LUT_AMPL_WIDTH - 1),
		21582 => to_unsigned(28782, LUT_AMPL_WIDTH - 1),
		21583 => to_unsigned(28780, LUT_AMPL_WIDTH - 1),
		21584 => to_unsigned(28779, LUT_AMPL_WIDTH - 1),
		21585 => to_unsigned(28777, LUT_AMPL_WIDTH - 1),
		21586 => to_unsigned(28776, LUT_AMPL_WIDTH - 1),
		21587 => to_unsigned(28774, LUT_AMPL_WIDTH - 1),
		21588 => to_unsigned(28773, LUT_AMPL_WIDTH - 1),
		21589 => to_unsigned(28771, LUT_AMPL_WIDTH - 1),
		21590 => to_unsigned(28770, LUT_AMPL_WIDTH - 1),
		21591 => to_unsigned(28768, LUT_AMPL_WIDTH - 1),
		21592 => to_unsigned(28767, LUT_AMPL_WIDTH - 1),
		21593 => to_unsigned(28765, LUT_AMPL_WIDTH - 1),
		21594 => to_unsigned(28764, LUT_AMPL_WIDTH - 1),
		21595 => to_unsigned(28762, LUT_AMPL_WIDTH - 1),
		21596 => to_unsigned(28761, LUT_AMPL_WIDTH - 1),
		21597 => to_unsigned(28759, LUT_AMPL_WIDTH - 1),
		21598 => to_unsigned(28758, LUT_AMPL_WIDTH - 1),
		21599 => to_unsigned(28756, LUT_AMPL_WIDTH - 1),
		21600 => to_unsigned(28755, LUT_AMPL_WIDTH - 1),
		21601 => to_unsigned(28753, LUT_AMPL_WIDTH - 1),
		21602 => to_unsigned(28752, LUT_AMPL_WIDTH - 1),
		21603 => to_unsigned(28750, LUT_AMPL_WIDTH - 1),
		21604 => to_unsigned(28748, LUT_AMPL_WIDTH - 1),
		21605 => to_unsigned(28747, LUT_AMPL_WIDTH - 1),
		21606 => to_unsigned(28745, LUT_AMPL_WIDTH - 1),
		21607 => to_unsigned(28744, LUT_AMPL_WIDTH - 1),
		21608 => to_unsigned(28742, LUT_AMPL_WIDTH - 1),
		21609 => to_unsigned(28741, LUT_AMPL_WIDTH - 1),
		21610 => to_unsigned(28739, LUT_AMPL_WIDTH - 1),
		21611 => to_unsigned(28738, LUT_AMPL_WIDTH - 1),
		21612 => to_unsigned(28736, LUT_AMPL_WIDTH - 1),
		21613 => to_unsigned(28735, LUT_AMPL_WIDTH - 1),
		21614 => to_unsigned(28733, LUT_AMPL_WIDTH - 1),
		21615 => to_unsigned(28732, LUT_AMPL_WIDTH - 1),
		21616 => to_unsigned(28730, LUT_AMPL_WIDTH - 1),
		21617 => to_unsigned(28729, LUT_AMPL_WIDTH - 1),
		21618 => to_unsigned(28727, LUT_AMPL_WIDTH - 1),
		21619 => to_unsigned(28726, LUT_AMPL_WIDTH - 1),
		21620 => to_unsigned(28724, LUT_AMPL_WIDTH - 1),
		21621 => to_unsigned(28723, LUT_AMPL_WIDTH - 1),
		21622 => to_unsigned(28721, LUT_AMPL_WIDTH - 1),
		21623 => to_unsigned(28720, LUT_AMPL_WIDTH - 1),
		21624 => to_unsigned(28718, LUT_AMPL_WIDTH - 1),
		21625 => to_unsigned(28717, LUT_AMPL_WIDTH - 1),
		21626 => to_unsigned(28715, LUT_AMPL_WIDTH - 1),
		21627 => to_unsigned(28714, LUT_AMPL_WIDTH - 1),
		21628 => to_unsigned(28712, LUT_AMPL_WIDTH - 1),
		21629 => to_unsigned(28711, LUT_AMPL_WIDTH - 1),
		21630 => to_unsigned(28709, LUT_AMPL_WIDTH - 1),
		21631 => to_unsigned(28708, LUT_AMPL_WIDTH - 1),
		21632 => to_unsigned(28706, LUT_AMPL_WIDTH - 1),
		21633 => to_unsigned(28705, LUT_AMPL_WIDTH - 1),
		21634 => to_unsigned(28703, LUT_AMPL_WIDTH - 1),
		21635 => to_unsigned(28702, LUT_AMPL_WIDTH - 1),
		21636 => to_unsigned(28700, LUT_AMPL_WIDTH - 1),
		21637 => to_unsigned(28699, LUT_AMPL_WIDTH - 1),
		21638 => to_unsigned(28697, LUT_AMPL_WIDTH - 1),
		21639 => to_unsigned(28696, LUT_AMPL_WIDTH - 1),
		21640 => to_unsigned(28694, LUT_AMPL_WIDTH - 1),
		21641 => to_unsigned(28693, LUT_AMPL_WIDTH - 1),
		21642 => to_unsigned(28691, LUT_AMPL_WIDTH - 1),
		21643 => to_unsigned(28690, LUT_AMPL_WIDTH - 1),
		21644 => to_unsigned(28688, LUT_AMPL_WIDTH - 1),
		21645 => to_unsigned(28686, LUT_AMPL_WIDTH - 1),
		21646 => to_unsigned(28685, LUT_AMPL_WIDTH - 1),
		21647 => to_unsigned(28683, LUT_AMPL_WIDTH - 1),
		21648 => to_unsigned(28682, LUT_AMPL_WIDTH - 1),
		21649 => to_unsigned(28680, LUT_AMPL_WIDTH - 1),
		21650 => to_unsigned(28679, LUT_AMPL_WIDTH - 1),
		21651 => to_unsigned(28677, LUT_AMPL_WIDTH - 1),
		21652 => to_unsigned(28676, LUT_AMPL_WIDTH - 1),
		21653 => to_unsigned(28674, LUT_AMPL_WIDTH - 1),
		21654 => to_unsigned(28673, LUT_AMPL_WIDTH - 1),
		21655 => to_unsigned(28671, LUT_AMPL_WIDTH - 1),
		21656 => to_unsigned(28670, LUT_AMPL_WIDTH - 1),
		21657 => to_unsigned(28668, LUT_AMPL_WIDTH - 1),
		21658 => to_unsigned(28667, LUT_AMPL_WIDTH - 1),
		21659 => to_unsigned(28665, LUT_AMPL_WIDTH - 1),
		21660 => to_unsigned(28664, LUT_AMPL_WIDTH - 1),
		21661 => to_unsigned(28662, LUT_AMPL_WIDTH - 1),
		21662 => to_unsigned(28661, LUT_AMPL_WIDTH - 1),
		21663 => to_unsigned(28659, LUT_AMPL_WIDTH - 1),
		21664 => to_unsigned(28658, LUT_AMPL_WIDTH - 1),
		21665 => to_unsigned(28656, LUT_AMPL_WIDTH - 1),
		21666 => to_unsigned(28655, LUT_AMPL_WIDTH - 1),
		21667 => to_unsigned(28653, LUT_AMPL_WIDTH - 1),
		21668 => to_unsigned(28651, LUT_AMPL_WIDTH - 1),
		21669 => to_unsigned(28650, LUT_AMPL_WIDTH - 1),
		21670 => to_unsigned(28648, LUT_AMPL_WIDTH - 1),
		21671 => to_unsigned(28647, LUT_AMPL_WIDTH - 1),
		21672 => to_unsigned(28645, LUT_AMPL_WIDTH - 1),
		21673 => to_unsigned(28644, LUT_AMPL_WIDTH - 1),
		21674 => to_unsigned(28642, LUT_AMPL_WIDTH - 1),
		21675 => to_unsigned(28641, LUT_AMPL_WIDTH - 1),
		21676 => to_unsigned(28639, LUT_AMPL_WIDTH - 1),
		21677 => to_unsigned(28638, LUT_AMPL_WIDTH - 1),
		21678 => to_unsigned(28636, LUT_AMPL_WIDTH - 1),
		21679 => to_unsigned(28635, LUT_AMPL_WIDTH - 1),
		21680 => to_unsigned(28633, LUT_AMPL_WIDTH - 1),
		21681 => to_unsigned(28632, LUT_AMPL_WIDTH - 1),
		21682 => to_unsigned(28630, LUT_AMPL_WIDTH - 1),
		21683 => to_unsigned(28629, LUT_AMPL_WIDTH - 1),
		21684 => to_unsigned(28627, LUT_AMPL_WIDTH - 1),
		21685 => to_unsigned(28626, LUT_AMPL_WIDTH - 1),
		21686 => to_unsigned(28624, LUT_AMPL_WIDTH - 1),
		21687 => to_unsigned(28622, LUT_AMPL_WIDTH - 1),
		21688 => to_unsigned(28621, LUT_AMPL_WIDTH - 1),
		21689 => to_unsigned(28619, LUT_AMPL_WIDTH - 1),
		21690 => to_unsigned(28618, LUT_AMPL_WIDTH - 1),
		21691 => to_unsigned(28616, LUT_AMPL_WIDTH - 1),
		21692 => to_unsigned(28615, LUT_AMPL_WIDTH - 1),
		21693 => to_unsigned(28613, LUT_AMPL_WIDTH - 1),
		21694 => to_unsigned(28612, LUT_AMPL_WIDTH - 1),
		21695 => to_unsigned(28610, LUT_AMPL_WIDTH - 1),
		21696 => to_unsigned(28609, LUT_AMPL_WIDTH - 1),
		21697 => to_unsigned(28607, LUT_AMPL_WIDTH - 1),
		21698 => to_unsigned(28606, LUT_AMPL_WIDTH - 1),
		21699 => to_unsigned(28604, LUT_AMPL_WIDTH - 1),
		21700 => to_unsigned(28603, LUT_AMPL_WIDTH - 1),
		21701 => to_unsigned(28601, LUT_AMPL_WIDTH - 1),
		21702 => to_unsigned(28600, LUT_AMPL_WIDTH - 1),
		21703 => to_unsigned(28598, LUT_AMPL_WIDTH - 1),
		21704 => to_unsigned(28596, LUT_AMPL_WIDTH - 1),
		21705 => to_unsigned(28595, LUT_AMPL_WIDTH - 1),
		21706 => to_unsigned(28593, LUT_AMPL_WIDTH - 1),
		21707 => to_unsigned(28592, LUT_AMPL_WIDTH - 1),
		21708 => to_unsigned(28590, LUT_AMPL_WIDTH - 1),
		21709 => to_unsigned(28589, LUT_AMPL_WIDTH - 1),
		21710 => to_unsigned(28587, LUT_AMPL_WIDTH - 1),
		21711 => to_unsigned(28586, LUT_AMPL_WIDTH - 1),
		21712 => to_unsigned(28584, LUT_AMPL_WIDTH - 1),
		21713 => to_unsigned(28583, LUT_AMPL_WIDTH - 1),
		21714 => to_unsigned(28581, LUT_AMPL_WIDTH - 1),
		21715 => to_unsigned(28580, LUT_AMPL_WIDTH - 1),
		21716 => to_unsigned(28578, LUT_AMPL_WIDTH - 1),
		21717 => to_unsigned(28576, LUT_AMPL_WIDTH - 1),
		21718 => to_unsigned(28575, LUT_AMPL_WIDTH - 1),
		21719 => to_unsigned(28573, LUT_AMPL_WIDTH - 1),
		21720 => to_unsigned(28572, LUT_AMPL_WIDTH - 1),
		21721 => to_unsigned(28570, LUT_AMPL_WIDTH - 1),
		21722 => to_unsigned(28569, LUT_AMPL_WIDTH - 1),
		21723 => to_unsigned(28567, LUT_AMPL_WIDTH - 1),
		21724 => to_unsigned(28566, LUT_AMPL_WIDTH - 1),
		21725 => to_unsigned(28564, LUT_AMPL_WIDTH - 1),
		21726 => to_unsigned(28563, LUT_AMPL_WIDTH - 1),
		21727 => to_unsigned(28561, LUT_AMPL_WIDTH - 1),
		21728 => to_unsigned(28560, LUT_AMPL_WIDTH - 1),
		21729 => to_unsigned(28558, LUT_AMPL_WIDTH - 1),
		21730 => to_unsigned(28556, LUT_AMPL_WIDTH - 1),
		21731 => to_unsigned(28555, LUT_AMPL_WIDTH - 1),
		21732 => to_unsigned(28553, LUT_AMPL_WIDTH - 1),
		21733 => to_unsigned(28552, LUT_AMPL_WIDTH - 1),
		21734 => to_unsigned(28550, LUT_AMPL_WIDTH - 1),
		21735 => to_unsigned(28549, LUT_AMPL_WIDTH - 1),
		21736 => to_unsigned(28547, LUT_AMPL_WIDTH - 1),
		21737 => to_unsigned(28546, LUT_AMPL_WIDTH - 1),
		21738 => to_unsigned(28544, LUT_AMPL_WIDTH - 1),
		21739 => to_unsigned(28543, LUT_AMPL_WIDTH - 1),
		21740 => to_unsigned(28541, LUT_AMPL_WIDTH - 1),
		21741 => to_unsigned(28540, LUT_AMPL_WIDTH - 1),
		21742 => to_unsigned(28538, LUT_AMPL_WIDTH - 1),
		21743 => to_unsigned(28536, LUT_AMPL_WIDTH - 1),
		21744 => to_unsigned(28535, LUT_AMPL_WIDTH - 1),
		21745 => to_unsigned(28533, LUT_AMPL_WIDTH - 1),
		21746 => to_unsigned(28532, LUT_AMPL_WIDTH - 1),
		21747 => to_unsigned(28530, LUT_AMPL_WIDTH - 1),
		21748 => to_unsigned(28529, LUT_AMPL_WIDTH - 1),
		21749 => to_unsigned(28527, LUT_AMPL_WIDTH - 1),
		21750 => to_unsigned(28526, LUT_AMPL_WIDTH - 1),
		21751 => to_unsigned(28524, LUT_AMPL_WIDTH - 1),
		21752 => to_unsigned(28523, LUT_AMPL_WIDTH - 1),
		21753 => to_unsigned(28521, LUT_AMPL_WIDTH - 1),
		21754 => to_unsigned(28519, LUT_AMPL_WIDTH - 1),
		21755 => to_unsigned(28518, LUT_AMPL_WIDTH - 1),
		21756 => to_unsigned(28516, LUT_AMPL_WIDTH - 1),
		21757 => to_unsigned(28515, LUT_AMPL_WIDTH - 1),
		21758 => to_unsigned(28513, LUT_AMPL_WIDTH - 1),
		21759 => to_unsigned(28512, LUT_AMPL_WIDTH - 1),
		21760 => to_unsigned(28510, LUT_AMPL_WIDTH - 1),
		21761 => to_unsigned(28509, LUT_AMPL_WIDTH - 1),
		21762 => to_unsigned(28507, LUT_AMPL_WIDTH - 1),
		21763 => to_unsigned(28505, LUT_AMPL_WIDTH - 1),
		21764 => to_unsigned(28504, LUT_AMPL_WIDTH - 1),
		21765 => to_unsigned(28502, LUT_AMPL_WIDTH - 1),
		21766 => to_unsigned(28501, LUT_AMPL_WIDTH - 1),
		21767 => to_unsigned(28499, LUT_AMPL_WIDTH - 1),
		21768 => to_unsigned(28498, LUT_AMPL_WIDTH - 1),
		21769 => to_unsigned(28496, LUT_AMPL_WIDTH - 1),
		21770 => to_unsigned(28495, LUT_AMPL_WIDTH - 1),
		21771 => to_unsigned(28493, LUT_AMPL_WIDTH - 1),
		21772 => to_unsigned(28492, LUT_AMPL_WIDTH - 1),
		21773 => to_unsigned(28490, LUT_AMPL_WIDTH - 1),
		21774 => to_unsigned(28488, LUT_AMPL_WIDTH - 1),
		21775 => to_unsigned(28487, LUT_AMPL_WIDTH - 1),
		21776 => to_unsigned(28485, LUT_AMPL_WIDTH - 1),
		21777 => to_unsigned(28484, LUT_AMPL_WIDTH - 1),
		21778 => to_unsigned(28482, LUT_AMPL_WIDTH - 1),
		21779 => to_unsigned(28481, LUT_AMPL_WIDTH - 1),
		21780 => to_unsigned(28479, LUT_AMPL_WIDTH - 1),
		21781 => to_unsigned(28478, LUT_AMPL_WIDTH - 1),
		21782 => to_unsigned(28476, LUT_AMPL_WIDTH - 1),
		21783 => to_unsigned(28474, LUT_AMPL_WIDTH - 1),
		21784 => to_unsigned(28473, LUT_AMPL_WIDTH - 1),
		21785 => to_unsigned(28471, LUT_AMPL_WIDTH - 1),
		21786 => to_unsigned(28470, LUT_AMPL_WIDTH - 1),
		21787 => to_unsigned(28468, LUT_AMPL_WIDTH - 1),
		21788 => to_unsigned(28467, LUT_AMPL_WIDTH - 1),
		21789 => to_unsigned(28465, LUT_AMPL_WIDTH - 1),
		21790 => to_unsigned(28464, LUT_AMPL_WIDTH - 1),
		21791 => to_unsigned(28462, LUT_AMPL_WIDTH - 1),
		21792 => to_unsigned(28460, LUT_AMPL_WIDTH - 1),
		21793 => to_unsigned(28459, LUT_AMPL_WIDTH - 1),
		21794 => to_unsigned(28457, LUT_AMPL_WIDTH - 1),
		21795 => to_unsigned(28456, LUT_AMPL_WIDTH - 1),
		21796 => to_unsigned(28454, LUT_AMPL_WIDTH - 1),
		21797 => to_unsigned(28453, LUT_AMPL_WIDTH - 1),
		21798 => to_unsigned(28451, LUT_AMPL_WIDTH - 1),
		21799 => to_unsigned(28450, LUT_AMPL_WIDTH - 1),
		21800 => to_unsigned(28448, LUT_AMPL_WIDTH - 1),
		21801 => to_unsigned(28446, LUT_AMPL_WIDTH - 1),
		21802 => to_unsigned(28445, LUT_AMPL_WIDTH - 1),
		21803 => to_unsigned(28443, LUT_AMPL_WIDTH - 1),
		21804 => to_unsigned(28442, LUT_AMPL_WIDTH - 1),
		21805 => to_unsigned(28440, LUT_AMPL_WIDTH - 1),
		21806 => to_unsigned(28439, LUT_AMPL_WIDTH - 1),
		21807 => to_unsigned(28437, LUT_AMPL_WIDTH - 1),
		21808 => to_unsigned(28436, LUT_AMPL_WIDTH - 1),
		21809 => to_unsigned(28434, LUT_AMPL_WIDTH - 1),
		21810 => to_unsigned(28432, LUT_AMPL_WIDTH - 1),
		21811 => to_unsigned(28431, LUT_AMPL_WIDTH - 1),
		21812 => to_unsigned(28429, LUT_AMPL_WIDTH - 1),
		21813 => to_unsigned(28428, LUT_AMPL_WIDTH - 1),
		21814 => to_unsigned(28426, LUT_AMPL_WIDTH - 1),
		21815 => to_unsigned(28425, LUT_AMPL_WIDTH - 1),
		21816 => to_unsigned(28423, LUT_AMPL_WIDTH - 1),
		21817 => to_unsigned(28421, LUT_AMPL_WIDTH - 1),
		21818 => to_unsigned(28420, LUT_AMPL_WIDTH - 1),
		21819 => to_unsigned(28418, LUT_AMPL_WIDTH - 1),
		21820 => to_unsigned(28417, LUT_AMPL_WIDTH - 1),
		21821 => to_unsigned(28415, LUT_AMPL_WIDTH - 1),
		21822 => to_unsigned(28414, LUT_AMPL_WIDTH - 1),
		21823 => to_unsigned(28412, LUT_AMPL_WIDTH - 1),
		21824 => to_unsigned(28411, LUT_AMPL_WIDTH - 1),
		21825 => to_unsigned(28409, LUT_AMPL_WIDTH - 1),
		21826 => to_unsigned(28407, LUT_AMPL_WIDTH - 1),
		21827 => to_unsigned(28406, LUT_AMPL_WIDTH - 1),
		21828 => to_unsigned(28404, LUT_AMPL_WIDTH - 1),
		21829 => to_unsigned(28403, LUT_AMPL_WIDTH - 1),
		21830 => to_unsigned(28401, LUT_AMPL_WIDTH - 1),
		21831 => to_unsigned(28400, LUT_AMPL_WIDTH - 1),
		21832 => to_unsigned(28398, LUT_AMPL_WIDTH - 1),
		21833 => to_unsigned(28396, LUT_AMPL_WIDTH - 1),
		21834 => to_unsigned(28395, LUT_AMPL_WIDTH - 1),
		21835 => to_unsigned(28393, LUT_AMPL_WIDTH - 1),
		21836 => to_unsigned(28392, LUT_AMPL_WIDTH - 1),
		21837 => to_unsigned(28390, LUT_AMPL_WIDTH - 1),
		21838 => to_unsigned(28389, LUT_AMPL_WIDTH - 1),
		21839 => to_unsigned(28387, LUT_AMPL_WIDTH - 1),
		21840 => to_unsigned(28385, LUT_AMPL_WIDTH - 1),
		21841 => to_unsigned(28384, LUT_AMPL_WIDTH - 1),
		21842 => to_unsigned(28382, LUT_AMPL_WIDTH - 1),
		21843 => to_unsigned(28381, LUT_AMPL_WIDTH - 1),
		21844 => to_unsigned(28379, LUT_AMPL_WIDTH - 1),
		21845 => to_unsigned(28378, LUT_AMPL_WIDTH - 1),
		21846 => to_unsigned(28376, LUT_AMPL_WIDTH - 1),
		21847 => to_unsigned(28374, LUT_AMPL_WIDTH - 1),
		21848 => to_unsigned(28373, LUT_AMPL_WIDTH - 1),
		21849 => to_unsigned(28371, LUT_AMPL_WIDTH - 1),
		21850 => to_unsigned(28370, LUT_AMPL_WIDTH - 1),
		21851 => to_unsigned(28368, LUT_AMPL_WIDTH - 1),
		21852 => to_unsigned(28367, LUT_AMPL_WIDTH - 1),
		21853 => to_unsigned(28365, LUT_AMPL_WIDTH - 1),
		21854 => to_unsigned(28363, LUT_AMPL_WIDTH - 1),
		21855 => to_unsigned(28362, LUT_AMPL_WIDTH - 1),
		21856 => to_unsigned(28360, LUT_AMPL_WIDTH - 1),
		21857 => to_unsigned(28359, LUT_AMPL_WIDTH - 1),
		21858 => to_unsigned(28357, LUT_AMPL_WIDTH - 1),
		21859 => to_unsigned(28356, LUT_AMPL_WIDTH - 1),
		21860 => to_unsigned(28354, LUT_AMPL_WIDTH - 1),
		21861 => to_unsigned(28352, LUT_AMPL_WIDTH - 1),
		21862 => to_unsigned(28351, LUT_AMPL_WIDTH - 1),
		21863 => to_unsigned(28349, LUT_AMPL_WIDTH - 1),
		21864 => to_unsigned(28348, LUT_AMPL_WIDTH - 1),
		21865 => to_unsigned(28346, LUT_AMPL_WIDTH - 1),
		21866 => to_unsigned(28345, LUT_AMPL_WIDTH - 1),
		21867 => to_unsigned(28343, LUT_AMPL_WIDTH - 1),
		21868 => to_unsigned(28341, LUT_AMPL_WIDTH - 1),
		21869 => to_unsigned(28340, LUT_AMPL_WIDTH - 1),
		21870 => to_unsigned(28338, LUT_AMPL_WIDTH - 1),
		21871 => to_unsigned(28337, LUT_AMPL_WIDTH - 1),
		21872 => to_unsigned(28335, LUT_AMPL_WIDTH - 1),
		21873 => to_unsigned(28333, LUT_AMPL_WIDTH - 1),
		21874 => to_unsigned(28332, LUT_AMPL_WIDTH - 1),
		21875 => to_unsigned(28330, LUT_AMPL_WIDTH - 1),
		21876 => to_unsigned(28329, LUT_AMPL_WIDTH - 1),
		21877 => to_unsigned(28327, LUT_AMPL_WIDTH - 1),
		21878 => to_unsigned(28326, LUT_AMPL_WIDTH - 1),
		21879 => to_unsigned(28324, LUT_AMPL_WIDTH - 1),
		21880 => to_unsigned(28322, LUT_AMPL_WIDTH - 1),
		21881 => to_unsigned(28321, LUT_AMPL_WIDTH - 1),
		21882 => to_unsigned(28319, LUT_AMPL_WIDTH - 1),
		21883 => to_unsigned(28318, LUT_AMPL_WIDTH - 1),
		21884 => to_unsigned(28316, LUT_AMPL_WIDTH - 1),
		21885 => to_unsigned(28315, LUT_AMPL_WIDTH - 1),
		21886 => to_unsigned(28313, LUT_AMPL_WIDTH - 1),
		21887 => to_unsigned(28311, LUT_AMPL_WIDTH - 1),
		21888 => to_unsigned(28310, LUT_AMPL_WIDTH - 1),
		21889 => to_unsigned(28308, LUT_AMPL_WIDTH - 1),
		21890 => to_unsigned(28307, LUT_AMPL_WIDTH - 1),
		21891 => to_unsigned(28305, LUT_AMPL_WIDTH - 1),
		21892 => to_unsigned(28303, LUT_AMPL_WIDTH - 1),
		21893 => to_unsigned(28302, LUT_AMPL_WIDTH - 1),
		21894 => to_unsigned(28300, LUT_AMPL_WIDTH - 1),
		21895 => to_unsigned(28299, LUT_AMPL_WIDTH - 1),
		21896 => to_unsigned(28297, LUT_AMPL_WIDTH - 1),
		21897 => to_unsigned(28296, LUT_AMPL_WIDTH - 1),
		21898 => to_unsigned(28294, LUT_AMPL_WIDTH - 1),
		21899 => to_unsigned(28292, LUT_AMPL_WIDTH - 1),
		21900 => to_unsigned(28291, LUT_AMPL_WIDTH - 1),
		21901 => to_unsigned(28289, LUT_AMPL_WIDTH - 1),
		21902 => to_unsigned(28288, LUT_AMPL_WIDTH - 1),
		21903 => to_unsigned(28286, LUT_AMPL_WIDTH - 1),
		21904 => to_unsigned(28284, LUT_AMPL_WIDTH - 1),
		21905 => to_unsigned(28283, LUT_AMPL_WIDTH - 1),
		21906 => to_unsigned(28281, LUT_AMPL_WIDTH - 1),
		21907 => to_unsigned(28280, LUT_AMPL_WIDTH - 1),
		21908 => to_unsigned(28278, LUT_AMPL_WIDTH - 1),
		21909 => to_unsigned(28277, LUT_AMPL_WIDTH - 1),
		21910 => to_unsigned(28275, LUT_AMPL_WIDTH - 1),
		21911 => to_unsigned(28273, LUT_AMPL_WIDTH - 1),
		21912 => to_unsigned(28272, LUT_AMPL_WIDTH - 1),
		21913 => to_unsigned(28270, LUT_AMPL_WIDTH - 1),
		21914 => to_unsigned(28269, LUT_AMPL_WIDTH - 1),
		21915 => to_unsigned(28267, LUT_AMPL_WIDTH - 1),
		21916 => to_unsigned(28265, LUT_AMPL_WIDTH - 1),
		21917 => to_unsigned(28264, LUT_AMPL_WIDTH - 1),
		21918 => to_unsigned(28262, LUT_AMPL_WIDTH - 1),
		21919 => to_unsigned(28261, LUT_AMPL_WIDTH - 1),
		21920 => to_unsigned(28259, LUT_AMPL_WIDTH - 1),
		21921 => to_unsigned(28257, LUT_AMPL_WIDTH - 1),
		21922 => to_unsigned(28256, LUT_AMPL_WIDTH - 1),
		21923 => to_unsigned(28254, LUT_AMPL_WIDTH - 1),
		21924 => to_unsigned(28253, LUT_AMPL_WIDTH - 1),
		21925 => to_unsigned(28251, LUT_AMPL_WIDTH - 1),
		21926 => to_unsigned(28249, LUT_AMPL_WIDTH - 1),
		21927 => to_unsigned(28248, LUT_AMPL_WIDTH - 1),
		21928 => to_unsigned(28246, LUT_AMPL_WIDTH - 1),
		21929 => to_unsigned(28245, LUT_AMPL_WIDTH - 1),
		21930 => to_unsigned(28243, LUT_AMPL_WIDTH - 1),
		21931 => to_unsigned(28242, LUT_AMPL_WIDTH - 1),
		21932 => to_unsigned(28240, LUT_AMPL_WIDTH - 1),
		21933 => to_unsigned(28238, LUT_AMPL_WIDTH - 1),
		21934 => to_unsigned(28237, LUT_AMPL_WIDTH - 1),
		21935 => to_unsigned(28235, LUT_AMPL_WIDTH - 1),
		21936 => to_unsigned(28234, LUT_AMPL_WIDTH - 1),
		21937 => to_unsigned(28232, LUT_AMPL_WIDTH - 1),
		21938 => to_unsigned(28230, LUT_AMPL_WIDTH - 1),
		21939 => to_unsigned(28229, LUT_AMPL_WIDTH - 1),
		21940 => to_unsigned(28227, LUT_AMPL_WIDTH - 1),
		21941 => to_unsigned(28226, LUT_AMPL_WIDTH - 1),
		21942 => to_unsigned(28224, LUT_AMPL_WIDTH - 1),
		21943 => to_unsigned(28222, LUT_AMPL_WIDTH - 1),
		21944 => to_unsigned(28221, LUT_AMPL_WIDTH - 1),
		21945 => to_unsigned(28219, LUT_AMPL_WIDTH - 1),
		21946 => to_unsigned(28218, LUT_AMPL_WIDTH - 1),
		21947 => to_unsigned(28216, LUT_AMPL_WIDTH - 1),
		21948 => to_unsigned(28214, LUT_AMPL_WIDTH - 1),
		21949 => to_unsigned(28213, LUT_AMPL_WIDTH - 1),
		21950 => to_unsigned(28211, LUT_AMPL_WIDTH - 1),
		21951 => to_unsigned(28210, LUT_AMPL_WIDTH - 1),
		21952 => to_unsigned(28208, LUT_AMPL_WIDTH - 1),
		21953 => to_unsigned(28206, LUT_AMPL_WIDTH - 1),
		21954 => to_unsigned(28205, LUT_AMPL_WIDTH - 1),
		21955 => to_unsigned(28203, LUT_AMPL_WIDTH - 1),
		21956 => to_unsigned(28202, LUT_AMPL_WIDTH - 1),
		21957 => to_unsigned(28200, LUT_AMPL_WIDTH - 1),
		21958 => to_unsigned(28198, LUT_AMPL_WIDTH - 1),
		21959 => to_unsigned(28197, LUT_AMPL_WIDTH - 1),
		21960 => to_unsigned(28195, LUT_AMPL_WIDTH - 1),
		21961 => to_unsigned(28194, LUT_AMPL_WIDTH - 1),
		21962 => to_unsigned(28192, LUT_AMPL_WIDTH - 1),
		21963 => to_unsigned(28190, LUT_AMPL_WIDTH - 1),
		21964 => to_unsigned(28189, LUT_AMPL_WIDTH - 1),
		21965 => to_unsigned(28187, LUT_AMPL_WIDTH - 1),
		21966 => to_unsigned(28186, LUT_AMPL_WIDTH - 1),
		21967 => to_unsigned(28184, LUT_AMPL_WIDTH - 1),
		21968 => to_unsigned(28182, LUT_AMPL_WIDTH - 1),
		21969 => to_unsigned(28181, LUT_AMPL_WIDTH - 1),
		21970 => to_unsigned(28179, LUT_AMPL_WIDTH - 1),
		21971 => to_unsigned(28178, LUT_AMPL_WIDTH - 1),
		21972 => to_unsigned(28176, LUT_AMPL_WIDTH - 1),
		21973 => to_unsigned(28174, LUT_AMPL_WIDTH - 1),
		21974 => to_unsigned(28173, LUT_AMPL_WIDTH - 1),
		21975 => to_unsigned(28171, LUT_AMPL_WIDTH - 1),
		21976 => to_unsigned(28170, LUT_AMPL_WIDTH - 1),
		21977 => to_unsigned(28168, LUT_AMPL_WIDTH - 1),
		21978 => to_unsigned(28166, LUT_AMPL_WIDTH - 1),
		21979 => to_unsigned(28165, LUT_AMPL_WIDTH - 1),
		21980 => to_unsigned(28163, LUT_AMPL_WIDTH - 1),
		21981 => to_unsigned(28162, LUT_AMPL_WIDTH - 1),
		21982 => to_unsigned(28160, LUT_AMPL_WIDTH - 1),
		21983 => to_unsigned(28158, LUT_AMPL_WIDTH - 1),
		21984 => to_unsigned(28157, LUT_AMPL_WIDTH - 1),
		21985 => to_unsigned(28155, LUT_AMPL_WIDTH - 1),
		21986 => to_unsigned(28154, LUT_AMPL_WIDTH - 1),
		21987 => to_unsigned(28152, LUT_AMPL_WIDTH - 1),
		21988 => to_unsigned(28150, LUT_AMPL_WIDTH - 1),
		21989 => to_unsigned(28149, LUT_AMPL_WIDTH - 1),
		21990 => to_unsigned(28147, LUT_AMPL_WIDTH - 1),
		21991 => to_unsigned(28145, LUT_AMPL_WIDTH - 1),
		21992 => to_unsigned(28144, LUT_AMPL_WIDTH - 1),
		21993 => to_unsigned(28142, LUT_AMPL_WIDTH - 1),
		21994 => to_unsigned(28141, LUT_AMPL_WIDTH - 1),
		21995 => to_unsigned(28139, LUT_AMPL_WIDTH - 1),
		21996 => to_unsigned(28137, LUT_AMPL_WIDTH - 1),
		21997 => to_unsigned(28136, LUT_AMPL_WIDTH - 1),
		21998 => to_unsigned(28134, LUT_AMPL_WIDTH - 1),
		21999 => to_unsigned(28133, LUT_AMPL_WIDTH - 1),
		22000 => to_unsigned(28131, LUT_AMPL_WIDTH - 1),
		22001 => to_unsigned(28129, LUT_AMPL_WIDTH - 1),
		22002 => to_unsigned(28128, LUT_AMPL_WIDTH - 1),
		22003 => to_unsigned(28126, LUT_AMPL_WIDTH - 1),
		22004 => to_unsigned(28125, LUT_AMPL_WIDTH - 1),
		22005 => to_unsigned(28123, LUT_AMPL_WIDTH - 1),
		22006 => to_unsigned(28121, LUT_AMPL_WIDTH - 1),
		22007 => to_unsigned(28120, LUT_AMPL_WIDTH - 1),
		22008 => to_unsigned(28118, LUT_AMPL_WIDTH - 1),
		22009 => to_unsigned(28116, LUT_AMPL_WIDTH - 1),
		22010 => to_unsigned(28115, LUT_AMPL_WIDTH - 1),
		22011 => to_unsigned(28113, LUT_AMPL_WIDTH - 1),
		22012 => to_unsigned(28112, LUT_AMPL_WIDTH - 1),
		22013 => to_unsigned(28110, LUT_AMPL_WIDTH - 1),
		22014 => to_unsigned(28108, LUT_AMPL_WIDTH - 1),
		22015 => to_unsigned(28107, LUT_AMPL_WIDTH - 1),
		22016 => to_unsigned(28105, LUT_AMPL_WIDTH - 1),
		22017 => to_unsigned(28104, LUT_AMPL_WIDTH - 1),
		22018 => to_unsigned(28102, LUT_AMPL_WIDTH - 1),
		22019 => to_unsigned(28100, LUT_AMPL_WIDTH - 1),
		22020 => to_unsigned(28099, LUT_AMPL_WIDTH - 1),
		22021 => to_unsigned(28097, LUT_AMPL_WIDTH - 1),
		22022 => to_unsigned(28095, LUT_AMPL_WIDTH - 1),
		22023 => to_unsigned(28094, LUT_AMPL_WIDTH - 1),
		22024 => to_unsigned(28092, LUT_AMPL_WIDTH - 1),
		22025 => to_unsigned(28091, LUT_AMPL_WIDTH - 1),
		22026 => to_unsigned(28089, LUT_AMPL_WIDTH - 1),
		22027 => to_unsigned(28087, LUT_AMPL_WIDTH - 1),
		22028 => to_unsigned(28086, LUT_AMPL_WIDTH - 1),
		22029 => to_unsigned(28084, LUT_AMPL_WIDTH - 1),
		22030 => to_unsigned(28083, LUT_AMPL_WIDTH - 1),
		22031 => to_unsigned(28081, LUT_AMPL_WIDTH - 1),
		22032 => to_unsigned(28079, LUT_AMPL_WIDTH - 1),
		22033 => to_unsigned(28078, LUT_AMPL_WIDTH - 1),
		22034 => to_unsigned(28076, LUT_AMPL_WIDTH - 1),
		22035 => to_unsigned(28074, LUT_AMPL_WIDTH - 1),
		22036 => to_unsigned(28073, LUT_AMPL_WIDTH - 1),
		22037 => to_unsigned(28071, LUT_AMPL_WIDTH - 1),
		22038 => to_unsigned(28070, LUT_AMPL_WIDTH - 1),
		22039 => to_unsigned(28068, LUT_AMPL_WIDTH - 1),
		22040 => to_unsigned(28066, LUT_AMPL_WIDTH - 1),
		22041 => to_unsigned(28065, LUT_AMPL_WIDTH - 1),
		22042 => to_unsigned(28063, LUT_AMPL_WIDTH - 1),
		22043 => to_unsigned(28061, LUT_AMPL_WIDTH - 1),
		22044 => to_unsigned(28060, LUT_AMPL_WIDTH - 1),
		22045 => to_unsigned(28058, LUT_AMPL_WIDTH - 1),
		22046 => to_unsigned(28057, LUT_AMPL_WIDTH - 1),
		22047 => to_unsigned(28055, LUT_AMPL_WIDTH - 1),
		22048 => to_unsigned(28053, LUT_AMPL_WIDTH - 1),
		22049 => to_unsigned(28052, LUT_AMPL_WIDTH - 1),
		22050 => to_unsigned(28050, LUT_AMPL_WIDTH - 1),
		22051 => to_unsigned(28049, LUT_AMPL_WIDTH - 1),
		22052 => to_unsigned(28047, LUT_AMPL_WIDTH - 1),
		22053 => to_unsigned(28045, LUT_AMPL_WIDTH - 1),
		22054 => to_unsigned(28044, LUT_AMPL_WIDTH - 1),
		22055 => to_unsigned(28042, LUT_AMPL_WIDTH - 1),
		22056 => to_unsigned(28040, LUT_AMPL_WIDTH - 1),
		22057 => to_unsigned(28039, LUT_AMPL_WIDTH - 1),
		22058 => to_unsigned(28037, LUT_AMPL_WIDTH - 1),
		22059 => to_unsigned(28036, LUT_AMPL_WIDTH - 1),
		22060 => to_unsigned(28034, LUT_AMPL_WIDTH - 1),
		22061 => to_unsigned(28032, LUT_AMPL_WIDTH - 1),
		22062 => to_unsigned(28031, LUT_AMPL_WIDTH - 1),
		22063 => to_unsigned(28029, LUT_AMPL_WIDTH - 1),
		22064 => to_unsigned(28027, LUT_AMPL_WIDTH - 1),
		22065 => to_unsigned(28026, LUT_AMPL_WIDTH - 1),
		22066 => to_unsigned(28024, LUT_AMPL_WIDTH - 1),
		22067 => to_unsigned(28022, LUT_AMPL_WIDTH - 1),
		22068 => to_unsigned(28021, LUT_AMPL_WIDTH - 1),
		22069 => to_unsigned(28019, LUT_AMPL_WIDTH - 1),
		22070 => to_unsigned(28018, LUT_AMPL_WIDTH - 1),
		22071 => to_unsigned(28016, LUT_AMPL_WIDTH - 1),
		22072 => to_unsigned(28014, LUT_AMPL_WIDTH - 1),
		22073 => to_unsigned(28013, LUT_AMPL_WIDTH - 1),
		22074 => to_unsigned(28011, LUT_AMPL_WIDTH - 1),
		22075 => to_unsigned(28009, LUT_AMPL_WIDTH - 1),
		22076 => to_unsigned(28008, LUT_AMPL_WIDTH - 1),
		22077 => to_unsigned(28006, LUT_AMPL_WIDTH - 1),
		22078 => to_unsigned(28005, LUT_AMPL_WIDTH - 1),
		22079 => to_unsigned(28003, LUT_AMPL_WIDTH - 1),
		22080 => to_unsigned(28001, LUT_AMPL_WIDTH - 1),
		22081 => to_unsigned(28000, LUT_AMPL_WIDTH - 1),
		22082 => to_unsigned(27998, LUT_AMPL_WIDTH - 1),
		22083 => to_unsigned(27996, LUT_AMPL_WIDTH - 1),
		22084 => to_unsigned(27995, LUT_AMPL_WIDTH - 1),
		22085 => to_unsigned(27993, LUT_AMPL_WIDTH - 1),
		22086 => to_unsigned(27992, LUT_AMPL_WIDTH - 1),
		22087 => to_unsigned(27990, LUT_AMPL_WIDTH - 1),
		22088 => to_unsigned(27988, LUT_AMPL_WIDTH - 1),
		22089 => to_unsigned(27987, LUT_AMPL_WIDTH - 1),
		22090 => to_unsigned(27985, LUT_AMPL_WIDTH - 1),
		22091 => to_unsigned(27983, LUT_AMPL_WIDTH - 1),
		22092 => to_unsigned(27982, LUT_AMPL_WIDTH - 1),
		22093 => to_unsigned(27980, LUT_AMPL_WIDTH - 1),
		22094 => to_unsigned(27978, LUT_AMPL_WIDTH - 1),
		22095 => to_unsigned(27977, LUT_AMPL_WIDTH - 1),
		22096 => to_unsigned(27975, LUT_AMPL_WIDTH - 1),
		22097 => to_unsigned(27974, LUT_AMPL_WIDTH - 1),
		22098 => to_unsigned(27972, LUT_AMPL_WIDTH - 1),
		22099 => to_unsigned(27970, LUT_AMPL_WIDTH - 1),
		22100 => to_unsigned(27969, LUT_AMPL_WIDTH - 1),
		22101 => to_unsigned(27967, LUT_AMPL_WIDTH - 1),
		22102 => to_unsigned(27965, LUT_AMPL_WIDTH - 1),
		22103 => to_unsigned(27964, LUT_AMPL_WIDTH - 1),
		22104 => to_unsigned(27962, LUT_AMPL_WIDTH - 1),
		22105 => to_unsigned(27960, LUT_AMPL_WIDTH - 1),
		22106 => to_unsigned(27959, LUT_AMPL_WIDTH - 1),
		22107 => to_unsigned(27957, LUT_AMPL_WIDTH - 1),
		22108 => to_unsigned(27956, LUT_AMPL_WIDTH - 1),
		22109 => to_unsigned(27954, LUT_AMPL_WIDTH - 1),
		22110 => to_unsigned(27952, LUT_AMPL_WIDTH - 1),
		22111 => to_unsigned(27951, LUT_AMPL_WIDTH - 1),
		22112 => to_unsigned(27949, LUT_AMPL_WIDTH - 1),
		22113 => to_unsigned(27947, LUT_AMPL_WIDTH - 1),
		22114 => to_unsigned(27946, LUT_AMPL_WIDTH - 1),
		22115 => to_unsigned(27944, LUT_AMPL_WIDTH - 1),
		22116 => to_unsigned(27942, LUT_AMPL_WIDTH - 1),
		22117 => to_unsigned(27941, LUT_AMPL_WIDTH - 1),
		22118 => to_unsigned(27939, LUT_AMPL_WIDTH - 1),
		22119 => to_unsigned(27937, LUT_AMPL_WIDTH - 1),
		22120 => to_unsigned(27936, LUT_AMPL_WIDTH - 1),
		22121 => to_unsigned(27934, LUT_AMPL_WIDTH - 1),
		22122 => to_unsigned(27933, LUT_AMPL_WIDTH - 1),
		22123 => to_unsigned(27931, LUT_AMPL_WIDTH - 1),
		22124 => to_unsigned(27929, LUT_AMPL_WIDTH - 1),
		22125 => to_unsigned(27928, LUT_AMPL_WIDTH - 1),
		22126 => to_unsigned(27926, LUT_AMPL_WIDTH - 1),
		22127 => to_unsigned(27924, LUT_AMPL_WIDTH - 1),
		22128 => to_unsigned(27923, LUT_AMPL_WIDTH - 1),
		22129 => to_unsigned(27921, LUT_AMPL_WIDTH - 1),
		22130 => to_unsigned(27919, LUT_AMPL_WIDTH - 1),
		22131 => to_unsigned(27918, LUT_AMPL_WIDTH - 1),
		22132 => to_unsigned(27916, LUT_AMPL_WIDTH - 1),
		22133 => to_unsigned(27914, LUT_AMPL_WIDTH - 1),
		22134 => to_unsigned(27913, LUT_AMPL_WIDTH - 1),
		22135 => to_unsigned(27911, LUT_AMPL_WIDTH - 1),
		22136 => to_unsigned(27910, LUT_AMPL_WIDTH - 1),
		22137 => to_unsigned(27908, LUT_AMPL_WIDTH - 1),
		22138 => to_unsigned(27906, LUT_AMPL_WIDTH - 1),
		22139 => to_unsigned(27905, LUT_AMPL_WIDTH - 1),
		22140 => to_unsigned(27903, LUT_AMPL_WIDTH - 1),
		22141 => to_unsigned(27901, LUT_AMPL_WIDTH - 1),
		22142 => to_unsigned(27900, LUT_AMPL_WIDTH - 1),
		22143 => to_unsigned(27898, LUT_AMPL_WIDTH - 1),
		22144 => to_unsigned(27896, LUT_AMPL_WIDTH - 1),
		22145 => to_unsigned(27895, LUT_AMPL_WIDTH - 1),
		22146 => to_unsigned(27893, LUT_AMPL_WIDTH - 1),
		22147 => to_unsigned(27891, LUT_AMPL_WIDTH - 1),
		22148 => to_unsigned(27890, LUT_AMPL_WIDTH - 1),
		22149 => to_unsigned(27888, LUT_AMPL_WIDTH - 1),
		22150 => to_unsigned(27886, LUT_AMPL_WIDTH - 1),
		22151 => to_unsigned(27885, LUT_AMPL_WIDTH - 1),
		22152 => to_unsigned(27883, LUT_AMPL_WIDTH - 1),
		22153 => to_unsigned(27882, LUT_AMPL_WIDTH - 1),
		22154 => to_unsigned(27880, LUT_AMPL_WIDTH - 1),
		22155 => to_unsigned(27878, LUT_AMPL_WIDTH - 1),
		22156 => to_unsigned(27877, LUT_AMPL_WIDTH - 1),
		22157 => to_unsigned(27875, LUT_AMPL_WIDTH - 1),
		22158 => to_unsigned(27873, LUT_AMPL_WIDTH - 1),
		22159 => to_unsigned(27872, LUT_AMPL_WIDTH - 1),
		22160 => to_unsigned(27870, LUT_AMPL_WIDTH - 1),
		22161 => to_unsigned(27868, LUT_AMPL_WIDTH - 1),
		22162 => to_unsigned(27867, LUT_AMPL_WIDTH - 1),
		22163 => to_unsigned(27865, LUT_AMPL_WIDTH - 1),
		22164 => to_unsigned(27863, LUT_AMPL_WIDTH - 1),
		22165 => to_unsigned(27862, LUT_AMPL_WIDTH - 1),
		22166 => to_unsigned(27860, LUT_AMPL_WIDTH - 1),
		22167 => to_unsigned(27858, LUT_AMPL_WIDTH - 1),
		22168 => to_unsigned(27857, LUT_AMPL_WIDTH - 1),
		22169 => to_unsigned(27855, LUT_AMPL_WIDTH - 1),
		22170 => to_unsigned(27853, LUT_AMPL_WIDTH - 1),
		22171 => to_unsigned(27852, LUT_AMPL_WIDTH - 1),
		22172 => to_unsigned(27850, LUT_AMPL_WIDTH - 1),
		22173 => to_unsigned(27848, LUT_AMPL_WIDTH - 1),
		22174 => to_unsigned(27847, LUT_AMPL_WIDTH - 1),
		22175 => to_unsigned(27845, LUT_AMPL_WIDTH - 1),
		22176 => to_unsigned(27843, LUT_AMPL_WIDTH - 1),
		22177 => to_unsigned(27842, LUT_AMPL_WIDTH - 1),
		22178 => to_unsigned(27840, LUT_AMPL_WIDTH - 1),
		22179 => to_unsigned(27839, LUT_AMPL_WIDTH - 1),
		22180 => to_unsigned(27837, LUT_AMPL_WIDTH - 1),
		22181 => to_unsigned(27835, LUT_AMPL_WIDTH - 1),
		22182 => to_unsigned(27834, LUT_AMPL_WIDTH - 1),
		22183 => to_unsigned(27832, LUT_AMPL_WIDTH - 1),
		22184 => to_unsigned(27830, LUT_AMPL_WIDTH - 1),
		22185 => to_unsigned(27829, LUT_AMPL_WIDTH - 1),
		22186 => to_unsigned(27827, LUT_AMPL_WIDTH - 1),
		22187 => to_unsigned(27825, LUT_AMPL_WIDTH - 1),
		22188 => to_unsigned(27824, LUT_AMPL_WIDTH - 1),
		22189 => to_unsigned(27822, LUT_AMPL_WIDTH - 1),
		22190 => to_unsigned(27820, LUT_AMPL_WIDTH - 1),
		22191 => to_unsigned(27819, LUT_AMPL_WIDTH - 1),
		22192 => to_unsigned(27817, LUT_AMPL_WIDTH - 1),
		22193 => to_unsigned(27815, LUT_AMPL_WIDTH - 1),
		22194 => to_unsigned(27814, LUT_AMPL_WIDTH - 1),
		22195 => to_unsigned(27812, LUT_AMPL_WIDTH - 1),
		22196 => to_unsigned(27810, LUT_AMPL_WIDTH - 1),
		22197 => to_unsigned(27809, LUT_AMPL_WIDTH - 1),
		22198 => to_unsigned(27807, LUT_AMPL_WIDTH - 1),
		22199 => to_unsigned(27805, LUT_AMPL_WIDTH - 1),
		22200 => to_unsigned(27804, LUT_AMPL_WIDTH - 1),
		22201 => to_unsigned(27802, LUT_AMPL_WIDTH - 1),
		22202 => to_unsigned(27800, LUT_AMPL_WIDTH - 1),
		22203 => to_unsigned(27799, LUT_AMPL_WIDTH - 1),
		22204 => to_unsigned(27797, LUT_AMPL_WIDTH - 1),
		22205 => to_unsigned(27795, LUT_AMPL_WIDTH - 1),
		22206 => to_unsigned(27794, LUT_AMPL_WIDTH - 1),
		22207 => to_unsigned(27792, LUT_AMPL_WIDTH - 1),
		22208 => to_unsigned(27790, LUT_AMPL_WIDTH - 1),
		22209 => to_unsigned(27789, LUT_AMPL_WIDTH - 1),
		22210 => to_unsigned(27787, LUT_AMPL_WIDTH - 1),
		22211 => to_unsigned(27785, LUT_AMPL_WIDTH - 1),
		22212 => to_unsigned(27784, LUT_AMPL_WIDTH - 1),
		22213 => to_unsigned(27782, LUT_AMPL_WIDTH - 1),
		22214 => to_unsigned(27780, LUT_AMPL_WIDTH - 1),
		22215 => to_unsigned(27779, LUT_AMPL_WIDTH - 1),
		22216 => to_unsigned(27777, LUT_AMPL_WIDTH - 1),
		22217 => to_unsigned(27775, LUT_AMPL_WIDTH - 1),
		22218 => to_unsigned(27774, LUT_AMPL_WIDTH - 1),
		22219 => to_unsigned(27772, LUT_AMPL_WIDTH - 1),
		22220 => to_unsigned(27770, LUT_AMPL_WIDTH - 1),
		22221 => to_unsigned(27769, LUT_AMPL_WIDTH - 1),
		22222 => to_unsigned(27767, LUT_AMPL_WIDTH - 1),
		22223 => to_unsigned(27765, LUT_AMPL_WIDTH - 1),
		22224 => to_unsigned(27764, LUT_AMPL_WIDTH - 1),
		22225 => to_unsigned(27762, LUT_AMPL_WIDTH - 1),
		22226 => to_unsigned(27760, LUT_AMPL_WIDTH - 1),
		22227 => to_unsigned(27759, LUT_AMPL_WIDTH - 1),
		22228 => to_unsigned(27757, LUT_AMPL_WIDTH - 1),
		22229 => to_unsigned(27755, LUT_AMPL_WIDTH - 1),
		22230 => to_unsigned(27754, LUT_AMPL_WIDTH - 1),
		22231 => to_unsigned(27752, LUT_AMPL_WIDTH - 1),
		22232 => to_unsigned(27750, LUT_AMPL_WIDTH - 1),
		22233 => to_unsigned(27749, LUT_AMPL_WIDTH - 1),
		22234 => to_unsigned(27747, LUT_AMPL_WIDTH - 1),
		22235 => to_unsigned(27745, LUT_AMPL_WIDTH - 1),
		22236 => to_unsigned(27744, LUT_AMPL_WIDTH - 1),
		22237 => to_unsigned(27742, LUT_AMPL_WIDTH - 1),
		22238 => to_unsigned(27740, LUT_AMPL_WIDTH - 1),
		22239 => to_unsigned(27739, LUT_AMPL_WIDTH - 1),
		22240 => to_unsigned(27737, LUT_AMPL_WIDTH - 1),
		22241 => to_unsigned(27735, LUT_AMPL_WIDTH - 1),
		22242 => to_unsigned(27734, LUT_AMPL_WIDTH - 1),
		22243 => to_unsigned(27732, LUT_AMPL_WIDTH - 1),
		22244 => to_unsigned(27730, LUT_AMPL_WIDTH - 1),
		22245 => to_unsigned(27729, LUT_AMPL_WIDTH - 1),
		22246 => to_unsigned(27727, LUT_AMPL_WIDTH - 1),
		22247 => to_unsigned(27725, LUT_AMPL_WIDTH - 1),
		22248 => to_unsigned(27724, LUT_AMPL_WIDTH - 1),
		22249 => to_unsigned(27722, LUT_AMPL_WIDTH - 1),
		22250 => to_unsigned(27720, LUT_AMPL_WIDTH - 1),
		22251 => to_unsigned(27719, LUT_AMPL_WIDTH - 1),
		22252 => to_unsigned(27717, LUT_AMPL_WIDTH - 1),
		22253 => to_unsigned(27715, LUT_AMPL_WIDTH - 1),
		22254 => to_unsigned(27714, LUT_AMPL_WIDTH - 1),
		22255 => to_unsigned(27712, LUT_AMPL_WIDTH - 1),
		22256 => to_unsigned(27710, LUT_AMPL_WIDTH - 1),
		22257 => to_unsigned(27708, LUT_AMPL_WIDTH - 1),
		22258 => to_unsigned(27707, LUT_AMPL_WIDTH - 1),
		22259 => to_unsigned(27705, LUT_AMPL_WIDTH - 1),
		22260 => to_unsigned(27703, LUT_AMPL_WIDTH - 1),
		22261 => to_unsigned(27702, LUT_AMPL_WIDTH - 1),
		22262 => to_unsigned(27700, LUT_AMPL_WIDTH - 1),
		22263 => to_unsigned(27698, LUT_AMPL_WIDTH - 1),
		22264 => to_unsigned(27697, LUT_AMPL_WIDTH - 1),
		22265 => to_unsigned(27695, LUT_AMPL_WIDTH - 1),
		22266 => to_unsigned(27693, LUT_AMPL_WIDTH - 1),
		22267 => to_unsigned(27692, LUT_AMPL_WIDTH - 1),
		22268 => to_unsigned(27690, LUT_AMPL_WIDTH - 1),
		22269 => to_unsigned(27688, LUT_AMPL_WIDTH - 1),
		22270 => to_unsigned(27687, LUT_AMPL_WIDTH - 1),
		22271 => to_unsigned(27685, LUT_AMPL_WIDTH - 1),
		22272 => to_unsigned(27683, LUT_AMPL_WIDTH - 1),
		22273 => to_unsigned(27682, LUT_AMPL_WIDTH - 1),
		22274 => to_unsigned(27680, LUT_AMPL_WIDTH - 1),
		22275 => to_unsigned(27678, LUT_AMPL_WIDTH - 1),
		22276 => to_unsigned(27677, LUT_AMPL_WIDTH - 1),
		22277 => to_unsigned(27675, LUT_AMPL_WIDTH - 1),
		22278 => to_unsigned(27673, LUT_AMPL_WIDTH - 1),
		22279 => to_unsigned(27672, LUT_AMPL_WIDTH - 1),
		22280 => to_unsigned(27670, LUT_AMPL_WIDTH - 1),
		22281 => to_unsigned(27668, LUT_AMPL_WIDTH - 1),
		22282 => to_unsigned(27666, LUT_AMPL_WIDTH - 1),
		22283 => to_unsigned(27665, LUT_AMPL_WIDTH - 1),
		22284 => to_unsigned(27663, LUT_AMPL_WIDTH - 1),
		22285 => to_unsigned(27661, LUT_AMPL_WIDTH - 1),
		22286 => to_unsigned(27660, LUT_AMPL_WIDTH - 1),
		22287 => to_unsigned(27658, LUT_AMPL_WIDTH - 1),
		22288 => to_unsigned(27656, LUT_AMPL_WIDTH - 1),
		22289 => to_unsigned(27655, LUT_AMPL_WIDTH - 1),
		22290 => to_unsigned(27653, LUT_AMPL_WIDTH - 1),
		22291 => to_unsigned(27651, LUT_AMPL_WIDTH - 1),
		22292 => to_unsigned(27650, LUT_AMPL_WIDTH - 1),
		22293 => to_unsigned(27648, LUT_AMPL_WIDTH - 1),
		22294 => to_unsigned(27646, LUT_AMPL_WIDTH - 1),
		22295 => to_unsigned(27645, LUT_AMPL_WIDTH - 1),
		22296 => to_unsigned(27643, LUT_AMPL_WIDTH - 1),
		22297 => to_unsigned(27641, LUT_AMPL_WIDTH - 1),
		22298 => to_unsigned(27640, LUT_AMPL_WIDTH - 1),
		22299 => to_unsigned(27638, LUT_AMPL_WIDTH - 1),
		22300 => to_unsigned(27636, LUT_AMPL_WIDTH - 1),
		22301 => to_unsigned(27634, LUT_AMPL_WIDTH - 1),
		22302 => to_unsigned(27633, LUT_AMPL_WIDTH - 1),
		22303 => to_unsigned(27631, LUT_AMPL_WIDTH - 1),
		22304 => to_unsigned(27629, LUT_AMPL_WIDTH - 1),
		22305 => to_unsigned(27628, LUT_AMPL_WIDTH - 1),
		22306 => to_unsigned(27626, LUT_AMPL_WIDTH - 1),
		22307 => to_unsigned(27624, LUT_AMPL_WIDTH - 1),
		22308 => to_unsigned(27623, LUT_AMPL_WIDTH - 1),
		22309 => to_unsigned(27621, LUT_AMPL_WIDTH - 1),
		22310 => to_unsigned(27619, LUT_AMPL_WIDTH - 1),
		22311 => to_unsigned(27618, LUT_AMPL_WIDTH - 1),
		22312 => to_unsigned(27616, LUT_AMPL_WIDTH - 1),
		22313 => to_unsigned(27614, LUT_AMPL_WIDTH - 1),
		22314 => to_unsigned(27613, LUT_AMPL_WIDTH - 1),
		22315 => to_unsigned(27611, LUT_AMPL_WIDTH - 1),
		22316 => to_unsigned(27609, LUT_AMPL_WIDTH - 1),
		22317 => to_unsigned(27607, LUT_AMPL_WIDTH - 1),
		22318 => to_unsigned(27606, LUT_AMPL_WIDTH - 1),
		22319 => to_unsigned(27604, LUT_AMPL_WIDTH - 1),
		22320 => to_unsigned(27602, LUT_AMPL_WIDTH - 1),
		22321 => to_unsigned(27601, LUT_AMPL_WIDTH - 1),
		22322 => to_unsigned(27599, LUT_AMPL_WIDTH - 1),
		22323 => to_unsigned(27597, LUT_AMPL_WIDTH - 1),
		22324 => to_unsigned(27596, LUT_AMPL_WIDTH - 1),
		22325 => to_unsigned(27594, LUT_AMPL_WIDTH - 1),
		22326 => to_unsigned(27592, LUT_AMPL_WIDTH - 1),
		22327 => to_unsigned(27590, LUT_AMPL_WIDTH - 1),
		22328 => to_unsigned(27589, LUT_AMPL_WIDTH - 1),
		22329 => to_unsigned(27587, LUT_AMPL_WIDTH - 1),
		22330 => to_unsigned(27585, LUT_AMPL_WIDTH - 1),
		22331 => to_unsigned(27584, LUT_AMPL_WIDTH - 1),
		22332 => to_unsigned(27582, LUT_AMPL_WIDTH - 1),
		22333 => to_unsigned(27580, LUT_AMPL_WIDTH - 1),
		22334 => to_unsigned(27579, LUT_AMPL_WIDTH - 1),
		22335 => to_unsigned(27577, LUT_AMPL_WIDTH - 1),
		22336 => to_unsigned(27575, LUT_AMPL_WIDTH - 1),
		22337 => to_unsigned(27574, LUT_AMPL_WIDTH - 1),
		22338 => to_unsigned(27572, LUT_AMPL_WIDTH - 1),
		22339 => to_unsigned(27570, LUT_AMPL_WIDTH - 1),
		22340 => to_unsigned(27568, LUT_AMPL_WIDTH - 1),
		22341 => to_unsigned(27567, LUT_AMPL_WIDTH - 1),
		22342 => to_unsigned(27565, LUT_AMPL_WIDTH - 1),
		22343 => to_unsigned(27563, LUT_AMPL_WIDTH - 1),
		22344 => to_unsigned(27562, LUT_AMPL_WIDTH - 1),
		22345 => to_unsigned(27560, LUT_AMPL_WIDTH - 1),
		22346 => to_unsigned(27558, LUT_AMPL_WIDTH - 1),
		22347 => to_unsigned(27557, LUT_AMPL_WIDTH - 1),
		22348 => to_unsigned(27555, LUT_AMPL_WIDTH - 1),
		22349 => to_unsigned(27553, LUT_AMPL_WIDTH - 1),
		22350 => to_unsigned(27551, LUT_AMPL_WIDTH - 1),
		22351 => to_unsigned(27550, LUT_AMPL_WIDTH - 1),
		22352 => to_unsigned(27548, LUT_AMPL_WIDTH - 1),
		22353 => to_unsigned(27546, LUT_AMPL_WIDTH - 1),
		22354 => to_unsigned(27545, LUT_AMPL_WIDTH - 1),
		22355 => to_unsigned(27543, LUT_AMPL_WIDTH - 1),
		22356 => to_unsigned(27541, LUT_AMPL_WIDTH - 1),
		22357 => to_unsigned(27540, LUT_AMPL_WIDTH - 1),
		22358 => to_unsigned(27538, LUT_AMPL_WIDTH - 1),
		22359 => to_unsigned(27536, LUT_AMPL_WIDTH - 1),
		22360 => to_unsigned(27534, LUT_AMPL_WIDTH - 1),
		22361 => to_unsigned(27533, LUT_AMPL_WIDTH - 1),
		22362 => to_unsigned(27531, LUT_AMPL_WIDTH - 1),
		22363 => to_unsigned(27529, LUT_AMPL_WIDTH - 1),
		22364 => to_unsigned(27528, LUT_AMPL_WIDTH - 1),
		22365 => to_unsigned(27526, LUT_AMPL_WIDTH - 1),
		22366 => to_unsigned(27524, LUT_AMPL_WIDTH - 1),
		22367 => to_unsigned(27523, LUT_AMPL_WIDTH - 1),
		22368 => to_unsigned(27521, LUT_AMPL_WIDTH - 1),
		22369 => to_unsigned(27519, LUT_AMPL_WIDTH - 1),
		22370 => to_unsigned(27517, LUT_AMPL_WIDTH - 1),
		22371 => to_unsigned(27516, LUT_AMPL_WIDTH - 1),
		22372 => to_unsigned(27514, LUT_AMPL_WIDTH - 1),
		22373 => to_unsigned(27512, LUT_AMPL_WIDTH - 1),
		22374 => to_unsigned(27511, LUT_AMPL_WIDTH - 1),
		22375 => to_unsigned(27509, LUT_AMPL_WIDTH - 1),
		22376 => to_unsigned(27507, LUT_AMPL_WIDTH - 1),
		22377 => to_unsigned(27505, LUT_AMPL_WIDTH - 1),
		22378 => to_unsigned(27504, LUT_AMPL_WIDTH - 1),
		22379 => to_unsigned(27502, LUT_AMPL_WIDTH - 1),
		22380 => to_unsigned(27500, LUT_AMPL_WIDTH - 1),
		22381 => to_unsigned(27499, LUT_AMPL_WIDTH - 1),
		22382 => to_unsigned(27497, LUT_AMPL_WIDTH - 1),
		22383 => to_unsigned(27495, LUT_AMPL_WIDTH - 1),
		22384 => to_unsigned(27493, LUT_AMPL_WIDTH - 1),
		22385 => to_unsigned(27492, LUT_AMPL_WIDTH - 1),
		22386 => to_unsigned(27490, LUT_AMPL_WIDTH - 1),
		22387 => to_unsigned(27488, LUT_AMPL_WIDTH - 1),
		22388 => to_unsigned(27487, LUT_AMPL_WIDTH - 1),
		22389 => to_unsigned(27485, LUT_AMPL_WIDTH - 1),
		22390 => to_unsigned(27483, LUT_AMPL_WIDTH - 1),
		22391 => to_unsigned(27482, LUT_AMPL_WIDTH - 1),
		22392 => to_unsigned(27480, LUT_AMPL_WIDTH - 1),
		22393 => to_unsigned(27478, LUT_AMPL_WIDTH - 1),
		22394 => to_unsigned(27476, LUT_AMPL_WIDTH - 1),
		22395 => to_unsigned(27475, LUT_AMPL_WIDTH - 1),
		22396 => to_unsigned(27473, LUT_AMPL_WIDTH - 1),
		22397 => to_unsigned(27471, LUT_AMPL_WIDTH - 1),
		22398 => to_unsigned(27470, LUT_AMPL_WIDTH - 1),
		22399 => to_unsigned(27468, LUT_AMPL_WIDTH - 1),
		22400 => to_unsigned(27466, LUT_AMPL_WIDTH - 1),
		22401 => to_unsigned(27464, LUT_AMPL_WIDTH - 1),
		22402 => to_unsigned(27463, LUT_AMPL_WIDTH - 1),
		22403 => to_unsigned(27461, LUT_AMPL_WIDTH - 1),
		22404 => to_unsigned(27459, LUT_AMPL_WIDTH - 1),
		22405 => to_unsigned(27458, LUT_AMPL_WIDTH - 1),
		22406 => to_unsigned(27456, LUT_AMPL_WIDTH - 1),
		22407 => to_unsigned(27454, LUT_AMPL_WIDTH - 1),
		22408 => to_unsigned(27452, LUT_AMPL_WIDTH - 1),
		22409 => to_unsigned(27451, LUT_AMPL_WIDTH - 1),
		22410 => to_unsigned(27449, LUT_AMPL_WIDTH - 1),
		22411 => to_unsigned(27447, LUT_AMPL_WIDTH - 1),
		22412 => to_unsigned(27446, LUT_AMPL_WIDTH - 1),
		22413 => to_unsigned(27444, LUT_AMPL_WIDTH - 1),
		22414 => to_unsigned(27442, LUT_AMPL_WIDTH - 1),
		22415 => to_unsigned(27440, LUT_AMPL_WIDTH - 1),
		22416 => to_unsigned(27439, LUT_AMPL_WIDTH - 1),
		22417 => to_unsigned(27437, LUT_AMPL_WIDTH - 1),
		22418 => to_unsigned(27435, LUT_AMPL_WIDTH - 1),
		22419 => to_unsigned(27434, LUT_AMPL_WIDTH - 1),
		22420 => to_unsigned(27432, LUT_AMPL_WIDTH - 1),
		22421 => to_unsigned(27430, LUT_AMPL_WIDTH - 1),
		22422 => to_unsigned(27428, LUT_AMPL_WIDTH - 1),
		22423 => to_unsigned(27427, LUT_AMPL_WIDTH - 1),
		22424 => to_unsigned(27425, LUT_AMPL_WIDTH - 1),
		22425 => to_unsigned(27423, LUT_AMPL_WIDTH - 1),
		22426 => to_unsigned(27421, LUT_AMPL_WIDTH - 1),
		22427 => to_unsigned(27420, LUT_AMPL_WIDTH - 1),
		22428 => to_unsigned(27418, LUT_AMPL_WIDTH - 1),
		22429 => to_unsigned(27416, LUT_AMPL_WIDTH - 1),
		22430 => to_unsigned(27415, LUT_AMPL_WIDTH - 1),
		22431 => to_unsigned(27413, LUT_AMPL_WIDTH - 1),
		22432 => to_unsigned(27411, LUT_AMPL_WIDTH - 1),
		22433 => to_unsigned(27409, LUT_AMPL_WIDTH - 1),
		22434 => to_unsigned(27408, LUT_AMPL_WIDTH - 1),
		22435 => to_unsigned(27406, LUT_AMPL_WIDTH - 1),
		22436 => to_unsigned(27404, LUT_AMPL_WIDTH - 1),
		22437 => to_unsigned(27403, LUT_AMPL_WIDTH - 1),
		22438 => to_unsigned(27401, LUT_AMPL_WIDTH - 1),
		22439 => to_unsigned(27399, LUT_AMPL_WIDTH - 1),
		22440 => to_unsigned(27397, LUT_AMPL_WIDTH - 1),
		22441 => to_unsigned(27396, LUT_AMPL_WIDTH - 1),
		22442 => to_unsigned(27394, LUT_AMPL_WIDTH - 1),
		22443 => to_unsigned(27392, LUT_AMPL_WIDTH - 1),
		22444 => to_unsigned(27390, LUT_AMPL_WIDTH - 1),
		22445 => to_unsigned(27389, LUT_AMPL_WIDTH - 1),
		22446 => to_unsigned(27387, LUT_AMPL_WIDTH - 1),
		22447 => to_unsigned(27385, LUT_AMPL_WIDTH - 1),
		22448 => to_unsigned(27384, LUT_AMPL_WIDTH - 1),
		22449 => to_unsigned(27382, LUT_AMPL_WIDTH - 1),
		22450 => to_unsigned(27380, LUT_AMPL_WIDTH - 1),
		22451 => to_unsigned(27378, LUT_AMPL_WIDTH - 1),
		22452 => to_unsigned(27377, LUT_AMPL_WIDTH - 1),
		22453 => to_unsigned(27375, LUT_AMPL_WIDTH - 1),
		22454 => to_unsigned(27373, LUT_AMPL_WIDTH - 1),
		22455 => to_unsigned(27372, LUT_AMPL_WIDTH - 1),
		22456 => to_unsigned(27370, LUT_AMPL_WIDTH - 1),
		22457 => to_unsigned(27368, LUT_AMPL_WIDTH - 1),
		22458 => to_unsigned(27366, LUT_AMPL_WIDTH - 1),
		22459 => to_unsigned(27365, LUT_AMPL_WIDTH - 1),
		22460 => to_unsigned(27363, LUT_AMPL_WIDTH - 1),
		22461 => to_unsigned(27361, LUT_AMPL_WIDTH - 1),
		22462 => to_unsigned(27359, LUT_AMPL_WIDTH - 1),
		22463 => to_unsigned(27358, LUT_AMPL_WIDTH - 1),
		22464 => to_unsigned(27356, LUT_AMPL_WIDTH - 1),
		22465 => to_unsigned(27354, LUT_AMPL_WIDTH - 1),
		22466 => to_unsigned(27352, LUT_AMPL_WIDTH - 1),
		22467 => to_unsigned(27351, LUT_AMPL_WIDTH - 1),
		22468 => to_unsigned(27349, LUT_AMPL_WIDTH - 1),
		22469 => to_unsigned(27347, LUT_AMPL_WIDTH - 1),
		22470 => to_unsigned(27346, LUT_AMPL_WIDTH - 1),
		22471 => to_unsigned(27344, LUT_AMPL_WIDTH - 1),
		22472 => to_unsigned(27342, LUT_AMPL_WIDTH - 1),
		22473 => to_unsigned(27340, LUT_AMPL_WIDTH - 1),
		22474 => to_unsigned(27339, LUT_AMPL_WIDTH - 1),
		22475 => to_unsigned(27337, LUT_AMPL_WIDTH - 1),
		22476 => to_unsigned(27335, LUT_AMPL_WIDTH - 1),
		22477 => to_unsigned(27333, LUT_AMPL_WIDTH - 1),
		22478 => to_unsigned(27332, LUT_AMPL_WIDTH - 1),
		22479 => to_unsigned(27330, LUT_AMPL_WIDTH - 1),
		22480 => to_unsigned(27328, LUT_AMPL_WIDTH - 1),
		22481 => to_unsigned(27327, LUT_AMPL_WIDTH - 1),
		22482 => to_unsigned(27325, LUT_AMPL_WIDTH - 1),
		22483 => to_unsigned(27323, LUT_AMPL_WIDTH - 1),
		22484 => to_unsigned(27321, LUT_AMPL_WIDTH - 1),
		22485 => to_unsigned(27320, LUT_AMPL_WIDTH - 1),
		22486 => to_unsigned(27318, LUT_AMPL_WIDTH - 1),
		22487 => to_unsigned(27316, LUT_AMPL_WIDTH - 1),
		22488 => to_unsigned(27314, LUT_AMPL_WIDTH - 1),
		22489 => to_unsigned(27313, LUT_AMPL_WIDTH - 1),
		22490 => to_unsigned(27311, LUT_AMPL_WIDTH - 1),
		22491 => to_unsigned(27309, LUT_AMPL_WIDTH - 1),
		22492 => to_unsigned(27307, LUT_AMPL_WIDTH - 1),
		22493 => to_unsigned(27306, LUT_AMPL_WIDTH - 1),
		22494 => to_unsigned(27304, LUT_AMPL_WIDTH - 1),
		22495 => to_unsigned(27302, LUT_AMPL_WIDTH - 1),
		22496 => to_unsigned(27300, LUT_AMPL_WIDTH - 1),
		22497 => to_unsigned(27299, LUT_AMPL_WIDTH - 1),
		22498 => to_unsigned(27297, LUT_AMPL_WIDTH - 1),
		22499 => to_unsigned(27295, LUT_AMPL_WIDTH - 1),
		22500 => to_unsigned(27294, LUT_AMPL_WIDTH - 1),
		22501 => to_unsigned(27292, LUT_AMPL_WIDTH - 1),
		22502 => to_unsigned(27290, LUT_AMPL_WIDTH - 1),
		22503 => to_unsigned(27288, LUT_AMPL_WIDTH - 1),
		22504 => to_unsigned(27287, LUT_AMPL_WIDTH - 1),
		22505 => to_unsigned(27285, LUT_AMPL_WIDTH - 1),
		22506 => to_unsigned(27283, LUT_AMPL_WIDTH - 1),
		22507 => to_unsigned(27281, LUT_AMPL_WIDTH - 1),
		22508 => to_unsigned(27280, LUT_AMPL_WIDTH - 1),
		22509 => to_unsigned(27278, LUT_AMPL_WIDTH - 1),
		22510 => to_unsigned(27276, LUT_AMPL_WIDTH - 1),
		22511 => to_unsigned(27274, LUT_AMPL_WIDTH - 1),
		22512 => to_unsigned(27273, LUT_AMPL_WIDTH - 1),
		22513 => to_unsigned(27271, LUT_AMPL_WIDTH - 1),
		22514 => to_unsigned(27269, LUT_AMPL_WIDTH - 1),
		22515 => to_unsigned(27267, LUT_AMPL_WIDTH - 1),
		22516 => to_unsigned(27266, LUT_AMPL_WIDTH - 1),
		22517 => to_unsigned(27264, LUT_AMPL_WIDTH - 1),
		22518 => to_unsigned(27262, LUT_AMPL_WIDTH - 1),
		22519 => to_unsigned(27260, LUT_AMPL_WIDTH - 1),
		22520 => to_unsigned(27259, LUT_AMPL_WIDTH - 1),
		22521 => to_unsigned(27257, LUT_AMPL_WIDTH - 1),
		22522 => to_unsigned(27255, LUT_AMPL_WIDTH - 1),
		22523 => to_unsigned(27253, LUT_AMPL_WIDTH - 1),
		22524 => to_unsigned(27252, LUT_AMPL_WIDTH - 1),
		22525 => to_unsigned(27250, LUT_AMPL_WIDTH - 1),
		22526 => to_unsigned(27248, LUT_AMPL_WIDTH - 1),
		22527 => to_unsigned(27247, LUT_AMPL_WIDTH - 1),
		22528 => to_unsigned(27245, LUT_AMPL_WIDTH - 1),
		22529 => to_unsigned(27243, LUT_AMPL_WIDTH - 1),
		22530 => to_unsigned(27241, LUT_AMPL_WIDTH - 1),
		22531 => to_unsigned(27240, LUT_AMPL_WIDTH - 1),
		22532 => to_unsigned(27238, LUT_AMPL_WIDTH - 1),
		22533 => to_unsigned(27236, LUT_AMPL_WIDTH - 1),
		22534 => to_unsigned(27234, LUT_AMPL_WIDTH - 1),
		22535 => to_unsigned(27233, LUT_AMPL_WIDTH - 1),
		22536 => to_unsigned(27231, LUT_AMPL_WIDTH - 1),
		22537 => to_unsigned(27229, LUT_AMPL_WIDTH - 1),
		22538 => to_unsigned(27227, LUT_AMPL_WIDTH - 1),
		22539 => to_unsigned(27226, LUT_AMPL_WIDTH - 1),
		22540 => to_unsigned(27224, LUT_AMPL_WIDTH - 1),
		22541 => to_unsigned(27222, LUT_AMPL_WIDTH - 1),
		22542 => to_unsigned(27220, LUT_AMPL_WIDTH - 1),
		22543 => to_unsigned(27219, LUT_AMPL_WIDTH - 1),
		22544 => to_unsigned(27217, LUT_AMPL_WIDTH - 1),
		22545 => to_unsigned(27215, LUT_AMPL_WIDTH - 1),
		22546 => to_unsigned(27213, LUT_AMPL_WIDTH - 1),
		22547 => to_unsigned(27212, LUT_AMPL_WIDTH - 1),
		22548 => to_unsigned(27210, LUT_AMPL_WIDTH - 1),
		22549 => to_unsigned(27208, LUT_AMPL_WIDTH - 1),
		22550 => to_unsigned(27206, LUT_AMPL_WIDTH - 1),
		22551 => to_unsigned(27205, LUT_AMPL_WIDTH - 1),
		22552 => to_unsigned(27203, LUT_AMPL_WIDTH - 1),
		22553 => to_unsigned(27201, LUT_AMPL_WIDTH - 1),
		22554 => to_unsigned(27199, LUT_AMPL_WIDTH - 1),
		22555 => to_unsigned(27198, LUT_AMPL_WIDTH - 1),
		22556 => to_unsigned(27196, LUT_AMPL_WIDTH - 1),
		22557 => to_unsigned(27194, LUT_AMPL_WIDTH - 1),
		22558 => to_unsigned(27192, LUT_AMPL_WIDTH - 1),
		22559 => to_unsigned(27191, LUT_AMPL_WIDTH - 1),
		22560 => to_unsigned(27189, LUT_AMPL_WIDTH - 1),
		22561 => to_unsigned(27187, LUT_AMPL_WIDTH - 1),
		22562 => to_unsigned(27185, LUT_AMPL_WIDTH - 1),
		22563 => to_unsigned(27184, LUT_AMPL_WIDTH - 1),
		22564 => to_unsigned(27182, LUT_AMPL_WIDTH - 1),
		22565 => to_unsigned(27180, LUT_AMPL_WIDTH - 1),
		22566 => to_unsigned(27178, LUT_AMPL_WIDTH - 1),
		22567 => to_unsigned(27177, LUT_AMPL_WIDTH - 1),
		22568 => to_unsigned(27175, LUT_AMPL_WIDTH - 1),
		22569 => to_unsigned(27173, LUT_AMPL_WIDTH - 1),
		22570 => to_unsigned(27171, LUT_AMPL_WIDTH - 1),
		22571 => to_unsigned(27169, LUT_AMPL_WIDTH - 1),
		22572 => to_unsigned(27168, LUT_AMPL_WIDTH - 1),
		22573 => to_unsigned(27166, LUT_AMPL_WIDTH - 1),
		22574 => to_unsigned(27164, LUT_AMPL_WIDTH - 1),
		22575 => to_unsigned(27162, LUT_AMPL_WIDTH - 1),
		22576 => to_unsigned(27161, LUT_AMPL_WIDTH - 1),
		22577 => to_unsigned(27159, LUT_AMPL_WIDTH - 1),
		22578 => to_unsigned(27157, LUT_AMPL_WIDTH - 1),
		22579 => to_unsigned(27155, LUT_AMPL_WIDTH - 1),
		22580 => to_unsigned(27154, LUT_AMPL_WIDTH - 1),
		22581 => to_unsigned(27152, LUT_AMPL_WIDTH - 1),
		22582 => to_unsigned(27150, LUT_AMPL_WIDTH - 1),
		22583 => to_unsigned(27148, LUT_AMPL_WIDTH - 1),
		22584 => to_unsigned(27147, LUT_AMPL_WIDTH - 1),
		22585 => to_unsigned(27145, LUT_AMPL_WIDTH - 1),
		22586 => to_unsigned(27143, LUT_AMPL_WIDTH - 1),
		22587 => to_unsigned(27141, LUT_AMPL_WIDTH - 1),
		22588 => to_unsigned(27140, LUT_AMPL_WIDTH - 1),
		22589 => to_unsigned(27138, LUT_AMPL_WIDTH - 1),
		22590 => to_unsigned(27136, LUT_AMPL_WIDTH - 1),
		22591 => to_unsigned(27134, LUT_AMPL_WIDTH - 1),
		22592 => to_unsigned(27133, LUT_AMPL_WIDTH - 1),
		22593 => to_unsigned(27131, LUT_AMPL_WIDTH - 1),
		22594 => to_unsigned(27129, LUT_AMPL_WIDTH - 1),
		22595 => to_unsigned(27127, LUT_AMPL_WIDTH - 1),
		22596 => to_unsigned(27126, LUT_AMPL_WIDTH - 1),
		22597 => to_unsigned(27124, LUT_AMPL_WIDTH - 1),
		22598 => to_unsigned(27122, LUT_AMPL_WIDTH - 1),
		22599 => to_unsigned(27120, LUT_AMPL_WIDTH - 1),
		22600 => to_unsigned(27118, LUT_AMPL_WIDTH - 1),
		22601 => to_unsigned(27117, LUT_AMPL_WIDTH - 1),
		22602 => to_unsigned(27115, LUT_AMPL_WIDTH - 1),
		22603 => to_unsigned(27113, LUT_AMPL_WIDTH - 1),
		22604 => to_unsigned(27111, LUT_AMPL_WIDTH - 1),
		22605 => to_unsigned(27110, LUT_AMPL_WIDTH - 1),
		22606 => to_unsigned(27108, LUT_AMPL_WIDTH - 1),
		22607 => to_unsigned(27106, LUT_AMPL_WIDTH - 1),
		22608 => to_unsigned(27104, LUT_AMPL_WIDTH - 1),
		22609 => to_unsigned(27103, LUT_AMPL_WIDTH - 1),
		22610 => to_unsigned(27101, LUT_AMPL_WIDTH - 1),
		22611 => to_unsigned(27099, LUT_AMPL_WIDTH - 1),
		22612 => to_unsigned(27097, LUT_AMPL_WIDTH - 1),
		22613 => to_unsigned(27096, LUT_AMPL_WIDTH - 1),
		22614 => to_unsigned(27094, LUT_AMPL_WIDTH - 1),
		22615 => to_unsigned(27092, LUT_AMPL_WIDTH - 1),
		22616 => to_unsigned(27090, LUT_AMPL_WIDTH - 1),
		22617 => to_unsigned(27088, LUT_AMPL_WIDTH - 1),
		22618 => to_unsigned(27087, LUT_AMPL_WIDTH - 1),
		22619 => to_unsigned(27085, LUT_AMPL_WIDTH - 1),
		22620 => to_unsigned(27083, LUT_AMPL_WIDTH - 1),
		22621 => to_unsigned(27081, LUT_AMPL_WIDTH - 1),
		22622 => to_unsigned(27080, LUT_AMPL_WIDTH - 1),
		22623 => to_unsigned(27078, LUT_AMPL_WIDTH - 1),
		22624 => to_unsigned(27076, LUT_AMPL_WIDTH - 1),
		22625 => to_unsigned(27074, LUT_AMPL_WIDTH - 1),
		22626 => to_unsigned(27073, LUT_AMPL_WIDTH - 1),
		22627 => to_unsigned(27071, LUT_AMPL_WIDTH - 1),
		22628 => to_unsigned(27069, LUT_AMPL_WIDTH - 1),
		22629 => to_unsigned(27067, LUT_AMPL_WIDTH - 1),
		22630 => to_unsigned(27065, LUT_AMPL_WIDTH - 1),
		22631 => to_unsigned(27064, LUT_AMPL_WIDTH - 1),
		22632 => to_unsigned(27062, LUT_AMPL_WIDTH - 1),
		22633 => to_unsigned(27060, LUT_AMPL_WIDTH - 1),
		22634 => to_unsigned(27058, LUT_AMPL_WIDTH - 1),
		22635 => to_unsigned(27057, LUT_AMPL_WIDTH - 1),
		22636 => to_unsigned(27055, LUT_AMPL_WIDTH - 1),
		22637 => to_unsigned(27053, LUT_AMPL_WIDTH - 1),
		22638 => to_unsigned(27051, LUT_AMPL_WIDTH - 1),
		22639 => to_unsigned(27049, LUT_AMPL_WIDTH - 1),
		22640 => to_unsigned(27048, LUT_AMPL_WIDTH - 1),
		22641 => to_unsigned(27046, LUT_AMPL_WIDTH - 1),
		22642 => to_unsigned(27044, LUT_AMPL_WIDTH - 1),
		22643 => to_unsigned(27042, LUT_AMPL_WIDTH - 1),
		22644 => to_unsigned(27041, LUT_AMPL_WIDTH - 1),
		22645 => to_unsigned(27039, LUT_AMPL_WIDTH - 1),
		22646 => to_unsigned(27037, LUT_AMPL_WIDTH - 1),
		22647 => to_unsigned(27035, LUT_AMPL_WIDTH - 1),
		22648 => to_unsigned(27034, LUT_AMPL_WIDTH - 1),
		22649 => to_unsigned(27032, LUT_AMPL_WIDTH - 1),
		22650 => to_unsigned(27030, LUT_AMPL_WIDTH - 1),
		22651 => to_unsigned(27028, LUT_AMPL_WIDTH - 1),
		22652 => to_unsigned(27026, LUT_AMPL_WIDTH - 1),
		22653 => to_unsigned(27025, LUT_AMPL_WIDTH - 1),
		22654 => to_unsigned(27023, LUT_AMPL_WIDTH - 1),
		22655 => to_unsigned(27021, LUT_AMPL_WIDTH - 1),
		22656 => to_unsigned(27019, LUT_AMPL_WIDTH - 1),
		22657 => to_unsigned(27018, LUT_AMPL_WIDTH - 1),
		22658 => to_unsigned(27016, LUT_AMPL_WIDTH - 1),
		22659 => to_unsigned(27014, LUT_AMPL_WIDTH - 1),
		22660 => to_unsigned(27012, LUT_AMPL_WIDTH - 1),
		22661 => to_unsigned(27010, LUT_AMPL_WIDTH - 1),
		22662 => to_unsigned(27009, LUT_AMPL_WIDTH - 1),
		22663 => to_unsigned(27007, LUT_AMPL_WIDTH - 1),
		22664 => to_unsigned(27005, LUT_AMPL_WIDTH - 1),
		22665 => to_unsigned(27003, LUT_AMPL_WIDTH - 1),
		22666 => to_unsigned(27002, LUT_AMPL_WIDTH - 1),
		22667 => to_unsigned(27000, LUT_AMPL_WIDTH - 1),
		22668 => to_unsigned(26998, LUT_AMPL_WIDTH - 1),
		22669 => to_unsigned(26996, LUT_AMPL_WIDTH - 1),
		22670 => to_unsigned(26994, LUT_AMPL_WIDTH - 1),
		22671 => to_unsigned(26993, LUT_AMPL_WIDTH - 1),
		22672 => to_unsigned(26991, LUT_AMPL_WIDTH - 1),
		22673 => to_unsigned(26989, LUT_AMPL_WIDTH - 1),
		22674 => to_unsigned(26987, LUT_AMPL_WIDTH - 1),
		22675 => to_unsigned(26986, LUT_AMPL_WIDTH - 1),
		22676 => to_unsigned(26984, LUT_AMPL_WIDTH - 1),
		22677 => to_unsigned(26982, LUT_AMPL_WIDTH - 1),
		22678 => to_unsigned(26980, LUT_AMPL_WIDTH - 1),
		22679 => to_unsigned(26978, LUT_AMPL_WIDTH - 1),
		22680 => to_unsigned(26977, LUT_AMPL_WIDTH - 1),
		22681 => to_unsigned(26975, LUT_AMPL_WIDTH - 1),
		22682 => to_unsigned(26973, LUT_AMPL_WIDTH - 1),
		22683 => to_unsigned(26971, LUT_AMPL_WIDTH - 1),
		22684 => to_unsigned(26969, LUT_AMPL_WIDTH - 1),
		22685 => to_unsigned(26968, LUT_AMPL_WIDTH - 1),
		22686 => to_unsigned(26966, LUT_AMPL_WIDTH - 1),
		22687 => to_unsigned(26964, LUT_AMPL_WIDTH - 1),
		22688 => to_unsigned(26962, LUT_AMPL_WIDTH - 1),
		22689 => to_unsigned(26961, LUT_AMPL_WIDTH - 1),
		22690 => to_unsigned(26959, LUT_AMPL_WIDTH - 1),
		22691 => to_unsigned(26957, LUT_AMPL_WIDTH - 1),
		22692 => to_unsigned(26955, LUT_AMPL_WIDTH - 1),
		22693 => to_unsigned(26953, LUT_AMPL_WIDTH - 1),
		22694 => to_unsigned(26952, LUT_AMPL_WIDTH - 1),
		22695 => to_unsigned(26950, LUT_AMPL_WIDTH - 1),
		22696 => to_unsigned(26948, LUT_AMPL_WIDTH - 1),
		22697 => to_unsigned(26946, LUT_AMPL_WIDTH - 1),
		22698 => to_unsigned(26944, LUT_AMPL_WIDTH - 1),
		22699 => to_unsigned(26943, LUT_AMPL_WIDTH - 1),
		22700 => to_unsigned(26941, LUT_AMPL_WIDTH - 1),
		22701 => to_unsigned(26939, LUT_AMPL_WIDTH - 1),
		22702 => to_unsigned(26937, LUT_AMPL_WIDTH - 1),
		22703 => to_unsigned(26936, LUT_AMPL_WIDTH - 1),
		22704 => to_unsigned(26934, LUT_AMPL_WIDTH - 1),
		22705 => to_unsigned(26932, LUT_AMPL_WIDTH - 1),
		22706 => to_unsigned(26930, LUT_AMPL_WIDTH - 1),
		22707 => to_unsigned(26928, LUT_AMPL_WIDTH - 1),
		22708 => to_unsigned(26927, LUT_AMPL_WIDTH - 1),
		22709 => to_unsigned(26925, LUT_AMPL_WIDTH - 1),
		22710 => to_unsigned(26923, LUT_AMPL_WIDTH - 1),
		22711 => to_unsigned(26921, LUT_AMPL_WIDTH - 1),
		22712 => to_unsigned(26919, LUT_AMPL_WIDTH - 1),
		22713 => to_unsigned(26918, LUT_AMPL_WIDTH - 1),
		22714 => to_unsigned(26916, LUT_AMPL_WIDTH - 1),
		22715 => to_unsigned(26914, LUT_AMPL_WIDTH - 1),
		22716 => to_unsigned(26912, LUT_AMPL_WIDTH - 1),
		22717 => to_unsigned(26910, LUT_AMPL_WIDTH - 1),
		22718 => to_unsigned(26909, LUT_AMPL_WIDTH - 1),
		22719 => to_unsigned(26907, LUT_AMPL_WIDTH - 1),
		22720 => to_unsigned(26905, LUT_AMPL_WIDTH - 1),
		22721 => to_unsigned(26903, LUT_AMPL_WIDTH - 1),
		22722 => to_unsigned(26901, LUT_AMPL_WIDTH - 1),
		22723 => to_unsigned(26900, LUT_AMPL_WIDTH - 1),
		22724 => to_unsigned(26898, LUT_AMPL_WIDTH - 1),
		22725 => to_unsigned(26896, LUT_AMPL_WIDTH - 1),
		22726 => to_unsigned(26894, LUT_AMPL_WIDTH - 1),
		22727 => to_unsigned(26893, LUT_AMPL_WIDTH - 1),
		22728 => to_unsigned(26891, LUT_AMPL_WIDTH - 1),
		22729 => to_unsigned(26889, LUT_AMPL_WIDTH - 1),
		22730 => to_unsigned(26887, LUT_AMPL_WIDTH - 1),
		22731 => to_unsigned(26885, LUT_AMPL_WIDTH - 1),
		22732 => to_unsigned(26884, LUT_AMPL_WIDTH - 1),
		22733 => to_unsigned(26882, LUT_AMPL_WIDTH - 1),
		22734 => to_unsigned(26880, LUT_AMPL_WIDTH - 1),
		22735 => to_unsigned(26878, LUT_AMPL_WIDTH - 1),
		22736 => to_unsigned(26876, LUT_AMPL_WIDTH - 1),
		22737 => to_unsigned(26875, LUT_AMPL_WIDTH - 1),
		22738 => to_unsigned(26873, LUT_AMPL_WIDTH - 1),
		22739 => to_unsigned(26871, LUT_AMPL_WIDTH - 1),
		22740 => to_unsigned(26869, LUT_AMPL_WIDTH - 1),
		22741 => to_unsigned(26867, LUT_AMPL_WIDTH - 1),
		22742 => to_unsigned(26866, LUT_AMPL_WIDTH - 1),
		22743 => to_unsigned(26864, LUT_AMPL_WIDTH - 1),
		22744 => to_unsigned(26862, LUT_AMPL_WIDTH - 1),
		22745 => to_unsigned(26860, LUT_AMPL_WIDTH - 1),
		22746 => to_unsigned(26858, LUT_AMPL_WIDTH - 1),
		22747 => to_unsigned(26857, LUT_AMPL_WIDTH - 1),
		22748 => to_unsigned(26855, LUT_AMPL_WIDTH - 1),
		22749 => to_unsigned(26853, LUT_AMPL_WIDTH - 1),
		22750 => to_unsigned(26851, LUT_AMPL_WIDTH - 1),
		22751 => to_unsigned(26849, LUT_AMPL_WIDTH - 1),
		22752 => to_unsigned(26848, LUT_AMPL_WIDTH - 1),
		22753 => to_unsigned(26846, LUT_AMPL_WIDTH - 1),
		22754 => to_unsigned(26844, LUT_AMPL_WIDTH - 1),
		22755 => to_unsigned(26842, LUT_AMPL_WIDTH - 1),
		22756 => to_unsigned(26840, LUT_AMPL_WIDTH - 1),
		22757 => to_unsigned(26839, LUT_AMPL_WIDTH - 1),
		22758 => to_unsigned(26837, LUT_AMPL_WIDTH - 1),
		22759 => to_unsigned(26835, LUT_AMPL_WIDTH - 1),
		22760 => to_unsigned(26833, LUT_AMPL_WIDTH - 1),
		22761 => to_unsigned(26831, LUT_AMPL_WIDTH - 1),
		22762 => to_unsigned(26830, LUT_AMPL_WIDTH - 1),
		22763 => to_unsigned(26828, LUT_AMPL_WIDTH - 1),
		22764 => to_unsigned(26826, LUT_AMPL_WIDTH - 1),
		22765 => to_unsigned(26824, LUT_AMPL_WIDTH - 1),
		22766 => to_unsigned(26822, LUT_AMPL_WIDTH - 1),
		22767 => to_unsigned(26821, LUT_AMPL_WIDTH - 1),
		22768 => to_unsigned(26819, LUT_AMPL_WIDTH - 1),
		22769 => to_unsigned(26817, LUT_AMPL_WIDTH - 1),
		22770 => to_unsigned(26815, LUT_AMPL_WIDTH - 1),
		22771 => to_unsigned(26813, LUT_AMPL_WIDTH - 1),
		22772 => to_unsigned(26811, LUT_AMPL_WIDTH - 1),
		22773 => to_unsigned(26810, LUT_AMPL_WIDTH - 1),
		22774 => to_unsigned(26808, LUT_AMPL_WIDTH - 1),
		22775 => to_unsigned(26806, LUT_AMPL_WIDTH - 1),
		22776 => to_unsigned(26804, LUT_AMPL_WIDTH - 1),
		22777 => to_unsigned(26802, LUT_AMPL_WIDTH - 1),
		22778 => to_unsigned(26801, LUT_AMPL_WIDTH - 1),
		22779 => to_unsigned(26799, LUT_AMPL_WIDTH - 1),
		22780 => to_unsigned(26797, LUT_AMPL_WIDTH - 1),
		22781 => to_unsigned(26795, LUT_AMPL_WIDTH - 1),
		22782 => to_unsigned(26793, LUT_AMPL_WIDTH - 1),
		22783 => to_unsigned(26792, LUT_AMPL_WIDTH - 1),
		22784 => to_unsigned(26790, LUT_AMPL_WIDTH - 1),
		22785 => to_unsigned(26788, LUT_AMPL_WIDTH - 1),
		22786 => to_unsigned(26786, LUT_AMPL_WIDTH - 1),
		22787 => to_unsigned(26784, LUT_AMPL_WIDTH - 1),
		22788 => to_unsigned(26783, LUT_AMPL_WIDTH - 1),
		22789 => to_unsigned(26781, LUT_AMPL_WIDTH - 1),
		22790 => to_unsigned(26779, LUT_AMPL_WIDTH - 1),
		22791 => to_unsigned(26777, LUT_AMPL_WIDTH - 1),
		22792 => to_unsigned(26775, LUT_AMPL_WIDTH - 1),
		22793 => to_unsigned(26774, LUT_AMPL_WIDTH - 1),
		22794 => to_unsigned(26772, LUT_AMPL_WIDTH - 1),
		22795 => to_unsigned(26770, LUT_AMPL_WIDTH - 1),
		22796 => to_unsigned(26768, LUT_AMPL_WIDTH - 1),
		22797 => to_unsigned(26766, LUT_AMPL_WIDTH - 1),
		22798 => to_unsigned(26764, LUT_AMPL_WIDTH - 1),
		22799 => to_unsigned(26763, LUT_AMPL_WIDTH - 1),
		22800 => to_unsigned(26761, LUT_AMPL_WIDTH - 1),
		22801 => to_unsigned(26759, LUT_AMPL_WIDTH - 1),
		22802 => to_unsigned(26757, LUT_AMPL_WIDTH - 1),
		22803 => to_unsigned(26755, LUT_AMPL_WIDTH - 1),
		22804 => to_unsigned(26754, LUT_AMPL_WIDTH - 1),
		22805 => to_unsigned(26752, LUT_AMPL_WIDTH - 1),
		22806 => to_unsigned(26750, LUT_AMPL_WIDTH - 1),
		22807 => to_unsigned(26748, LUT_AMPL_WIDTH - 1),
		22808 => to_unsigned(26746, LUT_AMPL_WIDTH - 1),
		22809 => to_unsigned(26745, LUT_AMPL_WIDTH - 1),
		22810 => to_unsigned(26743, LUT_AMPL_WIDTH - 1),
		22811 => to_unsigned(26741, LUT_AMPL_WIDTH - 1),
		22812 => to_unsigned(26739, LUT_AMPL_WIDTH - 1),
		22813 => to_unsigned(26737, LUT_AMPL_WIDTH - 1),
		22814 => to_unsigned(26735, LUT_AMPL_WIDTH - 1),
		22815 => to_unsigned(26734, LUT_AMPL_WIDTH - 1),
		22816 => to_unsigned(26732, LUT_AMPL_WIDTH - 1),
		22817 => to_unsigned(26730, LUT_AMPL_WIDTH - 1),
		22818 => to_unsigned(26728, LUT_AMPL_WIDTH - 1),
		22819 => to_unsigned(26726, LUT_AMPL_WIDTH - 1),
		22820 => to_unsigned(26725, LUT_AMPL_WIDTH - 1),
		22821 => to_unsigned(26723, LUT_AMPL_WIDTH - 1),
		22822 => to_unsigned(26721, LUT_AMPL_WIDTH - 1),
		22823 => to_unsigned(26719, LUT_AMPL_WIDTH - 1),
		22824 => to_unsigned(26717, LUT_AMPL_WIDTH - 1),
		22825 => to_unsigned(26715, LUT_AMPL_WIDTH - 1),
		22826 => to_unsigned(26714, LUT_AMPL_WIDTH - 1),
		22827 => to_unsigned(26712, LUT_AMPL_WIDTH - 1),
		22828 => to_unsigned(26710, LUT_AMPL_WIDTH - 1),
		22829 => to_unsigned(26708, LUT_AMPL_WIDTH - 1),
		22830 => to_unsigned(26706, LUT_AMPL_WIDTH - 1),
		22831 => to_unsigned(26705, LUT_AMPL_WIDTH - 1),
		22832 => to_unsigned(26703, LUT_AMPL_WIDTH - 1),
		22833 => to_unsigned(26701, LUT_AMPL_WIDTH - 1),
		22834 => to_unsigned(26699, LUT_AMPL_WIDTH - 1),
		22835 => to_unsigned(26697, LUT_AMPL_WIDTH - 1),
		22836 => to_unsigned(26695, LUT_AMPL_WIDTH - 1),
		22837 => to_unsigned(26694, LUT_AMPL_WIDTH - 1),
		22838 => to_unsigned(26692, LUT_AMPL_WIDTH - 1),
		22839 => to_unsigned(26690, LUT_AMPL_WIDTH - 1),
		22840 => to_unsigned(26688, LUT_AMPL_WIDTH - 1),
		22841 => to_unsigned(26686, LUT_AMPL_WIDTH - 1),
		22842 => to_unsigned(26684, LUT_AMPL_WIDTH - 1),
		22843 => to_unsigned(26683, LUT_AMPL_WIDTH - 1),
		22844 => to_unsigned(26681, LUT_AMPL_WIDTH - 1),
		22845 => to_unsigned(26679, LUT_AMPL_WIDTH - 1),
		22846 => to_unsigned(26677, LUT_AMPL_WIDTH - 1),
		22847 => to_unsigned(26675, LUT_AMPL_WIDTH - 1),
		22848 => to_unsigned(26674, LUT_AMPL_WIDTH - 1),
		22849 => to_unsigned(26672, LUT_AMPL_WIDTH - 1),
		22850 => to_unsigned(26670, LUT_AMPL_WIDTH - 1),
		22851 => to_unsigned(26668, LUT_AMPL_WIDTH - 1),
		22852 => to_unsigned(26666, LUT_AMPL_WIDTH - 1),
		22853 => to_unsigned(26664, LUT_AMPL_WIDTH - 1),
		22854 => to_unsigned(26663, LUT_AMPL_WIDTH - 1),
		22855 => to_unsigned(26661, LUT_AMPL_WIDTH - 1),
		22856 => to_unsigned(26659, LUT_AMPL_WIDTH - 1),
		22857 => to_unsigned(26657, LUT_AMPL_WIDTH - 1),
		22858 => to_unsigned(26655, LUT_AMPL_WIDTH - 1),
		22859 => to_unsigned(26653, LUT_AMPL_WIDTH - 1),
		22860 => to_unsigned(26652, LUT_AMPL_WIDTH - 1),
		22861 => to_unsigned(26650, LUT_AMPL_WIDTH - 1),
		22862 => to_unsigned(26648, LUT_AMPL_WIDTH - 1),
		22863 => to_unsigned(26646, LUT_AMPL_WIDTH - 1),
		22864 => to_unsigned(26644, LUT_AMPL_WIDTH - 1),
		22865 => to_unsigned(26642, LUT_AMPL_WIDTH - 1),
		22866 => to_unsigned(26641, LUT_AMPL_WIDTH - 1),
		22867 => to_unsigned(26639, LUT_AMPL_WIDTH - 1),
		22868 => to_unsigned(26637, LUT_AMPL_WIDTH - 1),
		22869 => to_unsigned(26635, LUT_AMPL_WIDTH - 1),
		22870 => to_unsigned(26633, LUT_AMPL_WIDTH - 1),
		22871 => to_unsigned(26631, LUT_AMPL_WIDTH - 1),
		22872 => to_unsigned(26630, LUT_AMPL_WIDTH - 1),
		22873 => to_unsigned(26628, LUT_AMPL_WIDTH - 1),
		22874 => to_unsigned(26626, LUT_AMPL_WIDTH - 1),
		22875 => to_unsigned(26624, LUT_AMPL_WIDTH - 1),
		22876 => to_unsigned(26622, LUT_AMPL_WIDTH - 1),
		22877 => to_unsigned(26621, LUT_AMPL_WIDTH - 1),
		22878 => to_unsigned(26619, LUT_AMPL_WIDTH - 1),
		22879 => to_unsigned(26617, LUT_AMPL_WIDTH - 1),
		22880 => to_unsigned(26615, LUT_AMPL_WIDTH - 1),
		22881 => to_unsigned(26613, LUT_AMPL_WIDTH - 1),
		22882 => to_unsigned(26611, LUT_AMPL_WIDTH - 1),
		22883 => to_unsigned(26610, LUT_AMPL_WIDTH - 1),
		22884 => to_unsigned(26608, LUT_AMPL_WIDTH - 1),
		22885 => to_unsigned(26606, LUT_AMPL_WIDTH - 1),
		22886 => to_unsigned(26604, LUT_AMPL_WIDTH - 1),
		22887 => to_unsigned(26602, LUT_AMPL_WIDTH - 1),
		22888 => to_unsigned(26600, LUT_AMPL_WIDTH - 1),
		22889 => to_unsigned(26599, LUT_AMPL_WIDTH - 1),
		22890 => to_unsigned(26597, LUT_AMPL_WIDTH - 1),
		22891 => to_unsigned(26595, LUT_AMPL_WIDTH - 1),
		22892 => to_unsigned(26593, LUT_AMPL_WIDTH - 1),
		22893 => to_unsigned(26591, LUT_AMPL_WIDTH - 1),
		22894 => to_unsigned(26589, LUT_AMPL_WIDTH - 1),
		22895 => to_unsigned(26588, LUT_AMPL_WIDTH - 1),
		22896 => to_unsigned(26586, LUT_AMPL_WIDTH - 1),
		22897 => to_unsigned(26584, LUT_AMPL_WIDTH - 1),
		22898 => to_unsigned(26582, LUT_AMPL_WIDTH - 1),
		22899 => to_unsigned(26580, LUT_AMPL_WIDTH - 1),
		22900 => to_unsigned(26578, LUT_AMPL_WIDTH - 1),
		22901 => to_unsigned(26576, LUT_AMPL_WIDTH - 1),
		22902 => to_unsigned(26575, LUT_AMPL_WIDTH - 1),
		22903 => to_unsigned(26573, LUT_AMPL_WIDTH - 1),
		22904 => to_unsigned(26571, LUT_AMPL_WIDTH - 1),
		22905 => to_unsigned(26569, LUT_AMPL_WIDTH - 1),
		22906 => to_unsigned(26567, LUT_AMPL_WIDTH - 1),
		22907 => to_unsigned(26565, LUT_AMPL_WIDTH - 1),
		22908 => to_unsigned(26564, LUT_AMPL_WIDTH - 1),
		22909 => to_unsigned(26562, LUT_AMPL_WIDTH - 1),
		22910 => to_unsigned(26560, LUT_AMPL_WIDTH - 1),
		22911 => to_unsigned(26558, LUT_AMPL_WIDTH - 1),
		22912 => to_unsigned(26556, LUT_AMPL_WIDTH - 1),
		22913 => to_unsigned(26554, LUT_AMPL_WIDTH - 1),
		22914 => to_unsigned(26553, LUT_AMPL_WIDTH - 1),
		22915 => to_unsigned(26551, LUT_AMPL_WIDTH - 1),
		22916 => to_unsigned(26549, LUT_AMPL_WIDTH - 1),
		22917 => to_unsigned(26547, LUT_AMPL_WIDTH - 1),
		22918 => to_unsigned(26545, LUT_AMPL_WIDTH - 1),
		22919 => to_unsigned(26543, LUT_AMPL_WIDTH - 1),
		22920 => to_unsigned(26542, LUT_AMPL_WIDTH - 1),
		22921 => to_unsigned(26540, LUT_AMPL_WIDTH - 1),
		22922 => to_unsigned(26538, LUT_AMPL_WIDTH - 1),
		22923 => to_unsigned(26536, LUT_AMPL_WIDTH - 1),
		22924 => to_unsigned(26534, LUT_AMPL_WIDTH - 1),
		22925 => to_unsigned(26532, LUT_AMPL_WIDTH - 1),
		22926 => to_unsigned(26530, LUT_AMPL_WIDTH - 1),
		22927 => to_unsigned(26529, LUT_AMPL_WIDTH - 1),
		22928 => to_unsigned(26527, LUT_AMPL_WIDTH - 1),
		22929 => to_unsigned(26525, LUT_AMPL_WIDTH - 1),
		22930 => to_unsigned(26523, LUT_AMPL_WIDTH - 1),
		22931 => to_unsigned(26521, LUT_AMPL_WIDTH - 1),
		22932 => to_unsigned(26519, LUT_AMPL_WIDTH - 1),
		22933 => to_unsigned(26518, LUT_AMPL_WIDTH - 1),
		22934 => to_unsigned(26516, LUT_AMPL_WIDTH - 1),
		22935 => to_unsigned(26514, LUT_AMPL_WIDTH - 1),
		22936 => to_unsigned(26512, LUT_AMPL_WIDTH - 1),
		22937 => to_unsigned(26510, LUT_AMPL_WIDTH - 1),
		22938 => to_unsigned(26508, LUT_AMPL_WIDTH - 1),
		22939 => to_unsigned(26506, LUT_AMPL_WIDTH - 1),
		22940 => to_unsigned(26505, LUT_AMPL_WIDTH - 1),
		22941 => to_unsigned(26503, LUT_AMPL_WIDTH - 1),
		22942 => to_unsigned(26501, LUT_AMPL_WIDTH - 1),
		22943 => to_unsigned(26499, LUT_AMPL_WIDTH - 1),
		22944 => to_unsigned(26497, LUT_AMPL_WIDTH - 1),
		22945 => to_unsigned(26495, LUT_AMPL_WIDTH - 1),
		22946 => to_unsigned(26494, LUT_AMPL_WIDTH - 1),
		22947 => to_unsigned(26492, LUT_AMPL_WIDTH - 1),
		22948 => to_unsigned(26490, LUT_AMPL_WIDTH - 1),
		22949 => to_unsigned(26488, LUT_AMPL_WIDTH - 1),
		22950 => to_unsigned(26486, LUT_AMPL_WIDTH - 1),
		22951 => to_unsigned(26484, LUT_AMPL_WIDTH - 1),
		22952 => to_unsigned(26482, LUT_AMPL_WIDTH - 1),
		22953 => to_unsigned(26481, LUT_AMPL_WIDTH - 1),
		22954 => to_unsigned(26479, LUT_AMPL_WIDTH - 1),
		22955 => to_unsigned(26477, LUT_AMPL_WIDTH - 1),
		22956 => to_unsigned(26475, LUT_AMPL_WIDTH - 1),
		22957 => to_unsigned(26473, LUT_AMPL_WIDTH - 1),
		22958 => to_unsigned(26471, LUT_AMPL_WIDTH - 1),
		22959 => to_unsigned(26469, LUT_AMPL_WIDTH - 1),
		22960 => to_unsigned(26468, LUT_AMPL_WIDTH - 1),
		22961 => to_unsigned(26466, LUT_AMPL_WIDTH - 1),
		22962 => to_unsigned(26464, LUT_AMPL_WIDTH - 1),
		22963 => to_unsigned(26462, LUT_AMPL_WIDTH - 1),
		22964 => to_unsigned(26460, LUT_AMPL_WIDTH - 1),
		22965 => to_unsigned(26458, LUT_AMPL_WIDTH - 1),
		22966 => to_unsigned(26457, LUT_AMPL_WIDTH - 1),
		22967 => to_unsigned(26455, LUT_AMPL_WIDTH - 1),
		22968 => to_unsigned(26453, LUT_AMPL_WIDTH - 1),
		22969 => to_unsigned(26451, LUT_AMPL_WIDTH - 1),
		22970 => to_unsigned(26449, LUT_AMPL_WIDTH - 1),
		22971 => to_unsigned(26447, LUT_AMPL_WIDTH - 1),
		22972 => to_unsigned(26445, LUT_AMPL_WIDTH - 1),
		22973 => to_unsigned(26444, LUT_AMPL_WIDTH - 1),
		22974 => to_unsigned(26442, LUT_AMPL_WIDTH - 1),
		22975 => to_unsigned(26440, LUT_AMPL_WIDTH - 1),
		22976 => to_unsigned(26438, LUT_AMPL_WIDTH - 1),
		22977 => to_unsigned(26436, LUT_AMPL_WIDTH - 1),
		22978 => to_unsigned(26434, LUT_AMPL_WIDTH - 1),
		22979 => to_unsigned(26432, LUT_AMPL_WIDTH - 1),
		22980 => to_unsigned(26431, LUT_AMPL_WIDTH - 1),
		22981 => to_unsigned(26429, LUT_AMPL_WIDTH - 1),
		22982 => to_unsigned(26427, LUT_AMPL_WIDTH - 1),
		22983 => to_unsigned(26425, LUT_AMPL_WIDTH - 1),
		22984 => to_unsigned(26423, LUT_AMPL_WIDTH - 1),
		22985 => to_unsigned(26421, LUT_AMPL_WIDTH - 1),
		22986 => to_unsigned(26419, LUT_AMPL_WIDTH - 1),
		22987 => to_unsigned(26418, LUT_AMPL_WIDTH - 1),
		22988 => to_unsigned(26416, LUT_AMPL_WIDTH - 1),
		22989 => to_unsigned(26414, LUT_AMPL_WIDTH - 1),
		22990 => to_unsigned(26412, LUT_AMPL_WIDTH - 1),
		22991 => to_unsigned(26410, LUT_AMPL_WIDTH - 1),
		22992 => to_unsigned(26408, LUT_AMPL_WIDTH - 1),
		22993 => to_unsigned(26406, LUT_AMPL_WIDTH - 1),
		22994 => to_unsigned(26405, LUT_AMPL_WIDTH - 1),
		22995 => to_unsigned(26403, LUT_AMPL_WIDTH - 1),
		22996 => to_unsigned(26401, LUT_AMPL_WIDTH - 1),
		22997 => to_unsigned(26399, LUT_AMPL_WIDTH - 1),
		22998 => to_unsigned(26397, LUT_AMPL_WIDTH - 1),
		22999 => to_unsigned(26395, LUT_AMPL_WIDTH - 1),
		23000 => to_unsigned(26393, LUT_AMPL_WIDTH - 1),
		23001 => to_unsigned(26392, LUT_AMPL_WIDTH - 1),
		23002 => to_unsigned(26390, LUT_AMPL_WIDTH - 1),
		23003 => to_unsigned(26388, LUT_AMPL_WIDTH - 1),
		23004 => to_unsigned(26386, LUT_AMPL_WIDTH - 1),
		23005 => to_unsigned(26384, LUT_AMPL_WIDTH - 1),
		23006 => to_unsigned(26382, LUT_AMPL_WIDTH - 1),
		23007 => to_unsigned(26380, LUT_AMPL_WIDTH - 1),
		23008 => to_unsigned(26378, LUT_AMPL_WIDTH - 1),
		23009 => to_unsigned(26377, LUT_AMPL_WIDTH - 1),
		23010 => to_unsigned(26375, LUT_AMPL_WIDTH - 1),
		23011 => to_unsigned(26373, LUT_AMPL_WIDTH - 1),
		23012 => to_unsigned(26371, LUT_AMPL_WIDTH - 1),
		23013 => to_unsigned(26369, LUT_AMPL_WIDTH - 1),
		23014 => to_unsigned(26367, LUT_AMPL_WIDTH - 1),
		23015 => to_unsigned(26365, LUT_AMPL_WIDTH - 1),
		23016 => to_unsigned(26364, LUT_AMPL_WIDTH - 1),
		23017 => to_unsigned(26362, LUT_AMPL_WIDTH - 1),
		23018 => to_unsigned(26360, LUT_AMPL_WIDTH - 1),
		23019 => to_unsigned(26358, LUT_AMPL_WIDTH - 1),
		23020 => to_unsigned(26356, LUT_AMPL_WIDTH - 1),
		23021 => to_unsigned(26354, LUT_AMPL_WIDTH - 1),
		23022 => to_unsigned(26352, LUT_AMPL_WIDTH - 1),
		23023 => to_unsigned(26350, LUT_AMPL_WIDTH - 1),
		23024 => to_unsigned(26349, LUT_AMPL_WIDTH - 1),
		23025 => to_unsigned(26347, LUT_AMPL_WIDTH - 1),
		23026 => to_unsigned(26345, LUT_AMPL_WIDTH - 1),
		23027 => to_unsigned(26343, LUT_AMPL_WIDTH - 1),
		23028 => to_unsigned(26341, LUT_AMPL_WIDTH - 1),
		23029 => to_unsigned(26339, LUT_AMPL_WIDTH - 1),
		23030 => to_unsigned(26337, LUT_AMPL_WIDTH - 1),
		23031 => to_unsigned(26336, LUT_AMPL_WIDTH - 1),
		23032 => to_unsigned(26334, LUT_AMPL_WIDTH - 1),
		23033 => to_unsigned(26332, LUT_AMPL_WIDTH - 1),
		23034 => to_unsigned(26330, LUT_AMPL_WIDTH - 1),
		23035 => to_unsigned(26328, LUT_AMPL_WIDTH - 1),
		23036 => to_unsigned(26326, LUT_AMPL_WIDTH - 1),
		23037 => to_unsigned(26324, LUT_AMPL_WIDTH - 1),
		23038 => to_unsigned(26322, LUT_AMPL_WIDTH - 1),
		23039 => to_unsigned(26321, LUT_AMPL_WIDTH - 1),
		23040 => to_unsigned(26319, LUT_AMPL_WIDTH - 1),
		23041 => to_unsigned(26317, LUT_AMPL_WIDTH - 1),
		23042 => to_unsigned(26315, LUT_AMPL_WIDTH - 1),
		23043 => to_unsigned(26313, LUT_AMPL_WIDTH - 1),
		23044 => to_unsigned(26311, LUT_AMPL_WIDTH - 1),
		23045 => to_unsigned(26309, LUT_AMPL_WIDTH - 1),
		23046 => to_unsigned(26307, LUT_AMPL_WIDTH - 1),
		23047 => to_unsigned(26306, LUT_AMPL_WIDTH - 1),
		23048 => to_unsigned(26304, LUT_AMPL_WIDTH - 1),
		23049 => to_unsigned(26302, LUT_AMPL_WIDTH - 1),
		23050 => to_unsigned(26300, LUT_AMPL_WIDTH - 1),
		23051 => to_unsigned(26298, LUT_AMPL_WIDTH - 1),
		23052 => to_unsigned(26296, LUT_AMPL_WIDTH - 1),
		23053 => to_unsigned(26294, LUT_AMPL_WIDTH - 1),
		23054 => to_unsigned(26292, LUT_AMPL_WIDTH - 1),
		23055 => to_unsigned(26291, LUT_AMPL_WIDTH - 1),
		23056 => to_unsigned(26289, LUT_AMPL_WIDTH - 1),
		23057 => to_unsigned(26287, LUT_AMPL_WIDTH - 1),
		23058 => to_unsigned(26285, LUT_AMPL_WIDTH - 1),
		23059 => to_unsigned(26283, LUT_AMPL_WIDTH - 1),
		23060 => to_unsigned(26281, LUT_AMPL_WIDTH - 1),
		23061 => to_unsigned(26279, LUT_AMPL_WIDTH - 1),
		23062 => to_unsigned(26277, LUT_AMPL_WIDTH - 1),
		23063 => to_unsigned(26276, LUT_AMPL_WIDTH - 1),
		23064 => to_unsigned(26274, LUT_AMPL_WIDTH - 1),
		23065 => to_unsigned(26272, LUT_AMPL_WIDTH - 1),
		23066 => to_unsigned(26270, LUT_AMPL_WIDTH - 1),
		23067 => to_unsigned(26268, LUT_AMPL_WIDTH - 1),
		23068 => to_unsigned(26266, LUT_AMPL_WIDTH - 1),
		23069 => to_unsigned(26264, LUT_AMPL_WIDTH - 1),
		23070 => to_unsigned(26262, LUT_AMPL_WIDTH - 1),
		23071 => to_unsigned(26261, LUT_AMPL_WIDTH - 1),
		23072 => to_unsigned(26259, LUT_AMPL_WIDTH - 1),
		23073 => to_unsigned(26257, LUT_AMPL_WIDTH - 1),
		23074 => to_unsigned(26255, LUT_AMPL_WIDTH - 1),
		23075 => to_unsigned(26253, LUT_AMPL_WIDTH - 1),
		23076 => to_unsigned(26251, LUT_AMPL_WIDTH - 1),
		23077 => to_unsigned(26249, LUT_AMPL_WIDTH - 1),
		23078 => to_unsigned(26247, LUT_AMPL_WIDTH - 1),
		23079 => to_unsigned(26246, LUT_AMPL_WIDTH - 1),
		23080 => to_unsigned(26244, LUT_AMPL_WIDTH - 1),
		23081 => to_unsigned(26242, LUT_AMPL_WIDTH - 1),
		23082 => to_unsigned(26240, LUT_AMPL_WIDTH - 1),
		23083 => to_unsigned(26238, LUT_AMPL_WIDTH - 1),
		23084 => to_unsigned(26236, LUT_AMPL_WIDTH - 1),
		23085 => to_unsigned(26234, LUT_AMPL_WIDTH - 1),
		23086 => to_unsigned(26232, LUT_AMPL_WIDTH - 1),
		23087 => to_unsigned(26230, LUT_AMPL_WIDTH - 1),
		23088 => to_unsigned(26229, LUT_AMPL_WIDTH - 1),
		23089 => to_unsigned(26227, LUT_AMPL_WIDTH - 1),
		23090 => to_unsigned(26225, LUT_AMPL_WIDTH - 1),
		23091 => to_unsigned(26223, LUT_AMPL_WIDTH - 1),
		23092 => to_unsigned(26221, LUT_AMPL_WIDTH - 1),
		23093 => to_unsigned(26219, LUT_AMPL_WIDTH - 1),
		23094 => to_unsigned(26217, LUT_AMPL_WIDTH - 1),
		23095 => to_unsigned(26215, LUT_AMPL_WIDTH - 1),
		23096 => to_unsigned(26214, LUT_AMPL_WIDTH - 1),
		23097 => to_unsigned(26212, LUT_AMPL_WIDTH - 1),
		23098 => to_unsigned(26210, LUT_AMPL_WIDTH - 1),
		23099 => to_unsigned(26208, LUT_AMPL_WIDTH - 1),
		23100 => to_unsigned(26206, LUT_AMPL_WIDTH - 1),
		23101 => to_unsigned(26204, LUT_AMPL_WIDTH - 1),
		23102 => to_unsigned(26202, LUT_AMPL_WIDTH - 1),
		23103 => to_unsigned(26200, LUT_AMPL_WIDTH - 1),
		23104 => to_unsigned(26198, LUT_AMPL_WIDTH - 1),
		23105 => to_unsigned(26197, LUT_AMPL_WIDTH - 1),
		23106 => to_unsigned(26195, LUT_AMPL_WIDTH - 1),
		23107 => to_unsigned(26193, LUT_AMPL_WIDTH - 1),
		23108 => to_unsigned(26191, LUT_AMPL_WIDTH - 1),
		23109 => to_unsigned(26189, LUT_AMPL_WIDTH - 1),
		23110 => to_unsigned(26187, LUT_AMPL_WIDTH - 1),
		23111 => to_unsigned(26185, LUT_AMPL_WIDTH - 1),
		23112 => to_unsigned(26183, LUT_AMPL_WIDTH - 1),
		23113 => to_unsigned(26181, LUT_AMPL_WIDTH - 1),
		23114 => to_unsigned(26180, LUT_AMPL_WIDTH - 1),
		23115 => to_unsigned(26178, LUT_AMPL_WIDTH - 1),
		23116 => to_unsigned(26176, LUT_AMPL_WIDTH - 1),
		23117 => to_unsigned(26174, LUT_AMPL_WIDTH - 1),
		23118 => to_unsigned(26172, LUT_AMPL_WIDTH - 1),
		23119 => to_unsigned(26170, LUT_AMPL_WIDTH - 1),
		23120 => to_unsigned(26168, LUT_AMPL_WIDTH - 1),
		23121 => to_unsigned(26166, LUT_AMPL_WIDTH - 1),
		23122 => to_unsigned(26164, LUT_AMPL_WIDTH - 1),
		23123 => to_unsigned(26163, LUT_AMPL_WIDTH - 1),
		23124 => to_unsigned(26161, LUT_AMPL_WIDTH - 1),
		23125 => to_unsigned(26159, LUT_AMPL_WIDTH - 1),
		23126 => to_unsigned(26157, LUT_AMPL_WIDTH - 1),
		23127 => to_unsigned(26155, LUT_AMPL_WIDTH - 1),
		23128 => to_unsigned(26153, LUT_AMPL_WIDTH - 1),
		23129 => to_unsigned(26151, LUT_AMPL_WIDTH - 1),
		23130 => to_unsigned(26149, LUT_AMPL_WIDTH - 1),
		23131 => to_unsigned(26147, LUT_AMPL_WIDTH - 1),
		23132 => to_unsigned(26146, LUT_AMPL_WIDTH - 1),
		23133 => to_unsigned(26144, LUT_AMPL_WIDTH - 1),
		23134 => to_unsigned(26142, LUT_AMPL_WIDTH - 1),
		23135 => to_unsigned(26140, LUT_AMPL_WIDTH - 1),
		23136 => to_unsigned(26138, LUT_AMPL_WIDTH - 1),
		23137 => to_unsigned(26136, LUT_AMPL_WIDTH - 1),
		23138 => to_unsigned(26134, LUT_AMPL_WIDTH - 1),
		23139 => to_unsigned(26132, LUT_AMPL_WIDTH - 1),
		23140 => to_unsigned(26130, LUT_AMPL_WIDTH - 1),
		23141 => to_unsigned(26128, LUT_AMPL_WIDTH - 1),
		23142 => to_unsigned(26127, LUT_AMPL_WIDTH - 1),
		23143 => to_unsigned(26125, LUT_AMPL_WIDTH - 1),
		23144 => to_unsigned(26123, LUT_AMPL_WIDTH - 1),
		23145 => to_unsigned(26121, LUT_AMPL_WIDTH - 1),
		23146 => to_unsigned(26119, LUT_AMPL_WIDTH - 1),
		23147 => to_unsigned(26117, LUT_AMPL_WIDTH - 1),
		23148 => to_unsigned(26115, LUT_AMPL_WIDTH - 1),
		23149 => to_unsigned(26113, LUT_AMPL_WIDTH - 1),
		23150 => to_unsigned(26111, LUT_AMPL_WIDTH - 1),
		23151 => to_unsigned(26109, LUT_AMPL_WIDTH - 1),
		23152 => to_unsigned(26108, LUT_AMPL_WIDTH - 1),
		23153 => to_unsigned(26106, LUT_AMPL_WIDTH - 1),
		23154 => to_unsigned(26104, LUT_AMPL_WIDTH - 1),
		23155 => to_unsigned(26102, LUT_AMPL_WIDTH - 1),
		23156 => to_unsigned(26100, LUT_AMPL_WIDTH - 1),
		23157 => to_unsigned(26098, LUT_AMPL_WIDTH - 1),
		23158 => to_unsigned(26096, LUT_AMPL_WIDTH - 1),
		23159 => to_unsigned(26094, LUT_AMPL_WIDTH - 1),
		23160 => to_unsigned(26092, LUT_AMPL_WIDTH - 1),
		23161 => to_unsigned(26090, LUT_AMPL_WIDTH - 1),
		23162 => to_unsigned(26089, LUT_AMPL_WIDTH - 1),
		23163 => to_unsigned(26087, LUT_AMPL_WIDTH - 1),
		23164 => to_unsigned(26085, LUT_AMPL_WIDTH - 1),
		23165 => to_unsigned(26083, LUT_AMPL_WIDTH - 1),
		23166 => to_unsigned(26081, LUT_AMPL_WIDTH - 1),
		23167 => to_unsigned(26079, LUT_AMPL_WIDTH - 1),
		23168 => to_unsigned(26077, LUT_AMPL_WIDTH - 1),
		23169 => to_unsigned(26075, LUT_AMPL_WIDTH - 1),
		23170 => to_unsigned(26073, LUT_AMPL_WIDTH - 1),
		23171 => to_unsigned(26071, LUT_AMPL_WIDTH - 1),
		23172 => to_unsigned(26070, LUT_AMPL_WIDTH - 1),
		23173 => to_unsigned(26068, LUT_AMPL_WIDTH - 1),
		23174 => to_unsigned(26066, LUT_AMPL_WIDTH - 1),
		23175 => to_unsigned(26064, LUT_AMPL_WIDTH - 1),
		23176 => to_unsigned(26062, LUT_AMPL_WIDTH - 1),
		23177 => to_unsigned(26060, LUT_AMPL_WIDTH - 1),
		23178 => to_unsigned(26058, LUT_AMPL_WIDTH - 1),
		23179 => to_unsigned(26056, LUT_AMPL_WIDTH - 1),
		23180 => to_unsigned(26054, LUT_AMPL_WIDTH - 1),
		23181 => to_unsigned(26052, LUT_AMPL_WIDTH - 1),
		23182 => to_unsigned(26051, LUT_AMPL_WIDTH - 1),
		23183 => to_unsigned(26049, LUT_AMPL_WIDTH - 1),
		23184 => to_unsigned(26047, LUT_AMPL_WIDTH - 1),
		23185 => to_unsigned(26045, LUT_AMPL_WIDTH - 1),
		23186 => to_unsigned(26043, LUT_AMPL_WIDTH - 1),
		23187 => to_unsigned(26041, LUT_AMPL_WIDTH - 1),
		23188 => to_unsigned(26039, LUT_AMPL_WIDTH - 1),
		23189 => to_unsigned(26037, LUT_AMPL_WIDTH - 1),
		23190 => to_unsigned(26035, LUT_AMPL_WIDTH - 1),
		23191 => to_unsigned(26033, LUT_AMPL_WIDTH - 1),
		23192 => to_unsigned(26031, LUT_AMPL_WIDTH - 1),
		23193 => to_unsigned(26030, LUT_AMPL_WIDTH - 1),
		23194 => to_unsigned(26028, LUT_AMPL_WIDTH - 1),
		23195 => to_unsigned(26026, LUT_AMPL_WIDTH - 1),
		23196 => to_unsigned(26024, LUT_AMPL_WIDTH - 1),
		23197 => to_unsigned(26022, LUT_AMPL_WIDTH - 1),
		23198 => to_unsigned(26020, LUT_AMPL_WIDTH - 1),
		23199 => to_unsigned(26018, LUT_AMPL_WIDTH - 1),
		23200 => to_unsigned(26016, LUT_AMPL_WIDTH - 1),
		23201 => to_unsigned(26014, LUT_AMPL_WIDTH - 1),
		23202 => to_unsigned(26012, LUT_AMPL_WIDTH - 1),
		23203 => to_unsigned(26010, LUT_AMPL_WIDTH - 1),
		23204 => to_unsigned(26009, LUT_AMPL_WIDTH - 1),
		23205 => to_unsigned(26007, LUT_AMPL_WIDTH - 1),
		23206 => to_unsigned(26005, LUT_AMPL_WIDTH - 1),
		23207 => to_unsigned(26003, LUT_AMPL_WIDTH - 1),
		23208 => to_unsigned(26001, LUT_AMPL_WIDTH - 1),
		23209 => to_unsigned(25999, LUT_AMPL_WIDTH - 1),
		23210 => to_unsigned(25997, LUT_AMPL_WIDTH - 1),
		23211 => to_unsigned(25995, LUT_AMPL_WIDTH - 1),
		23212 => to_unsigned(25993, LUT_AMPL_WIDTH - 1),
		23213 => to_unsigned(25991, LUT_AMPL_WIDTH - 1),
		23214 => to_unsigned(25989, LUT_AMPL_WIDTH - 1),
		23215 => to_unsigned(25988, LUT_AMPL_WIDTH - 1),
		23216 => to_unsigned(25986, LUT_AMPL_WIDTH - 1),
		23217 => to_unsigned(25984, LUT_AMPL_WIDTH - 1),
		23218 => to_unsigned(25982, LUT_AMPL_WIDTH - 1),
		23219 => to_unsigned(25980, LUT_AMPL_WIDTH - 1),
		23220 => to_unsigned(25978, LUT_AMPL_WIDTH - 1),
		23221 => to_unsigned(25976, LUT_AMPL_WIDTH - 1),
		23222 => to_unsigned(25974, LUT_AMPL_WIDTH - 1),
		23223 => to_unsigned(25972, LUT_AMPL_WIDTH - 1),
		23224 => to_unsigned(25970, LUT_AMPL_WIDTH - 1),
		23225 => to_unsigned(25968, LUT_AMPL_WIDTH - 1),
		23226 => to_unsigned(25966, LUT_AMPL_WIDTH - 1),
		23227 => to_unsigned(25965, LUT_AMPL_WIDTH - 1),
		23228 => to_unsigned(25963, LUT_AMPL_WIDTH - 1),
		23229 => to_unsigned(25961, LUT_AMPL_WIDTH - 1),
		23230 => to_unsigned(25959, LUT_AMPL_WIDTH - 1),
		23231 => to_unsigned(25957, LUT_AMPL_WIDTH - 1),
		23232 => to_unsigned(25955, LUT_AMPL_WIDTH - 1),
		23233 => to_unsigned(25953, LUT_AMPL_WIDTH - 1),
		23234 => to_unsigned(25951, LUT_AMPL_WIDTH - 1),
		23235 => to_unsigned(25949, LUT_AMPL_WIDTH - 1),
		23236 => to_unsigned(25947, LUT_AMPL_WIDTH - 1),
		23237 => to_unsigned(25945, LUT_AMPL_WIDTH - 1),
		23238 => to_unsigned(25943, LUT_AMPL_WIDTH - 1),
		23239 => to_unsigned(25942, LUT_AMPL_WIDTH - 1),
		23240 => to_unsigned(25940, LUT_AMPL_WIDTH - 1),
		23241 => to_unsigned(25938, LUT_AMPL_WIDTH - 1),
		23242 => to_unsigned(25936, LUT_AMPL_WIDTH - 1),
		23243 => to_unsigned(25934, LUT_AMPL_WIDTH - 1),
		23244 => to_unsigned(25932, LUT_AMPL_WIDTH - 1),
		23245 => to_unsigned(25930, LUT_AMPL_WIDTH - 1),
		23246 => to_unsigned(25928, LUT_AMPL_WIDTH - 1),
		23247 => to_unsigned(25926, LUT_AMPL_WIDTH - 1),
		23248 => to_unsigned(25924, LUT_AMPL_WIDTH - 1),
		23249 => to_unsigned(25922, LUT_AMPL_WIDTH - 1),
		23250 => to_unsigned(25920, LUT_AMPL_WIDTH - 1),
		23251 => to_unsigned(25918, LUT_AMPL_WIDTH - 1),
		23252 => to_unsigned(25917, LUT_AMPL_WIDTH - 1),
		23253 => to_unsigned(25915, LUT_AMPL_WIDTH - 1),
		23254 => to_unsigned(25913, LUT_AMPL_WIDTH - 1),
		23255 => to_unsigned(25911, LUT_AMPL_WIDTH - 1),
		23256 => to_unsigned(25909, LUT_AMPL_WIDTH - 1),
		23257 => to_unsigned(25907, LUT_AMPL_WIDTH - 1),
		23258 => to_unsigned(25905, LUT_AMPL_WIDTH - 1),
		23259 => to_unsigned(25903, LUT_AMPL_WIDTH - 1),
		23260 => to_unsigned(25901, LUT_AMPL_WIDTH - 1),
		23261 => to_unsigned(25899, LUT_AMPL_WIDTH - 1),
		23262 => to_unsigned(25897, LUT_AMPL_WIDTH - 1),
		23263 => to_unsigned(25895, LUT_AMPL_WIDTH - 1),
		23264 => to_unsigned(25893, LUT_AMPL_WIDTH - 1),
		23265 => to_unsigned(25892, LUT_AMPL_WIDTH - 1),
		23266 => to_unsigned(25890, LUT_AMPL_WIDTH - 1),
		23267 => to_unsigned(25888, LUT_AMPL_WIDTH - 1),
		23268 => to_unsigned(25886, LUT_AMPL_WIDTH - 1),
		23269 => to_unsigned(25884, LUT_AMPL_WIDTH - 1),
		23270 => to_unsigned(25882, LUT_AMPL_WIDTH - 1),
		23271 => to_unsigned(25880, LUT_AMPL_WIDTH - 1),
		23272 => to_unsigned(25878, LUT_AMPL_WIDTH - 1),
		23273 => to_unsigned(25876, LUT_AMPL_WIDTH - 1),
		23274 => to_unsigned(25874, LUT_AMPL_WIDTH - 1),
		23275 => to_unsigned(25872, LUT_AMPL_WIDTH - 1),
		23276 => to_unsigned(25870, LUT_AMPL_WIDTH - 1),
		23277 => to_unsigned(25868, LUT_AMPL_WIDTH - 1),
		23278 => to_unsigned(25866, LUT_AMPL_WIDTH - 1),
		23279 => to_unsigned(25865, LUT_AMPL_WIDTH - 1),
		23280 => to_unsigned(25863, LUT_AMPL_WIDTH - 1),
		23281 => to_unsigned(25861, LUT_AMPL_WIDTH - 1),
		23282 => to_unsigned(25859, LUT_AMPL_WIDTH - 1),
		23283 => to_unsigned(25857, LUT_AMPL_WIDTH - 1),
		23284 => to_unsigned(25855, LUT_AMPL_WIDTH - 1),
		23285 => to_unsigned(25853, LUT_AMPL_WIDTH - 1),
		23286 => to_unsigned(25851, LUT_AMPL_WIDTH - 1),
		23287 => to_unsigned(25849, LUT_AMPL_WIDTH - 1),
		23288 => to_unsigned(25847, LUT_AMPL_WIDTH - 1),
		23289 => to_unsigned(25845, LUT_AMPL_WIDTH - 1),
		23290 => to_unsigned(25843, LUT_AMPL_WIDTH - 1),
		23291 => to_unsigned(25841, LUT_AMPL_WIDTH - 1),
		23292 => to_unsigned(25839, LUT_AMPL_WIDTH - 1),
		23293 => to_unsigned(25838, LUT_AMPL_WIDTH - 1),
		23294 => to_unsigned(25836, LUT_AMPL_WIDTH - 1),
		23295 => to_unsigned(25834, LUT_AMPL_WIDTH - 1),
		23296 => to_unsigned(25832, LUT_AMPL_WIDTH - 1),
		23297 => to_unsigned(25830, LUT_AMPL_WIDTH - 1),
		23298 => to_unsigned(25828, LUT_AMPL_WIDTH - 1),
		23299 => to_unsigned(25826, LUT_AMPL_WIDTH - 1),
		23300 => to_unsigned(25824, LUT_AMPL_WIDTH - 1),
		23301 => to_unsigned(25822, LUT_AMPL_WIDTH - 1),
		23302 => to_unsigned(25820, LUT_AMPL_WIDTH - 1),
		23303 => to_unsigned(25818, LUT_AMPL_WIDTH - 1),
		23304 => to_unsigned(25816, LUT_AMPL_WIDTH - 1),
		23305 => to_unsigned(25814, LUT_AMPL_WIDTH - 1),
		23306 => to_unsigned(25812, LUT_AMPL_WIDTH - 1),
		23307 => to_unsigned(25810, LUT_AMPL_WIDTH - 1),
		23308 => to_unsigned(25809, LUT_AMPL_WIDTH - 1),
		23309 => to_unsigned(25807, LUT_AMPL_WIDTH - 1),
		23310 => to_unsigned(25805, LUT_AMPL_WIDTH - 1),
		23311 => to_unsigned(25803, LUT_AMPL_WIDTH - 1),
		23312 => to_unsigned(25801, LUT_AMPL_WIDTH - 1),
		23313 => to_unsigned(25799, LUT_AMPL_WIDTH - 1),
		23314 => to_unsigned(25797, LUT_AMPL_WIDTH - 1),
		23315 => to_unsigned(25795, LUT_AMPL_WIDTH - 1),
		23316 => to_unsigned(25793, LUT_AMPL_WIDTH - 1),
		23317 => to_unsigned(25791, LUT_AMPL_WIDTH - 1),
		23318 => to_unsigned(25789, LUT_AMPL_WIDTH - 1),
		23319 => to_unsigned(25787, LUT_AMPL_WIDTH - 1),
		23320 => to_unsigned(25785, LUT_AMPL_WIDTH - 1),
		23321 => to_unsigned(25783, LUT_AMPL_WIDTH - 1),
		23322 => to_unsigned(25781, LUT_AMPL_WIDTH - 1),
		23323 => to_unsigned(25779, LUT_AMPL_WIDTH - 1),
		23324 => to_unsigned(25778, LUT_AMPL_WIDTH - 1),
		23325 => to_unsigned(25776, LUT_AMPL_WIDTH - 1),
		23326 => to_unsigned(25774, LUT_AMPL_WIDTH - 1),
		23327 => to_unsigned(25772, LUT_AMPL_WIDTH - 1),
		23328 => to_unsigned(25770, LUT_AMPL_WIDTH - 1),
		23329 => to_unsigned(25768, LUT_AMPL_WIDTH - 1),
		23330 => to_unsigned(25766, LUT_AMPL_WIDTH - 1),
		23331 => to_unsigned(25764, LUT_AMPL_WIDTH - 1),
		23332 => to_unsigned(25762, LUT_AMPL_WIDTH - 1),
		23333 => to_unsigned(25760, LUT_AMPL_WIDTH - 1),
		23334 => to_unsigned(25758, LUT_AMPL_WIDTH - 1),
		23335 => to_unsigned(25756, LUT_AMPL_WIDTH - 1),
		23336 => to_unsigned(25754, LUT_AMPL_WIDTH - 1),
		23337 => to_unsigned(25752, LUT_AMPL_WIDTH - 1),
		23338 => to_unsigned(25750, LUT_AMPL_WIDTH - 1),
		23339 => to_unsigned(25748, LUT_AMPL_WIDTH - 1),
		23340 => to_unsigned(25746, LUT_AMPL_WIDTH - 1),
		23341 => to_unsigned(25745, LUT_AMPL_WIDTH - 1),
		23342 => to_unsigned(25743, LUT_AMPL_WIDTH - 1),
		23343 => to_unsigned(25741, LUT_AMPL_WIDTH - 1),
		23344 => to_unsigned(25739, LUT_AMPL_WIDTH - 1),
		23345 => to_unsigned(25737, LUT_AMPL_WIDTH - 1),
		23346 => to_unsigned(25735, LUT_AMPL_WIDTH - 1),
		23347 => to_unsigned(25733, LUT_AMPL_WIDTH - 1),
		23348 => to_unsigned(25731, LUT_AMPL_WIDTH - 1),
		23349 => to_unsigned(25729, LUT_AMPL_WIDTH - 1),
		23350 => to_unsigned(25727, LUT_AMPL_WIDTH - 1),
		23351 => to_unsigned(25725, LUT_AMPL_WIDTH - 1),
		23352 => to_unsigned(25723, LUT_AMPL_WIDTH - 1),
		23353 => to_unsigned(25721, LUT_AMPL_WIDTH - 1),
		23354 => to_unsigned(25719, LUT_AMPL_WIDTH - 1),
		23355 => to_unsigned(25717, LUT_AMPL_WIDTH - 1),
		23356 => to_unsigned(25715, LUT_AMPL_WIDTH - 1),
		23357 => to_unsigned(25713, LUT_AMPL_WIDTH - 1),
		23358 => to_unsigned(25711, LUT_AMPL_WIDTH - 1),
		23359 => to_unsigned(25710, LUT_AMPL_WIDTH - 1),
		23360 => to_unsigned(25708, LUT_AMPL_WIDTH - 1),
		23361 => to_unsigned(25706, LUT_AMPL_WIDTH - 1),
		23362 => to_unsigned(25704, LUT_AMPL_WIDTH - 1),
		23363 => to_unsigned(25702, LUT_AMPL_WIDTH - 1),
		23364 => to_unsigned(25700, LUT_AMPL_WIDTH - 1),
		23365 => to_unsigned(25698, LUT_AMPL_WIDTH - 1),
		23366 => to_unsigned(25696, LUT_AMPL_WIDTH - 1),
		23367 => to_unsigned(25694, LUT_AMPL_WIDTH - 1),
		23368 => to_unsigned(25692, LUT_AMPL_WIDTH - 1),
		23369 => to_unsigned(25690, LUT_AMPL_WIDTH - 1),
		23370 => to_unsigned(25688, LUT_AMPL_WIDTH - 1),
		23371 => to_unsigned(25686, LUT_AMPL_WIDTH - 1),
		23372 => to_unsigned(25684, LUT_AMPL_WIDTH - 1),
		23373 => to_unsigned(25682, LUT_AMPL_WIDTH - 1),
		23374 => to_unsigned(25680, LUT_AMPL_WIDTH - 1),
		23375 => to_unsigned(25678, LUT_AMPL_WIDTH - 1),
		23376 => to_unsigned(25676, LUT_AMPL_WIDTH - 1),
		23377 => to_unsigned(25674, LUT_AMPL_WIDTH - 1),
		23378 => to_unsigned(25672, LUT_AMPL_WIDTH - 1),
		23379 => to_unsigned(25671, LUT_AMPL_WIDTH - 1),
		23380 => to_unsigned(25669, LUT_AMPL_WIDTH - 1),
		23381 => to_unsigned(25667, LUT_AMPL_WIDTH - 1),
		23382 => to_unsigned(25665, LUT_AMPL_WIDTH - 1),
		23383 => to_unsigned(25663, LUT_AMPL_WIDTH - 1),
		23384 => to_unsigned(25661, LUT_AMPL_WIDTH - 1),
		23385 => to_unsigned(25659, LUT_AMPL_WIDTH - 1),
		23386 => to_unsigned(25657, LUT_AMPL_WIDTH - 1),
		23387 => to_unsigned(25655, LUT_AMPL_WIDTH - 1),
		23388 => to_unsigned(25653, LUT_AMPL_WIDTH - 1),
		23389 => to_unsigned(25651, LUT_AMPL_WIDTH - 1),
		23390 => to_unsigned(25649, LUT_AMPL_WIDTH - 1),
		23391 => to_unsigned(25647, LUT_AMPL_WIDTH - 1),
		23392 => to_unsigned(25645, LUT_AMPL_WIDTH - 1),
		23393 => to_unsigned(25643, LUT_AMPL_WIDTH - 1),
		23394 => to_unsigned(25641, LUT_AMPL_WIDTH - 1),
		23395 => to_unsigned(25639, LUT_AMPL_WIDTH - 1),
		23396 => to_unsigned(25637, LUT_AMPL_WIDTH - 1),
		23397 => to_unsigned(25635, LUT_AMPL_WIDTH - 1),
		23398 => to_unsigned(25633, LUT_AMPL_WIDTH - 1),
		23399 => to_unsigned(25631, LUT_AMPL_WIDTH - 1),
		23400 => to_unsigned(25629, LUT_AMPL_WIDTH - 1),
		23401 => to_unsigned(25628, LUT_AMPL_WIDTH - 1),
		23402 => to_unsigned(25626, LUT_AMPL_WIDTH - 1),
		23403 => to_unsigned(25624, LUT_AMPL_WIDTH - 1),
		23404 => to_unsigned(25622, LUT_AMPL_WIDTH - 1),
		23405 => to_unsigned(25620, LUT_AMPL_WIDTH - 1),
		23406 => to_unsigned(25618, LUT_AMPL_WIDTH - 1),
		23407 => to_unsigned(25616, LUT_AMPL_WIDTH - 1),
		23408 => to_unsigned(25614, LUT_AMPL_WIDTH - 1),
		23409 => to_unsigned(25612, LUT_AMPL_WIDTH - 1),
		23410 => to_unsigned(25610, LUT_AMPL_WIDTH - 1),
		23411 => to_unsigned(25608, LUT_AMPL_WIDTH - 1),
		23412 => to_unsigned(25606, LUT_AMPL_WIDTH - 1),
		23413 => to_unsigned(25604, LUT_AMPL_WIDTH - 1),
		23414 => to_unsigned(25602, LUT_AMPL_WIDTH - 1),
		23415 => to_unsigned(25600, LUT_AMPL_WIDTH - 1),
		23416 => to_unsigned(25598, LUT_AMPL_WIDTH - 1),
		23417 => to_unsigned(25596, LUT_AMPL_WIDTH - 1),
		23418 => to_unsigned(25594, LUT_AMPL_WIDTH - 1),
		23419 => to_unsigned(25592, LUT_AMPL_WIDTH - 1),
		23420 => to_unsigned(25590, LUT_AMPL_WIDTH - 1),
		23421 => to_unsigned(25588, LUT_AMPL_WIDTH - 1),
		23422 => to_unsigned(25586, LUT_AMPL_WIDTH - 1),
		23423 => to_unsigned(25584, LUT_AMPL_WIDTH - 1),
		23424 => to_unsigned(25582, LUT_AMPL_WIDTH - 1),
		23425 => to_unsigned(25580, LUT_AMPL_WIDTH - 1),
		23426 => to_unsigned(25578, LUT_AMPL_WIDTH - 1),
		23427 => to_unsigned(25577, LUT_AMPL_WIDTH - 1),
		23428 => to_unsigned(25575, LUT_AMPL_WIDTH - 1),
		23429 => to_unsigned(25573, LUT_AMPL_WIDTH - 1),
		23430 => to_unsigned(25571, LUT_AMPL_WIDTH - 1),
		23431 => to_unsigned(25569, LUT_AMPL_WIDTH - 1),
		23432 => to_unsigned(25567, LUT_AMPL_WIDTH - 1),
		23433 => to_unsigned(25565, LUT_AMPL_WIDTH - 1),
		23434 => to_unsigned(25563, LUT_AMPL_WIDTH - 1),
		23435 => to_unsigned(25561, LUT_AMPL_WIDTH - 1),
		23436 => to_unsigned(25559, LUT_AMPL_WIDTH - 1),
		23437 => to_unsigned(25557, LUT_AMPL_WIDTH - 1),
		23438 => to_unsigned(25555, LUT_AMPL_WIDTH - 1),
		23439 => to_unsigned(25553, LUT_AMPL_WIDTH - 1),
		23440 => to_unsigned(25551, LUT_AMPL_WIDTH - 1),
		23441 => to_unsigned(25549, LUT_AMPL_WIDTH - 1),
		23442 => to_unsigned(25547, LUT_AMPL_WIDTH - 1),
		23443 => to_unsigned(25545, LUT_AMPL_WIDTH - 1),
		23444 => to_unsigned(25543, LUT_AMPL_WIDTH - 1),
		23445 => to_unsigned(25541, LUT_AMPL_WIDTH - 1),
		23446 => to_unsigned(25539, LUT_AMPL_WIDTH - 1),
		23447 => to_unsigned(25537, LUT_AMPL_WIDTH - 1),
		23448 => to_unsigned(25535, LUT_AMPL_WIDTH - 1),
		23449 => to_unsigned(25533, LUT_AMPL_WIDTH - 1),
		23450 => to_unsigned(25531, LUT_AMPL_WIDTH - 1),
		23451 => to_unsigned(25529, LUT_AMPL_WIDTH - 1),
		23452 => to_unsigned(25527, LUT_AMPL_WIDTH - 1),
		23453 => to_unsigned(25525, LUT_AMPL_WIDTH - 1),
		23454 => to_unsigned(25523, LUT_AMPL_WIDTH - 1),
		23455 => to_unsigned(25521, LUT_AMPL_WIDTH - 1),
		23456 => to_unsigned(25519, LUT_AMPL_WIDTH - 1),
		23457 => to_unsigned(25518, LUT_AMPL_WIDTH - 1),
		23458 => to_unsigned(25516, LUT_AMPL_WIDTH - 1),
		23459 => to_unsigned(25514, LUT_AMPL_WIDTH - 1),
		23460 => to_unsigned(25512, LUT_AMPL_WIDTH - 1),
		23461 => to_unsigned(25510, LUT_AMPL_WIDTH - 1),
		23462 => to_unsigned(25508, LUT_AMPL_WIDTH - 1),
		23463 => to_unsigned(25506, LUT_AMPL_WIDTH - 1),
		23464 => to_unsigned(25504, LUT_AMPL_WIDTH - 1),
		23465 => to_unsigned(25502, LUT_AMPL_WIDTH - 1),
		23466 => to_unsigned(25500, LUT_AMPL_WIDTH - 1),
		23467 => to_unsigned(25498, LUT_AMPL_WIDTH - 1),
		23468 => to_unsigned(25496, LUT_AMPL_WIDTH - 1),
		23469 => to_unsigned(25494, LUT_AMPL_WIDTH - 1),
		23470 => to_unsigned(25492, LUT_AMPL_WIDTH - 1),
		23471 => to_unsigned(25490, LUT_AMPL_WIDTH - 1),
		23472 => to_unsigned(25488, LUT_AMPL_WIDTH - 1),
		23473 => to_unsigned(25486, LUT_AMPL_WIDTH - 1),
		23474 => to_unsigned(25484, LUT_AMPL_WIDTH - 1),
		23475 => to_unsigned(25482, LUT_AMPL_WIDTH - 1),
		23476 => to_unsigned(25480, LUT_AMPL_WIDTH - 1),
		23477 => to_unsigned(25478, LUT_AMPL_WIDTH - 1),
		23478 => to_unsigned(25476, LUT_AMPL_WIDTH - 1),
		23479 => to_unsigned(25474, LUT_AMPL_WIDTH - 1),
		23480 => to_unsigned(25472, LUT_AMPL_WIDTH - 1),
		23481 => to_unsigned(25470, LUT_AMPL_WIDTH - 1),
		23482 => to_unsigned(25468, LUT_AMPL_WIDTH - 1),
		23483 => to_unsigned(25466, LUT_AMPL_WIDTH - 1),
		23484 => to_unsigned(25464, LUT_AMPL_WIDTH - 1),
		23485 => to_unsigned(25462, LUT_AMPL_WIDTH - 1),
		23486 => to_unsigned(25460, LUT_AMPL_WIDTH - 1),
		23487 => to_unsigned(25458, LUT_AMPL_WIDTH - 1),
		23488 => to_unsigned(25456, LUT_AMPL_WIDTH - 1),
		23489 => to_unsigned(25454, LUT_AMPL_WIDTH - 1),
		23490 => to_unsigned(25452, LUT_AMPL_WIDTH - 1),
		23491 => to_unsigned(25450, LUT_AMPL_WIDTH - 1),
		23492 => to_unsigned(25448, LUT_AMPL_WIDTH - 1),
		23493 => to_unsigned(25446, LUT_AMPL_WIDTH - 1),
		23494 => to_unsigned(25444, LUT_AMPL_WIDTH - 1),
		23495 => to_unsigned(25442, LUT_AMPL_WIDTH - 1),
		23496 => to_unsigned(25440, LUT_AMPL_WIDTH - 1),
		23497 => to_unsigned(25438, LUT_AMPL_WIDTH - 1),
		23498 => to_unsigned(25437, LUT_AMPL_WIDTH - 1),
		23499 => to_unsigned(25435, LUT_AMPL_WIDTH - 1),
		23500 => to_unsigned(25433, LUT_AMPL_WIDTH - 1),
		23501 => to_unsigned(25431, LUT_AMPL_WIDTH - 1),
		23502 => to_unsigned(25429, LUT_AMPL_WIDTH - 1),
		23503 => to_unsigned(25427, LUT_AMPL_WIDTH - 1),
		23504 => to_unsigned(25425, LUT_AMPL_WIDTH - 1),
		23505 => to_unsigned(25423, LUT_AMPL_WIDTH - 1),
		23506 => to_unsigned(25421, LUT_AMPL_WIDTH - 1),
		23507 => to_unsigned(25419, LUT_AMPL_WIDTH - 1),
		23508 => to_unsigned(25417, LUT_AMPL_WIDTH - 1),
		23509 => to_unsigned(25415, LUT_AMPL_WIDTH - 1),
		23510 => to_unsigned(25413, LUT_AMPL_WIDTH - 1),
		23511 => to_unsigned(25411, LUT_AMPL_WIDTH - 1),
		23512 => to_unsigned(25409, LUT_AMPL_WIDTH - 1),
		23513 => to_unsigned(25407, LUT_AMPL_WIDTH - 1),
		23514 => to_unsigned(25405, LUT_AMPL_WIDTH - 1),
		23515 => to_unsigned(25403, LUT_AMPL_WIDTH - 1),
		23516 => to_unsigned(25401, LUT_AMPL_WIDTH - 1),
		23517 => to_unsigned(25399, LUT_AMPL_WIDTH - 1),
		23518 => to_unsigned(25397, LUT_AMPL_WIDTH - 1),
		23519 => to_unsigned(25395, LUT_AMPL_WIDTH - 1),
		23520 => to_unsigned(25393, LUT_AMPL_WIDTH - 1),
		23521 => to_unsigned(25391, LUT_AMPL_WIDTH - 1),
		23522 => to_unsigned(25389, LUT_AMPL_WIDTH - 1),
		23523 => to_unsigned(25387, LUT_AMPL_WIDTH - 1),
		23524 => to_unsigned(25385, LUT_AMPL_WIDTH - 1),
		23525 => to_unsigned(25383, LUT_AMPL_WIDTH - 1),
		23526 => to_unsigned(25381, LUT_AMPL_WIDTH - 1),
		23527 => to_unsigned(25379, LUT_AMPL_WIDTH - 1),
		23528 => to_unsigned(25377, LUT_AMPL_WIDTH - 1),
		23529 => to_unsigned(25375, LUT_AMPL_WIDTH - 1),
		23530 => to_unsigned(25373, LUT_AMPL_WIDTH - 1),
		23531 => to_unsigned(25371, LUT_AMPL_WIDTH - 1),
		23532 => to_unsigned(25369, LUT_AMPL_WIDTH - 1),
		23533 => to_unsigned(25367, LUT_AMPL_WIDTH - 1),
		23534 => to_unsigned(25365, LUT_AMPL_WIDTH - 1),
		23535 => to_unsigned(25363, LUT_AMPL_WIDTH - 1),
		23536 => to_unsigned(25361, LUT_AMPL_WIDTH - 1),
		23537 => to_unsigned(25359, LUT_AMPL_WIDTH - 1),
		23538 => to_unsigned(25357, LUT_AMPL_WIDTH - 1),
		23539 => to_unsigned(25355, LUT_AMPL_WIDTH - 1),
		23540 => to_unsigned(25353, LUT_AMPL_WIDTH - 1),
		23541 => to_unsigned(25351, LUT_AMPL_WIDTH - 1),
		23542 => to_unsigned(25349, LUT_AMPL_WIDTH - 1),
		23543 => to_unsigned(25347, LUT_AMPL_WIDTH - 1),
		23544 => to_unsigned(25345, LUT_AMPL_WIDTH - 1),
		23545 => to_unsigned(25343, LUT_AMPL_WIDTH - 1),
		23546 => to_unsigned(25341, LUT_AMPL_WIDTH - 1),
		23547 => to_unsigned(25339, LUT_AMPL_WIDTH - 1),
		23548 => to_unsigned(25337, LUT_AMPL_WIDTH - 1),
		23549 => to_unsigned(25335, LUT_AMPL_WIDTH - 1),
		23550 => to_unsigned(25333, LUT_AMPL_WIDTH - 1),
		23551 => to_unsigned(25331, LUT_AMPL_WIDTH - 1),
		23552 => to_unsigned(25329, LUT_AMPL_WIDTH - 1),
		23553 => to_unsigned(25327, LUT_AMPL_WIDTH - 1),
		23554 => to_unsigned(25325, LUT_AMPL_WIDTH - 1),
		23555 => to_unsigned(25323, LUT_AMPL_WIDTH - 1),
		23556 => to_unsigned(25321, LUT_AMPL_WIDTH - 1),
		23557 => to_unsigned(25319, LUT_AMPL_WIDTH - 1),
		23558 => to_unsigned(25317, LUT_AMPL_WIDTH - 1),
		23559 => to_unsigned(25315, LUT_AMPL_WIDTH - 1),
		23560 => to_unsigned(25313, LUT_AMPL_WIDTH - 1),
		23561 => to_unsigned(25311, LUT_AMPL_WIDTH - 1),
		23562 => to_unsigned(25309, LUT_AMPL_WIDTH - 1),
		23563 => to_unsigned(25307, LUT_AMPL_WIDTH - 1),
		23564 => to_unsigned(25305, LUT_AMPL_WIDTH - 1),
		23565 => to_unsigned(25303, LUT_AMPL_WIDTH - 1),
		23566 => to_unsigned(25301, LUT_AMPL_WIDTH - 1),
		23567 => to_unsigned(25299, LUT_AMPL_WIDTH - 1),
		23568 => to_unsigned(25297, LUT_AMPL_WIDTH - 1),
		23569 => to_unsigned(25295, LUT_AMPL_WIDTH - 1),
		23570 => to_unsigned(25293, LUT_AMPL_WIDTH - 1),
		23571 => to_unsigned(25291, LUT_AMPL_WIDTH - 1),
		23572 => to_unsigned(25289, LUT_AMPL_WIDTH - 1),
		23573 => to_unsigned(25287, LUT_AMPL_WIDTH - 1),
		23574 => to_unsigned(25285, LUT_AMPL_WIDTH - 1),
		23575 => to_unsigned(25283, LUT_AMPL_WIDTH - 1),
		23576 => to_unsigned(25281, LUT_AMPL_WIDTH - 1),
		23577 => to_unsigned(25279, LUT_AMPL_WIDTH - 1),
		23578 => to_unsigned(25277, LUT_AMPL_WIDTH - 1),
		23579 => to_unsigned(25275, LUT_AMPL_WIDTH - 1),
		23580 => to_unsigned(25273, LUT_AMPL_WIDTH - 1),
		23581 => to_unsigned(25271, LUT_AMPL_WIDTH - 1),
		23582 => to_unsigned(25269, LUT_AMPL_WIDTH - 1),
		23583 => to_unsigned(25267, LUT_AMPL_WIDTH - 1),
		23584 => to_unsigned(25265, LUT_AMPL_WIDTH - 1),
		23585 => to_unsigned(25263, LUT_AMPL_WIDTH - 1),
		23586 => to_unsigned(25261, LUT_AMPL_WIDTH - 1),
		23587 => to_unsigned(25259, LUT_AMPL_WIDTH - 1),
		23588 => to_unsigned(25257, LUT_AMPL_WIDTH - 1),
		23589 => to_unsigned(25255, LUT_AMPL_WIDTH - 1),
		23590 => to_unsigned(25253, LUT_AMPL_WIDTH - 1),
		23591 => to_unsigned(25251, LUT_AMPL_WIDTH - 1),
		23592 => to_unsigned(25249, LUT_AMPL_WIDTH - 1),
		23593 => to_unsigned(25247, LUT_AMPL_WIDTH - 1),
		23594 => to_unsigned(25245, LUT_AMPL_WIDTH - 1),
		23595 => to_unsigned(25243, LUT_AMPL_WIDTH - 1),
		23596 => to_unsigned(25241, LUT_AMPL_WIDTH - 1),
		23597 => to_unsigned(25239, LUT_AMPL_WIDTH - 1),
		23598 => to_unsigned(25237, LUT_AMPL_WIDTH - 1),
		23599 => to_unsigned(25235, LUT_AMPL_WIDTH - 1),
		23600 => to_unsigned(25233, LUT_AMPL_WIDTH - 1),
		23601 => to_unsigned(25231, LUT_AMPL_WIDTH - 1),
		23602 => to_unsigned(25229, LUT_AMPL_WIDTH - 1),
		23603 => to_unsigned(25227, LUT_AMPL_WIDTH - 1),
		23604 => to_unsigned(25225, LUT_AMPL_WIDTH - 1),
		23605 => to_unsigned(25223, LUT_AMPL_WIDTH - 1),
		23606 => to_unsigned(25221, LUT_AMPL_WIDTH - 1),
		23607 => to_unsigned(25219, LUT_AMPL_WIDTH - 1),
		23608 => to_unsigned(25217, LUT_AMPL_WIDTH - 1),
		23609 => to_unsigned(25215, LUT_AMPL_WIDTH - 1),
		23610 => to_unsigned(25213, LUT_AMPL_WIDTH - 1),
		23611 => to_unsigned(25211, LUT_AMPL_WIDTH - 1),
		23612 => to_unsigned(25209, LUT_AMPL_WIDTH - 1),
		23613 => to_unsigned(25207, LUT_AMPL_WIDTH - 1),
		23614 => to_unsigned(25205, LUT_AMPL_WIDTH - 1),
		23615 => to_unsigned(25203, LUT_AMPL_WIDTH - 1),
		23616 => to_unsigned(25201, LUT_AMPL_WIDTH - 1),
		23617 => to_unsigned(25199, LUT_AMPL_WIDTH - 1),
		23618 => to_unsigned(25197, LUT_AMPL_WIDTH - 1),
		23619 => to_unsigned(25195, LUT_AMPL_WIDTH - 1),
		23620 => to_unsigned(25193, LUT_AMPL_WIDTH - 1),
		23621 => to_unsigned(25191, LUT_AMPL_WIDTH - 1),
		23622 => to_unsigned(25189, LUT_AMPL_WIDTH - 1),
		23623 => to_unsigned(25187, LUT_AMPL_WIDTH - 1),
		23624 => to_unsigned(25185, LUT_AMPL_WIDTH - 1),
		23625 => to_unsigned(25183, LUT_AMPL_WIDTH - 1),
		23626 => to_unsigned(25181, LUT_AMPL_WIDTH - 1),
		23627 => to_unsigned(25179, LUT_AMPL_WIDTH - 1),
		23628 => to_unsigned(25177, LUT_AMPL_WIDTH - 1),
		23629 => to_unsigned(25175, LUT_AMPL_WIDTH - 1),
		23630 => to_unsigned(25173, LUT_AMPL_WIDTH - 1),
		23631 => to_unsigned(25171, LUT_AMPL_WIDTH - 1),
		23632 => to_unsigned(25169, LUT_AMPL_WIDTH - 1),
		23633 => to_unsigned(25167, LUT_AMPL_WIDTH - 1),
		23634 => to_unsigned(25165, LUT_AMPL_WIDTH - 1),
		23635 => to_unsigned(25163, LUT_AMPL_WIDTH - 1),
		23636 => to_unsigned(25161, LUT_AMPL_WIDTH - 1),
		23637 => to_unsigned(25159, LUT_AMPL_WIDTH - 1),
		23638 => to_unsigned(25157, LUT_AMPL_WIDTH - 1),
		23639 => to_unsigned(25155, LUT_AMPL_WIDTH - 1),
		23640 => to_unsigned(25153, LUT_AMPL_WIDTH - 1),
		23641 => to_unsigned(25151, LUT_AMPL_WIDTH - 1),
		23642 => to_unsigned(25149, LUT_AMPL_WIDTH - 1),
		23643 => to_unsigned(25147, LUT_AMPL_WIDTH - 1),
		23644 => to_unsigned(25145, LUT_AMPL_WIDTH - 1),
		23645 => to_unsigned(25143, LUT_AMPL_WIDTH - 1),
		23646 => to_unsigned(25141, LUT_AMPL_WIDTH - 1),
		23647 => to_unsigned(25139, LUT_AMPL_WIDTH - 1),
		23648 => to_unsigned(25137, LUT_AMPL_WIDTH - 1),
		23649 => to_unsigned(25135, LUT_AMPL_WIDTH - 1),
		23650 => to_unsigned(25133, LUT_AMPL_WIDTH - 1),
		23651 => to_unsigned(25131, LUT_AMPL_WIDTH - 1),
		23652 => to_unsigned(25129, LUT_AMPL_WIDTH - 1),
		23653 => to_unsigned(25127, LUT_AMPL_WIDTH - 1),
		23654 => to_unsigned(25125, LUT_AMPL_WIDTH - 1),
		23655 => to_unsigned(25123, LUT_AMPL_WIDTH - 1),
		23656 => to_unsigned(25121, LUT_AMPL_WIDTH - 1),
		23657 => to_unsigned(25119, LUT_AMPL_WIDTH - 1),
		23658 => to_unsigned(25117, LUT_AMPL_WIDTH - 1),
		23659 => to_unsigned(25115, LUT_AMPL_WIDTH - 1),
		23660 => to_unsigned(25113, LUT_AMPL_WIDTH - 1),
		23661 => to_unsigned(25111, LUT_AMPL_WIDTH - 1),
		23662 => to_unsigned(25109, LUT_AMPL_WIDTH - 1),
		23663 => to_unsigned(25107, LUT_AMPL_WIDTH - 1),
		23664 => to_unsigned(25105, LUT_AMPL_WIDTH - 1),
		23665 => to_unsigned(25103, LUT_AMPL_WIDTH - 1),
		23666 => to_unsigned(25101, LUT_AMPL_WIDTH - 1),
		23667 => to_unsigned(25099, LUT_AMPL_WIDTH - 1),
		23668 => to_unsigned(25096, LUT_AMPL_WIDTH - 1),
		23669 => to_unsigned(25094, LUT_AMPL_WIDTH - 1),
		23670 => to_unsigned(25092, LUT_AMPL_WIDTH - 1),
		23671 => to_unsigned(25090, LUT_AMPL_WIDTH - 1),
		23672 => to_unsigned(25088, LUT_AMPL_WIDTH - 1),
		23673 => to_unsigned(25086, LUT_AMPL_WIDTH - 1),
		23674 => to_unsigned(25084, LUT_AMPL_WIDTH - 1),
		23675 => to_unsigned(25082, LUT_AMPL_WIDTH - 1),
		23676 => to_unsigned(25080, LUT_AMPL_WIDTH - 1),
		23677 => to_unsigned(25078, LUT_AMPL_WIDTH - 1),
		23678 => to_unsigned(25076, LUT_AMPL_WIDTH - 1),
		23679 => to_unsigned(25074, LUT_AMPL_WIDTH - 1),
		23680 => to_unsigned(25072, LUT_AMPL_WIDTH - 1),
		23681 => to_unsigned(25070, LUT_AMPL_WIDTH - 1),
		23682 => to_unsigned(25068, LUT_AMPL_WIDTH - 1),
		23683 => to_unsigned(25066, LUT_AMPL_WIDTH - 1),
		23684 => to_unsigned(25064, LUT_AMPL_WIDTH - 1),
		23685 => to_unsigned(25062, LUT_AMPL_WIDTH - 1),
		23686 => to_unsigned(25060, LUT_AMPL_WIDTH - 1),
		23687 => to_unsigned(25058, LUT_AMPL_WIDTH - 1),
		23688 => to_unsigned(25056, LUT_AMPL_WIDTH - 1),
		23689 => to_unsigned(25054, LUT_AMPL_WIDTH - 1),
		23690 => to_unsigned(25052, LUT_AMPL_WIDTH - 1),
		23691 => to_unsigned(25050, LUT_AMPL_WIDTH - 1),
		23692 => to_unsigned(25048, LUT_AMPL_WIDTH - 1),
		23693 => to_unsigned(25046, LUT_AMPL_WIDTH - 1),
		23694 => to_unsigned(25044, LUT_AMPL_WIDTH - 1),
		23695 => to_unsigned(25042, LUT_AMPL_WIDTH - 1),
		23696 => to_unsigned(25040, LUT_AMPL_WIDTH - 1),
		23697 => to_unsigned(25038, LUT_AMPL_WIDTH - 1),
		23698 => to_unsigned(25036, LUT_AMPL_WIDTH - 1),
		23699 => to_unsigned(25034, LUT_AMPL_WIDTH - 1),
		23700 => to_unsigned(25032, LUT_AMPL_WIDTH - 1),
		23701 => to_unsigned(25030, LUT_AMPL_WIDTH - 1),
		23702 => to_unsigned(25028, LUT_AMPL_WIDTH - 1),
		23703 => to_unsigned(25026, LUT_AMPL_WIDTH - 1),
		23704 => to_unsigned(25024, LUT_AMPL_WIDTH - 1),
		23705 => to_unsigned(25022, LUT_AMPL_WIDTH - 1),
		23706 => to_unsigned(25020, LUT_AMPL_WIDTH - 1),
		23707 => to_unsigned(25018, LUT_AMPL_WIDTH - 1),
		23708 => to_unsigned(25016, LUT_AMPL_WIDTH - 1),
		23709 => to_unsigned(25013, LUT_AMPL_WIDTH - 1),
		23710 => to_unsigned(25011, LUT_AMPL_WIDTH - 1),
		23711 => to_unsigned(25009, LUT_AMPL_WIDTH - 1),
		23712 => to_unsigned(25007, LUT_AMPL_WIDTH - 1),
		23713 => to_unsigned(25005, LUT_AMPL_WIDTH - 1),
		23714 => to_unsigned(25003, LUT_AMPL_WIDTH - 1),
		23715 => to_unsigned(25001, LUT_AMPL_WIDTH - 1),
		23716 => to_unsigned(24999, LUT_AMPL_WIDTH - 1),
		23717 => to_unsigned(24997, LUT_AMPL_WIDTH - 1),
		23718 => to_unsigned(24995, LUT_AMPL_WIDTH - 1),
		23719 => to_unsigned(24993, LUT_AMPL_WIDTH - 1),
		23720 => to_unsigned(24991, LUT_AMPL_WIDTH - 1),
		23721 => to_unsigned(24989, LUT_AMPL_WIDTH - 1),
		23722 => to_unsigned(24987, LUT_AMPL_WIDTH - 1),
		23723 => to_unsigned(24985, LUT_AMPL_WIDTH - 1),
		23724 => to_unsigned(24983, LUT_AMPL_WIDTH - 1),
		23725 => to_unsigned(24981, LUT_AMPL_WIDTH - 1),
		23726 => to_unsigned(24979, LUT_AMPL_WIDTH - 1),
		23727 => to_unsigned(24977, LUT_AMPL_WIDTH - 1),
		23728 => to_unsigned(24975, LUT_AMPL_WIDTH - 1),
		23729 => to_unsigned(24973, LUT_AMPL_WIDTH - 1),
		23730 => to_unsigned(24971, LUT_AMPL_WIDTH - 1),
		23731 => to_unsigned(24969, LUT_AMPL_WIDTH - 1),
		23732 => to_unsigned(24967, LUT_AMPL_WIDTH - 1),
		23733 => to_unsigned(24965, LUT_AMPL_WIDTH - 1),
		23734 => to_unsigned(24963, LUT_AMPL_WIDTH - 1),
		23735 => to_unsigned(24961, LUT_AMPL_WIDTH - 1),
		23736 => to_unsigned(24959, LUT_AMPL_WIDTH - 1),
		23737 => to_unsigned(24957, LUT_AMPL_WIDTH - 1),
		23738 => to_unsigned(24955, LUT_AMPL_WIDTH - 1),
		23739 => to_unsigned(24953, LUT_AMPL_WIDTH - 1),
		23740 => to_unsigned(24950, LUT_AMPL_WIDTH - 1),
		23741 => to_unsigned(24948, LUT_AMPL_WIDTH - 1),
		23742 => to_unsigned(24946, LUT_AMPL_WIDTH - 1),
		23743 => to_unsigned(24944, LUT_AMPL_WIDTH - 1),
		23744 => to_unsigned(24942, LUT_AMPL_WIDTH - 1),
		23745 => to_unsigned(24940, LUT_AMPL_WIDTH - 1),
		23746 => to_unsigned(24938, LUT_AMPL_WIDTH - 1),
		23747 => to_unsigned(24936, LUT_AMPL_WIDTH - 1),
		23748 => to_unsigned(24934, LUT_AMPL_WIDTH - 1),
		23749 => to_unsigned(24932, LUT_AMPL_WIDTH - 1),
		23750 => to_unsigned(24930, LUT_AMPL_WIDTH - 1),
		23751 => to_unsigned(24928, LUT_AMPL_WIDTH - 1),
		23752 => to_unsigned(24926, LUT_AMPL_WIDTH - 1),
		23753 => to_unsigned(24924, LUT_AMPL_WIDTH - 1),
		23754 => to_unsigned(24922, LUT_AMPL_WIDTH - 1),
		23755 => to_unsigned(24920, LUT_AMPL_WIDTH - 1),
		23756 => to_unsigned(24918, LUT_AMPL_WIDTH - 1),
		23757 => to_unsigned(24916, LUT_AMPL_WIDTH - 1),
		23758 => to_unsigned(24914, LUT_AMPL_WIDTH - 1),
		23759 => to_unsigned(24912, LUT_AMPL_WIDTH - 1),
		23760 => to_unsigned(24910, LUT_AMPL_WIDTH - 1),
		23761 => to_unsigned(24908, LUT_AMPL_WIDTH - 1),
		23762 => to_unsigned(24906, LUT_AMPL_WIDTH - 1),
		23763 => to_unsigned(24904, LUT_AMPL_WIDTH - 1),
		23764 => to_unsigned(24902, LUT_AMPL_WIDTH - 1),
		23765 => to_unsigned(24899, LUT_AMPL_WIDTH - 1),
		23766 => to_unsigned(24897, LUT_AMPL_WIDTH - 1),
		23767 => to_unsigned(24895, LUT_AMPL_WIDTH - 1),
		23768 => to_unsigned(24893, LUT_AMPL_WIDTH - 1),
		23769 => to_unsigned(24891, LUT_AMPL_WIDTH - 1),
		23770 => to_unsigned(24889, LUT_AMPL_WIDTH - 1),
		23771 => to_unsigned(24887, LUT_AMPL_WIDTH - 1),
		23772 => to_unsigned(24885, LUT_AMPL_WIDTH - 1),
		23773 => to_unsigned(24883, LUT_AMPL_WIDTH - 1),
		23774 => to_unsigned(24881, LUT_AMPL_WIDTH - 1),
		23775 => to_unsigned(24879, LUT_AMPL_WIDTH - 1),
		23776 => to_unsigned(24877, LUT_AMPL_WIDTH - 1),
		23777 => to_unsigned(24875, LUT_AMPL_WIDTH - 1),
		23778 => to_unsigned(24873, LUT_AMPL_WIDTH - 1),
		23779 => to_unsigned(24871, LUT_AMPL_WIDTH - 1),
		23780 => to_unsigned(24869, LUT_AMPL_WIDTH - 1),
		23781 => to_unsigned(24867, LUT_AMPL_WIDTH - 1),
		23782 => to_unsigned(24865, LUT_AMPL_WIDTH - 1),
		23783 => to_unsigned(24863, LUT_AMPL_WIDTH - 1),
		23784 => to_unsigned(24861, LUT_AMPL_WIDTH - 1),
		23785 => to_unsigned(24859, LUT_AMPL_WIDTH - 1),
		23786 => to_unsigned(24857, LUT_AMPL_WIDTH - 1),
		23787 => to_unsigned(24855, LUT_AMPL_WIDTH - 1),
		23788 => to_unsigned(24852, LUT_AMPL_WIDTH - 1),
		23789 => to_unsigned(24850, LUT_AMPL_WIDTH - 1),
		23790 => to_unsigned(24848, LUT_AMPL_WIDTH - 1),
		23791 => to_unsigned(24846, LUT_AMPL_WIDTH - 1),
		23792 => to_unsigned(24844, LUT_AMPL_WIDTH - 1),
		23793 => to_unsigned(24842, LUT_AMPL_WIDTH - 1),
		23794 => to_unsigned(24840, LUT_AMPL_WIDTH - 1),
		23795 => to_unsigned(24838, LUT_AMPL_WIDTH - 1),
		23796 => to_unsigned(24836, LUT_AMPL_WIDTH - 1),
		23797 => to_unsigned(24834, LUT_AMPL_WIDTH - 1),
		23798 => to_unsigned(24832, LUT_AMPL_WIDTH - 1),
		23799 => to_unsigned(24830, LUT_AMPL_WIDTH - 1),
		23800 => to_unsigned(24828, LUT_AMPL_WIDTH - 1),
		23801 => to_unsigned(24826, LUT_AMPL_WIDTH - 1),
		23802 => to_unsigned(24824, LUT_AMPL_WIDTH - 1),
		23803 => to_unsigned(24822, LUT_AMPL_WIDTH - 1),
		23804 => to_unsigned(24820, LUT_AMPL_WIDTH - 1),
		23805 => to_unsigned(24818, LUT_AMPL_WIDTH - 1),
		23806 => to_unsigned(24816, LUT_AMPL_WIDTH - 1),
		23807 => to_unsigned(24814, LUT_AMPL_WIDTH - 1),
		23808 => to_unsigned(24811, LUT_AMPL_WIDTH - 1),
		23809 => to_unsigned(24809, LUT_AMPL_WIDTH - 1),
		23810 => to_unsigned(24807, LUT_AMPL_WIDTH - 1),
		23811 => to_unsigned(24805, LUT_AMPL_WIDTH - 1),
		23812 => to_unsigned(24803, LUT_AMPL_WIDTH - 1),
		23813 => to_unsigned(24801, LUT_AMPL_WIDTH - 1),
		23814 => to_unsigned(24799, LUT_AMPL_WIDTH - 1),
		23815 => to_unsigned(24797, LUT_AMPL_WIDTH - 1),
		23816 => to_unsigned(24795, LUT_AMPL_WIDTH - 1),
		23817 => to_unsigned(24793, LUT_AMPL_WIDTH - 1),
		23818 => to_unsigned(24791, LUT_AMPL_WIDTH - 1),
		23819 => to_unsigned(24789, LUT_AMPL_WIDTH - 1),
		23820 => to_unsigned(24787, LUT_AMPL_WIDTH - 1),
		23821 => to_unsigned(24785, LUT_AMPL_WIDTH - 1),
		23822 => to_unsigned(24783, LUT_AMPL_WIDTH - 1),
		23823 => to_unsigned(24781, LUT_AMPL_WIDTH - 1),
		23824 => to_unsigned(24779, LUT_AMPL_WIDTH - 1),
		23825 => to_unsigned(24777, LUT_AMPL_WIDTH - 1),
		23826 => to_unsigned(24774, LUT_AMPL_WIDTH - 1),
		23827 => to_unsigned(24772, LUT_AMPL_WIDTH - 1),
		23828 => to_unsigned(24770, LUT_AMPL_WIDTH - 1),
		23829 => to_unsigned(24768, LUT_AMPL_WIDTH - 1),
		23830 => to_unsigned(24766, LUT_AMPL_WIDTH - 1),
		23831 => to_unsigned(24764, LUT_AMPL_WIDTH - 1),
		23832 => to_unsigned(24762, LUT_AMPL_WIDTH - 1),
		23833 => to_unsigned(24760, LUT_AMPL_WIDTH - 1),
		23834 => to_unsigned(24758, LUT_AMPL_WIDTH - 1),
		23835 => to_unsigned(24756, LUT_AMPL_WIDTH - 1),
		23836 => to_unsigned(24754, LUT_AMPL_WIDTH - 1),
		23837 => to_unsigned(24752, LUT_AMPL_WIDTH - 1),
		23838 => to_unsigned(24750, LUT_AMPL_WIDTH - 1),
		23839 => to_unsigned(24748, LUT_AMPL_WIDTH - 1),
		23840 => to_unsigned(24746, LUT_AMPL_WIDTH - 1),
		23841 => to_unsigned(24744, LUT_AMPL_WIDTH - 1),
		23842 => to_unsigned(24742, LUT_AMPL_WIDTH - 1),
		23843 => to_unsigned(24740, LUT_AMPL_WIDTH - 1),
		23844 => to_unsigned(24737, LUT_AMPL_WIDTH - 1),
		23845 => to_unsigned(24735, LUT_AMPL_WIDTH - 1),
		23846 => to_unsigned(24733, LUT_AMPL_WIDTH - 1),
		23847 => to_unsigned(24731, LUT_AMPL_WIDTH - 1),
		23848 => to_unsigned(24729, LUT_AMPL_WIDTH - 1),
		23849 => to_unsigned(24727, LUT_AMPL_WIDTH - 1),
		23850 => to_unsigned(24725, LUT_AMPL_WIDTH - 1),
		23851 => to_unsigned(24723, LUT_AMPL_WIDTH - 1),
		23852 => to_unsigned(24721, LUT_AMPL_WIDTH - 1),
		23853 => to_unsigned(24719, LUT_AMPL_WIDTH - 1),
		23854 => to_unsigned(24717, LUT_AMPL_WIDTH - 1),
		23855 => to_unsigned(24715, LUT_AMPL_WIDTH - 1),
		23856 => to_unsigned(24713, LUT_AMPL_WIDTH - 1),
		23857 => to_unsigned(24711, LUT_AMPL_WIDTH - 1),
		23858 => to_unsigned(24709, LUT_AMPL_WIDTH - 1),
		23859 => to_unsigned(24707, LUT_AMPL_WIDTH - 1),
		23860 => to_unsigned(24704, LUT_AMPL_WIDTH - 1),
		23861 => to_unsigned(24702, LUT_AMPL_WIDTH - 1),
		23862 => to_unsigned(24700, LUT_AMPL_WIDTH - 1),
		23863 => to_unsigned(24698, LUT_AMPL_WIDTH - 1),
		23864 => to_unsigned(24696, LUT_AMPL_WIDTH - 1),
		23865 => to_unsigned(24694, LUT_AMPL_WIDTH - 1),
		23866 => to_unsigned(24692, LUT_AMPL_WIDTH - 1),
		23867 => to_unsigned(24690, LUT_AMPL_WIDTH - 1),
		23868 => to_unsigned(24688, LUT_AMPL_WIDTH - 1),
		23869 => to_unsigned(24686, LUT_AMPL_WIDTH - 1),
		23870 => to_unsigned(24684, LUT_AMPL_WIDTH - 1),
		23871 => to_unsigned(24682, LUT_AMPL_WIDTH - 1),
		23872 => to_unsigned(24680, LUT_AMPL_WIDTH - 1),
		23873 => to_unsigned(24678, LUT_AMPL_WIDTH - 1),
		23874 => to_unsigned(24676, LUT_AMPL_WIDTH - 1),
		23875 => to_unsigned(24673, LUT_AMPL_WIDTH - 1),
		23876 => to_unsigned(24671, LUT_AMPL_WIDTH - 1),
		23877 => to_unsigned(24669, LUT_AMPL_WIDTH - 1),
		23878 => to_unsigned(24667, LUT_AMPL_WIDTH - 1),
		23879 => to_unsigned(24665, LUT_AMPL_WIDTH - 1),
		23880 => to_unsigned(24663, LUT_AMPL_WIDTH - 1),
		23881 => to_unsigned(24661, LUT_AMPL_WIDTH - 1),
		23882 => to_unsigned(24659, LUT_AMPL_WIDTH - 1),
		23883 => to_unsigned(24657, LUT_AMPL_WIDTH - 1),
		23884 => to_unsigned(24655, LUT_AMPL_WIDTH - 1),
		23885 => to_unsigned(24653, LUT_AMPL_WIDTH - 1),
		23886 => to_unsigned(24651, LUT_AMPL_WIDTH - 1),
		23887 => to_unsigned(24649, LUT_AMPL_WIDTH - 1),
		23888 => to_unsigned(24647, LUT_AMPL_WIDTH - 1),
		23889 => to_unsigned(24645, LUT_AMPL_WIDTH - 1),
		23890 => to_unsigned(24642, LUT_AMPL_WIDTH - 1),
		23891 => to_unsigned(24640, LUT_AMPL_WIDTH - 1),
		23892 => to_unsigned(24638, LUT_AMPL_WIDTH - 1),
		23893 => to_unsigned(24636, LUT_AMPL_WIDTH - 1),
		23894 => to_unsigned(24634, LUT_AMPL_WIDTH - 1),
		23895 => to_unsigned(24632, LUT_AMPL_WIDTH - 1),
		23896 => to_unsigned(24630, LUT_AMPL_WIDTH - 1),
		23897 => to_unsigned(24628, LUT_AMPL_WIDTH - 1),
		23898 => to_unsigned(24626, LUT_AMPL_WIDTH - 1),
		23899 => to_unsigned(24624, LUT_AMPL_WIDTH - 1),
		23900 => to_unsigned(24622, LUT_AMPL_WIDTH - 1),
		23901 => to_unsigned(24620, LUT_AMPL_WIDTH - 1),
		23902 => to_unsigned(24618, LUT_AMPL_WIDTH - 1),
		23903 => to_unsigned(24616, LUT_AMPL_WIDTH - 1),
		23904 => to_unsigned(24613, LUT_AMPL_WIDTH - 1),
		23905 => to_unsigned(24611, LUT_AMPL_WIDTH - 1),
		23906 => to_unsigned(24609, LUT_AMPL_WIDTH - 1),
		23907 => to_unsigned(24607, LUT_AMPL_WIDTH - 1),
		23908 => to_unsigned(24605, LUT_AMPL_WIDTH - 1),
		23909 => to_unsigned(24603, LUT_AMPL_WIDTH - 1),
		23910 => to_unsigned(24601, LUT_AMPL_WIDTH - 1),
		23911 => to_unsigned(24599, LUT_AMPL_WIDTH - 1),
		23912 => to_unsigned(24597, LUT_AMPL_WIDTH - 1),
		23913 => to_unsigned(24595, LUT_AMPL_WIDTH - 1),
		23914 => to_unsigned(24593, LUT_AMPL_WIDTH - 1),
		23915 => to_unsigned(24591, LUT_AMPL_WIDTH - 1),
		23916 => to_unsigned(24589, LUT_AMPL_WIDTH - 1),
		23917 => to_unsigned(24586, LUT_AMPL_WIDTH - 1),
		23918 => to_unsigned(24584, LUT_AMPL_WIDTH - 1),
		23919 => to_unsigned(24582, LUT_AMPL_WIDTH - 1),
		23920 => to_unsigned(24580, LUT_AMPL_WIDTH - 1),
		23921 => to_unsigned(24578, LUT_AMPL_WIDTH - 1),
		23922 => to_unsigned(24576, LUT_AMPL_WIDTH - 1),
		23923 => to_unsigned(24574, LUT_AMPL_WIDTH - 1),
		23924 => to_unsigned(24572, LUT_AMPL_WIDTH - 1),
		23925 => to_unsigned(24570, LUT_AMPL_WIDTH - 1),
		23926 => to_unsigned(24568, LUT_AMPL_WIDTH - 1),
		23927 => to_unsigned(24566, LUT_AMPL_WIDTH - 1),
		23928 => to_unsigned(24564, LUT_AMPL_WIDTH - 1),
		23929 => to_unsigned(24562, LUT_AMPL_WIDTH - 1),
		23930 => to_unsigned(24559, LUT_AMPL_WIDTH - 1),
		23931 => to_unsigned(24557, LUT_AMPL_WIDTH - 1),
		23932 => to_unsigned(24555, LUT_AMPL_WIDTH - 1),
		23933 => to_unsigned(24553, LUT_AMPL_WIDTH - 1),
		23934 => to_unsigned(24551, LUT_AMPL_WIDTH - 1),
		23935 => to_unsigned(24549, LUT_AMPL_WIDTH - 1),
		23936 => to_unsigned(24547, LUT_AMPL_WIDTH - 1),
		23937 => to_unsigned(24545, LUT_AMPL_WIDTH - 1),
		23938 => to_unsigned(24543, LUT_AMPL_WIDTH - 1),
		23939 => to_unsigned(24541, LUT_AMPL_WIDTH - 1),
		23940 => to_unsigned(24539, LUT_AMPL_WIDTH - 1),
		23941 => to_unsigned(24537, LUT_AMPL_WIDTH - 1),
		23942 => to_unsigned(24534, LUT_AMPL_WIDTH - 1),
		23943 => to_unsigned(24532, LUT_AMPL_WIDTH - 1),
		23944 => to_unsigned(24530, LUT_AMPL_WIDTH - 1),
		23945 => to_unsigned(24528, LUT_AMPL_WIDTH - 1),
		23946 => to_unsigned(24526, LUT_AMPL_WIDTH - 1),
		23947 => to_unsigned(24524, LUT_AMPL_WIDTH - 1),
		23948 => to_unsigned(24522, LUT_AMPL_WIDTH - 1),
		23949 => to_unsigned(24520, LUT_AMPL_WIDTH - 1),
		23950 => to_unsigned(24518, LUT_AMPL_WIDTH - 1),
		23951 => to_unsigned(24516, LUT_AMPL_WIDTH - 1),
		23952 => to_unsigned(24514, LUT_AMPL_WIDTH - 1),
		23953 => to_unsigned(24512, LUT_AMPL_WIDTH - 1),
		23954 => to_unsigned(24509, LUT_AMPL_WIDTH - 1),
		23955 => to_unsigned(24507, LUT_AMPL_WIDTH - 1),
		23956 => to_unsigned(24505, LUT_AMPL_WIDTH - 1),
		23957 => to_unsigned(24503, LUT_AMPL_WIDTH - 1),
		23958 => to_unsigned(24501, LUT_AMPL_WIDTH - 1),
		23959 => to_unsigned(24499, LUT_AMPL_WIDTH - 1),
		23960 => to_unsigned(24497, LUT_AMPL_WIDTH - 1),
		23961 => to_unsigned(24495, LUT_AMPL_WIDTH - 1),
		23962 => to_unsigned(24493, LUT_AMPL_WIDTH - 1),
		23963 => to_unsigned(24491, LUT_AMPL_WIDTH - 1),
		23964 => to_unsigned(24489, LUT_AMPL_WIDTH - 1),
		23965 => to_unsigned(24487, LUT_AMPL_WIDTH - 1),
		23966 => to_unsigned(24484, LUT_AMPL_WIDTH - 1),
		23967 => to_unsigned(24482, LUT_AMPL_WIDTH - 1),
		23968 => to_unsigned(24480, LUT_AMPL_WIDTH - 1),
		23969 => to_unsigned(24478, LUT_AMPL_WIDTH - 1),
		23970 => to_unsigned(24476, LUT_AMPL_WIDTH - 1),
		23971 => to_unsigned(24474, LUT_AMPL_WIDTH - 1),
		23972 => to_unsigned(24472, LUT_AMPL_WIDTH - 1),
		23973 => to_unsigned(24470, LUT_AMPL_WIDTH - 1),
		23974 => to_unsigned(24468, LUT_AMPL_WIDTH - 1),
		23975 => to_unsigned(24466, LUT_AMPL_WIDTH - 1),
		23976 => to_unsigned(24464, LUT_AMPL_WIDTH - 1),
		23977 => to_unsigned(24461, LUT_AMPL_WIDTH - 1),
		23978 => to_unsigned(24459, LUT_AMPL_WIDTH - 1),
		23979 => to_unsigned(24457, LUT_AMPL_WIDTH - 1),
		23980 => to_unsigned(24455, LUT_AMPL_WIDTH - 1),
		23981 => to_unsigned(24453, LUT_AMPL_WIDTH - 1),
		23982 => to_unsigned(24451, LUT_AMPL_WIDTH - 1),
		23983 => to_unsigned(24449, LUT_AMPL_WIDTH - 1),
		23984 => to_unsigned(24447, LUT_AMPL_WIDTH - 1),
		23985 => to_unsigned(24445, LUT_AMPL_WIDTH - 1),
		23986 => to_unsigned(24443, LUT_AMPL_WIDTH - 1),
		23987 => to_unsigned(24441, LUT_AMPL_WIDTH - 1),
		23988 => to_unsigned(24438, LUT_AMPL_WIDTH - 1),
		23989 => to_unsigned(24436, LUT_AMPL_WIDTH - 1),
		23990 => to_unsigned(24434, LUT_AMPL_WIDTH - 1),
		23991 => to_unsigned(24432, LUT_AMPL_WIDTH - 1),
		23992 => to_unsigned(24430, LUT_AMPL_WIDTH - 1),
		23993 => to_unsigned(24428, LUT_AMPL_WIDTH - 1),
		23994 => to_unsigned(24426, LUT_AMPL_WIDTH - 1),
		23995 => to_unsigned(24424, LUT_AMPL_WIDTH - 1),
		23996 => to_unsigned(24422, LUT_AMPL_WIDTH - 1),
		23997 => to_unsigned(24420, LUT_AMPL_WIDTH - 1),
		23998 => to_unsigned(24417, LUT_AMPL_WIDTH - 1),
		23999 => to_unsigned(24415, LUT_AMPL_WIDTH - 1),
		24000 => to_unsigned(24413, LUT_AMPL_WIDTH - 1),
		24001 => to_unsigned(24411, LUT_AMPL_WIDTH - 1),
		24002 => to_unsigned(24409, LUT_AMPL_WIDTH - 1),
		24003 => to_unsigned(24407, LUT_AMPL_WIDTH - 1),
		24004 => to_unsigned(24405, LUT_AMPL_WIDTH - 1),
		24005 => to_unsigned(24403, LUT_AMPL_WIDTH - 1),
		24006 => to_unsigned(24401, LUT_AMPL_WIDTH - 1),
		24007 => to_unsigned(24399, LUT_AMPL_WIDTH - 1),
		24008 => to_unsigned(24397, LUT_AMPL_WIDTH - 1),
		24009 => to_unsigned(24394, LUT_AMPL_WIDTH - 1),
		24010 => to_unsigned(24392, LUT_AMPL_WIDTH - 1),
		24011 => to_unsigned(24390, LUT_AMPL_WIDTH - 1),
		24012 => to_unsigned(24388, LUT_AMPL_WIDTH - 1),
		24013 => to_unsigned(24386, LUT_AMPL_WIDTH - 1),
		24014 => to_unsigned(24384, LUT_AMPL_WIDTH - 1),
		24015 => to_unsigned(24382, LUT_AMPL_WIDTH - 1),
		24016 => to_unsigned(24380, LUT_AMPL_WIDTH - 1),
		24017 => to_unsigned(24378, LUT_AMPL_WIDTH - 1),
		24018 => to_unsigned(24376, LUT_AMPL_WIDTH - 1),
		24019 => to_unsigned(24373, LUT_AMPL_WIDTH - 1),
		24020 => to_unsigned(24371, LUT_AMPL_WIDTH - 1),
		24021 => to_unsigned(24369, LUT_AMPL_WIDTH - 1),
		24022 => to_unsigned(24367, LUT_AMPL_WIDTH - 1),
		24023 => to_unsigned(24365, LUT_AMPL_WIDTH - 1),
		24024 => to_unsigned(24363, LUT_AMPL_WIDTH - 1),
		24025 => to_unsigned(24361, LUT_AMPL_WIDTH - 1),
		24026 => to_unsigned(24359, LUT_AMPL_WIDTH - 1),
		24027 => to_unsigned(24357, LUT_AMPL_WIDTH - 1),
		24028 => to_unsigned(24355, LUT_AMPL_WIDTH - 1),
		24029 => to_unsigned(24352, LUT_AMPL_WIDTH - 1),
		24030 => to_unsigned(24350, LUT_AMPL_WIDTH - 1),
		24031 => to_unsigned(24348, LUT_AMPL_WIDTH - 1),
		24032 => to_unsigned(24346, LUT_AMPL_WIDTH - 1),
		24033 => to_unsigned(24344, LUT_AMPL_WIDTH - 1),
		24034 => to_unsigned(24342, LUT_AMPL_WIDTH - 1),
		24035 => to_unsigned(24340, LUT_AMPL_WIDTH - 1),
		24036 => to_unsigned(24338, LUT_AMPL_WIDTH - 1),
		24037 => to_unsigned(24336, LUT_AMPL_WIDTH - 1),
		24038 => to_unsigned(24334, LUT_AMPL_WIDTH - 1),
		24039 => to_unsigned(24331, LUT_AMPL_WIDTH - 1),
		24040 => to_unsigned(24329, LUT_AMPL_WIDTH - 1),
		24041 => to_unsigned(24327, LUT_AMPL_WIDTH - 1),
		24042 => to_unsigned(24325, LUT_AMPL_WIDTH - 1),
		24043 => to_unsigned(24323, LUT_AMPL_WIDTH - 1),
		24044 => to_unsigned(24321, LUT_AMPL_WIDTH - 1),
		24045 => to_unsigned(24319, LUT_AMPL_WIDTH - 1),
		24046 => to_unsigned(24317, LUT_AMPL_WIDTH - 1),
		24047 => to_unsigned(24315, LUT_AMPL_WIDTH - 1),
		24048 => to_unsigned(24312, LUT_AMPL_WIDTH - 1),
		24049 => to_unsigned(24310, LUT_AMPL_WIDTH - 1),
		24050 => to_unsigned(24308, LUT_AMPL_WIDTH - 1),
		24051 => to_unsigned(24306, LUT_AMPL_WIDTH - 1),
		24052 => to_unsigned(24304, LUT_AMPL_WIDTH - 1),
		24053 => to_unsigned(24302, LUT_AMPL_WIDTH - 1),
		24054 => to_unsigned(24300, LUT_AMPL_WIDTH - 1),
		24055 => to_unsigned(24298, LUT_AMPL_WIDTH - 1),
		24056 => to_unsigned(24296, LUT_AMPL_WIDTH - 1),
		24057 => to_unsigned(24294, LUT_AMPL_WIDTH - 1),
		24058 => to_unsigned(24291, LUT_AMPL_WIDTH - 1),
		24059 => to_unsigned(24289, LUT_AMPL_WIDTH - 1),
		24060 => to_unsigned(24287, LUT_AMPL_WIDTH - 1),
		24061 => to_unsigned(24285, LUT_AMPL_WIDTH - 1),
		24062 => to_unsigned(24283, LUT_AMPL_WIDTH - 1),
		24063 => to_unsigned(24281, LUT_AMPL_WIDTH - 1),
		24064 => to_unsigned(24279, LUT_AMPL_WIDTH - 1),
		24065 => to_unsigned(24277, LUT_AMPL_WIDTH - 1),
		24066 => to_unsigned(24275, LUT_AMPL_WIDTH - 1),
		24067 => to_unsigned(24272, LUT_AMPL_WIDTH - 1),
		24068 => to_unsigned(24270, LUT_AMPL_WIDTH - 1),
		24069 => to_unsigned(24268, LUT_AMPL_WIDTH - 1),
		24070 => to_unsigned(24266, LUT_AMPL_WIDTH - 1),
		24071 => to_unsigned(24264, LUT_AMPL_WIDTH - 1),
		24072 => to_unsigned(24262, LUT_AMPL_WIDTH - 1),
		24073 => to_unsigned(24260, LUT_AMPL_WIDTH - 1),
		24074 => to_unsigned(24258, LUT_AMPL_WIDTH - 1),
		24075 => to_unsigned(24256, LUT_AMPL_WIDTH - 1),
		24076 => to_unsigned(24253, LUT_AMPL_WIDTH - 1),
		24077 => to_unsigned(24251, LUT_AMPL_WIDTH - 1),
		24078 => to_unsigned(24249, LUT_AMPL_WIDTH - 1),
		24079 => to_unsigned(24247, LUT_AMPL_WIDTH - 1),
		24080 => to_unsigned(24245, LUT_AMPL_WIDTH - 1),
		24081 => to_unsigned(24243, LUT_AMPL_WIDTH - 1),
		24082 => to_unsigned(24241, LUT_AMPL_WIDTH - 1),
		24083 => to_unsigned(24239, LUT_AMPL_WIDTH - 1),
		24084 => to_unsigned(24237, LUT_AMPL_WIDTH - 1),
		24085 => to_unsigned(24234, LUT_AMPL_WIDTH - 1),
		24086 => to_unsigned(24232, LUT_AMPL_WIDTH - 1),
		24087 => to_unsigned(24230, LUT_AMPL_WIDTH - 1),
		24088 => to_unsigned(24228, LUT_AMPL_WIDTH - 1),
		24089 => to_unsigned(24226, LUT_AMPL_WIDTH - 1),
		24090 => to_unsigned(24224, LUT_AMPL_WIDTH - 1),
		24091 => to_unsigned(24222, LUT_AMPL_WIDTH - 1),
		24092 => to_unsigned(24220, LUT_AMPL_WIDTH - 1),
		24093 => to_unsigned(24217, LUT_AMPL_WIDTH - 1),
		24094 => to_unsigned(24215, LUT_AMPL_WIDTH - 1),
		24095 => to_unsigned(24213, LUT_AMPL_WIDTH - 1),
		24096 => to_unsigned(24211, LUT_AMPL_WIDTH - 1),
		24097 => to_unsigned(24209, LUT_AMPL_WIDTH - 1),
		24098 => to_unsigned(24207, LUT_AMPL_WIDTH - 1),
		24099 => to_unsigned(24205, LUT_AMPL_WIDTH - 1),
		24100 => to_unsigned(24203, LUT_AMPL_WIDTH - 1),
		24101 => to_unsigned(24201, LUT_AMPL_WIDTH - 1),
		24102 => to_unsigned(24198, LUT_AMPL_WIDTH - 1),
		24103 => to_unsigned(24196, LUT_AMPL_WIDTH - 1),
		24104 => to_unsigned(24194, LUT_AMPL_WIDTH - 1),
		24105 => to_unsigned(24192, LUT_AMPL_WIDTH - 1),
		24106 => to_unsigned(24190, LUT_AMPL_WIDTH - 1),
		24107 => to_unsigned(24188, LUT_AMPL_WIDTH - 1),
		24108 => to_unsigned(24186, LUT_AMPL_WIDTH - 1),
		24109 => to_unsigned(24184, LUT_AMPL_WIDTH - 1),
		24110 => to_unsigned(24181, LUT_AMPL_WIDTH - 1),
		24111 => to_unsigned(24179, LUT_AMPL_WIDTH - 1),
		24112 => to_unsigned(24177, LUT_AMPL_WIDTH - 1),
		24113 => to_unsigned(24175, LUT_AMPL_WIDTH - 1),
		24114 => to_unsigned(24173, LUT_AMPL_WIDTH - 1),
		24115 => to_unsigned(24171, LUT_AMPL_WIDTH - 1),
		24116 => to_unsigned(24169, LUT_AMPL_WIDTH - 1),
		24117 => to_unsigned(24167, LUT_AMPL_WIDTH - 1),
		24118 => to_unsigned(24164, LUT_AMPL_WIDTH - 1),
		24119 => to_unsigned(24162, LUT_AMPL_WIDTH - 1),
		24120 => to_unsigned(24160, LUT_AMPL_WIDTH - 1),
		24121 => to_unsigned(24158, LUT_AMPL_WIDTH - 1),
		24122 => to_unsigned(24156, LUT_AMPL_WIDTH - 1),
		24123 => to_unsigned(24154, LUT_AMPL_WIDTH - 1),
		24124 => to_unsigned(24152, LUT_AMPL_WIDTH - 1),
		24125 => to_unsigned(24150, LUT_AMPL_WIDTH - 1),
		24126 => to_unsigned(24148, LUT_AMPL_WIDTH - 1),
		24127 => to_unsigned(24145, LUT_AMPL_WIDTH - 1),
		24128 => to_unsigned(24143, LUT_AMPL_WIDTH - 1),
		24129 => to_unsigned(24141, LUT_AMPL_WIDTH - 1),
		24130 => to_unsigned(24139, LUT_AMPL_WIDTH - 1),
		24131 => to_unsigned(24137, LUT_AMPL_WIDTH - 1),
		24132 => to_unsigned(24135, LUT_AMPL_WIDTH - 1),
		24133 => to_unsigned(24133, LUT_AMPL_WIDTH - 1),
		24134 => to_unsigned(24131, LUT_AMPL_WIDTH - 1),
		24135 => to_unsigned(24128, LUT_AMPL_WIDTH - 1),
		24136 => to_unsigned(24126, LUT_AMPL_WIDTH - 1),
		24137 => to_unsigned(24124, LUT_AMPL_WIDTH - 1),
		24138 => to_unsigned(24122, LUT_AMPL_WIDTH - 1),
		24139 => to_unsigned(24120, LUT_AMPL_WIDTH - 1),
		24140 => to_unsigned(24118, LUT_AMPL_WIDTH - 1),
		24141 => to_unsigned(24116, LUT_AMPL_WIDTH - 1),
		24142 => to_unsigned(24114, LUT_AMPL_WIDTH - 1),
		24143 => to_unsigned(24111, LUT_AMPL_WIDTH - 1),
		24144 => to_unsigned(24109, LUT_AMPL_WIDTH - 1),
		24145 => to_unsigned(24107, LUT_AMPL_WIDTH - 1),
		24146 => to_unsigned(24105, LUT_AMPL_WIDTH - 1),
		24147 => to_unsigned(24103, LUT_AMPL_WIDTH - 1),
		24148 => to_unsigned(24101, LUT_AMPL_WIDTH - 1),
		24149 => to_unsigned(24099, LUT_AMPL_WIDTH - 1),
		24150 => to_unsigned(24096, LUT_AMPL_WIDTH - 1),
		24151 => to_unsigned(24094, LUT_AMPL_WIDTH - 1),
		24152 => to_unsigned(24092, LUT_AMPL_WIDTH - 1),
		24153 => to_unsigned(24090, LUT_AMPL_WIDTH - 1),
		24154 => to_unsigned(24088, LUT_AMPL_WIDTH - 1),
		24155 => to_unsigned(24086, LUT_AMPL_WIDTH - 1),
		24156 => to_unsigned(24084, LUT_AMPL_WIDTH - 1),
		24157 => to_unsigned(24082, LUT_AMPL_WIDTH - 1),
		24158 => to_unsigned(24079, LUT_AMPL_WIDTH - 1),
		24159 => to_unsigned(24077, LUT_AMPL_WIDTH - 1),
		24160 => to_unsigned(24075, LUT_AMPL_WIDTH - 1),
		24161 => to_unsigned(24073, LUT_AMPL_WIDTH - 1),
		24162 => to_unsigned(24071, LUT_AMPL_WIDTH - 1),
		24163 => to_unsigned(24069, LUT_AMPL_WIDTH - 1),
		24164 => to_unsigned(24067, LUT_AMPL_WIDTH - 1),
		24165 => to_unsigned(24065, LUT_AMPL_WIDTH - 1),
		24166 => to_unsigned(24062, LUT_AMPL_WIDTH - 1),
		24167 => to_unsigned(24060, LUT_AMPL_WIDTH - 1),
		24168 => to_unsigned(24058, LUT_AMPL_WIDTH - 1),
		24169 => to_unsigned(24056, LUT_AMPL_WIDTH - 1),
		24170 => to_unsigned(24054, LUT_AMPL_WIDTH - 1),
		24171 => to_unsigned(24052, LUT_AMPL_WIDTH - 1),
		24172 => to_unsigned(24050, LUT_AMPL_WIDTH - 1),
		24173 => to_unsigned(24047, LUT_AMPL_WIDTH - 1),
		24174 => to_unsigned(24045, LUT_AMPL_WIDTH - 1),
		24175 => to_unsigned(24043, LUT_AMPL_WIDTH - 1),
		24176 => to_unsigned(24041, LUT_AMPL_WIDTH - 1),
		24177 => to_unsigned(24039, LUT_AMPL_WIDTH - 1),
		24178 => to_unsigned(24037, LUT_AMPL_WIDTH - 1),
		24179 => to_unsigned(24035, LUT_AMPL_WIDTH - 1),
		24180 => to_unsigned(24033, LUT_AMPL_WIDTH - 1),
		24181 => to_unsigned(24030, LUT_AMPL_WIDTH - 1),
		24182 => to_unsigned(24028, LUT_AMPL_WIDTH - 1),
		24183 => to_unsigned(24026, LUT_AMPL_WIDTH - 1),
		24184 => to_unsigned(24024, LUT_AMPL_WIDTH - 1),
		24185 => to_unsigned(24022, LUT_AMPL_WIDTH - 1),
		24186 => to_unsigned(24020, LUT_AMPL_WIDTH - 1),
		24187 => to_unsigned(24018, LUT_AMPL_WIDTH - 1),
		24188 => to_unsigned(24015, LUT_AMPL_WIDTH - 1),
		24189 => to_unsigned(24013, LUT_AMPL_WIDTH - 1),
		24190 => to_unsigned(24011, LUT_AMPL_WIDTH - 1),
		24191 => to_unsigned(24009, LUT_AMPL_WIDTH - 1),
		24192 => to_unsigned(24007, LUT_AMPL_WIDTH - 1),
		24193 => to_unsigned(24005, LUT_AMPL_WIDTH - 1),
		24194 => to_unsigned(24003, LUT_AMPL_WIDTH - 1),
		24195 => to_unsigned(24000, LUT_AMPL_WIDTH - 1),
		24196 => to_unsigned(23998, LUT_AMPL_WIDTH - 1),
		24197 => to_unsigned(23996, LUT_AMPL_WIDTH - 1),
		24198 => to_unsigned(23994, LUT_AMPL_WIDTH - 1),
		24199 => to_unsigned(23992, LUT_AMPL_WIDTH - 1),
		24200 => to_unsigned(23990, LUT_AMPL_WIDTH - 1),
		24201 => to_unsigned(23988, LUT_AMPL_WIDTH - 1),
		24202 => to_unsigned(23985, LUT_AMPL_WIDTH - 1),
		24203 => to_unsigned(23983, LUT_AMPL_WIDTH - 1),
		24204 => to_unsigned(23981, LUT_AMPL_WIDTH - 1),
		24205 => to_unsigned(23979, LUT_AMPL_WIDTH - 1),
		24206 => to_unsigned(23977, LUT_AMPL_WIDTH - 1),
		24207 => to_unsigned(23975, LUT_AMPL_WIDTH - 1),
		24208 => to_unsigned(23973, LUT_AMPL_WIDTH - 1),
		24209 => to_unsigned(23971, LUT_AMPL_WIDTH - 1),
		24210 => to_unsigned(23968, LUT_AMPL_WIDTH - 1),
		24211 => to_unsigned(23966, LUT_AMPL_WIDTH - 1),
		24212 => to_unsigned(23964, LUT_AMPL_WIDTH - 1),
		24213 => to_unsigned(23962, LUT_AMPL_WIDTH - 1),
		24214 => to_unsigned(23960, LUT_AMPL_WIDTH - 1),
		24215 => to_unsigned(23958, LUT_AMPL_WIDTH - 1),
		24216 => to_unsigned(23956, LUT_AMPL_WIDTH - 1),
		24217 => to_unsigned(23953, LUT_AMPL_WIDTH - 1),
		24218 => to_unsigned(23951, LUT_AMPL_WIDTH - 1),
		24219 => to_unsigned(23949, LUT_AMPL_WIDTH - 1),
		24220 => to_unsigned(23947, LUT_AMPL_WIDTH - 1),
		24221 => to_unsigned(23945, LUT_AMPL_WIDTH - 1),
		24222 => to_unsigned(23943, LUT_AMPL_WIDTH - 1),
		24223 => to_unsigned(23940, LUT_AMPL_WIDTH - 1),
		24224 => to_unsigned(23938, LUT_AMPL_WIDTH - 1),
		24225 => to_unsigned(23936, LUT_AMPL_WIDTH - 1),
		24226 => to_unsigned(23934, LUT_AMPL_WIDTH - 1),
		24227 => to_unsigned(23932, LUT_AMPL_WIDTH - 1),
		24228 => to_unsigned(23930, LUT_AMPL_WIDTH - 1),
		24229 => to_unsigned(23928, LUT_AMPL_WIDTH - 1),
		24230 => to_unsigned(23925, LUT_AMPL_WIDTH - 1),
		24231 => to_unsigned(23923, LUT_AMPL_WIDTH - 1),
		24232 => to_unsigned(23921, LUT_AMPL_WIDTH - 1),
		24233 => to_unsigned(23919, LUT_AMPL_WIDTH - 1),
		24234 => to_unsigned(23917, LUT_AMPL_WIDTH - 1),
		24235 => to_unsigned(23915, LUT_AMPL_WIDTH - 1),
		24236 => to_unsigned(23913, LUT_AMPL_WIDTH - 1),
		24237 => to_unsigned(23910, LUT_AMPL_WIDTH - 1),
		24238 => to_unsigned(23908, LUT_AMPL_WIDTH - 1),
		24239 => to_unsigned(23906, LUT_AMPL_WIDTH - 1),
		24240 => to_unsigned(23904, LUT_AMPL_WIDTH - 1),
		24241 => to_unsigned(23902, LUT_AMPL_WIDTH - 1),
		24242 => to_unsigned(23900, LUT_AMPL_WIDTH - 1),
		24243 => to_unsigned(23898, LUT_AMPL_WIDTH - 1),
		24244 => to_unsigned(23895, LUT_AMPL_WIDTH - 1),
		24245 => to_unsigned(23893, LUT_AMPL_WIDTH - 1),
		24246 => to_unsigned(23891, LUT_AMPL_WIDTH - 1),
		24247 => to_unsigned(23889, LUT_AMPL_WIDTH - 1),
		24248 => to_unsigned(23887, LUT_AMPL_WIDTH - 1),
		24249 => to_unsigned(23885, LUT_AMPL_WIDTH - 1),
		24250 => to_unsigned(23883, LUT_AMPL_WIDTH - 1),
		24251 => to_unsigned(23880, LUT_AMPL_WIDTH - 1),
		24252 => to_unsigned(23878, LUT_AMPL_WIDTH - 1),
		24253 => to_unsigned(23876, LUT_AMPL_WIDTH - 1),
		24254 => to_unsigned(23874, LUT_AMPL_WIDTH - 1),
		24255 => to_unsigned(23872, LUT_AMPL_WIDTH - 1),
		24256 => to_unsigned(23870, LUT_AMPL_WIDTH - 1),
		24257 => to_unsigned(23867, LUT_AMPL_WIDTH - 1),
		24258 => to_unsigned(23865, LUT_AMPL_WIDTH - 1),
		24259 => to_unsigned(23863, LUT_AMPL_WIDTH - 1),
		24260 => to_unsigned(23861, LUT_AMPL_WIDTH - 1),
		24261 => to_unsigned(23859, LUT_AMPL_WIDTH - 1),
		24262 => to_unsigned(23857, LUT_AMPL_WIDTH - 1),
		24263 => to_unsigned(23855, LUT_AMPL_WIDTH - 1),
		24264 => to_unsigned(23852, LUT_AMPL_WIDTH - 1),
		24265 => to_unsigned(23850, LUT_AMPL_WIDTH - 1),
		24266 => to_unsigned(23848, LUT_AMPL_WIDTH - 1),
		24267 => to_unsigned(23846, LUT_AMPL_WIDTH - 1),
		24268 => to_unsigned(23844, LUT_AMPL_WIDTH - 1),
		24269 => to_unsigned(23842, LUT_AMPL_WIDTH - 1),
		24270 => to_unsigned(23839, LUT_AMPL_WIDTH - 1),
		24271 => to_unsigned(23837, LUT_AMPL_WIDTH - 1),
		24272 => to_unsigned(23835, LUT_AMPL_WIDTH - 1),
		24273 => to_unsigned(23833, LUT_AMPL_WIDTH - 1),
		24274 => to_unsigned(23831, LUT_AMPL_WIDTH - 1),
		24275 => to_unsigned(23829, LUT_AMPL_WIDTH - 1),
		24276 => to_unsigned(23827, LUT_AMPL_WIDTH - 1),
		24277 => to_unsigned(23824, LUT_AMPL_WIDTH - 1),
		24278 => to_unsigned(23822, LUT_AMPL_WIDTH - 1),
		24279 => to_unsigned(23820, LUT_AMPL_WIDTH - 1),
		24280 => to_unsigned(23818, LUT_AMPL_WIDTH - 1),
		24281 => to_unsigned(23816, LUT_AMPL_WIDTH - 1),
		24282 => to_unsigned(23814, LUT_AMPL_WIDTH - 1),
		24283 => to_unsigned(23811, LUT_AMPL_WIDTH - 1),
		24284 => to_unsigned(23809, LUT_AMPL_WIDTH - 1),
		24285 => to_unsigned(23807, LUT_AMPL_WIDTH - 1),
		24286 => to_unsigned(23805, LUT_AMPL_WIDTH - 1),
		24287 => to_unsigned(23803, LUT_AMPL_WIDTH - 1),
		24288 => to_unsigned(23801, LUT_AMPL_WIDTH - 1),
		24289 => to_unsigned(23798, LUT_AMPL_WIDTH - 1),
		24290 => to_unsigned(23796, LUT_AMPL_WIDTH - 1),
		24291 => to_unsigned(23794, LUT_AMPL_WIDTH - 1),
		24292 => to_unsigned(23792, LUT_AMPL_WIDTH - 1),
		24293 => to_unsigned(23790, LUT_AMPL_WIDTH - 1),
		24294 => to_unsigned(23788, LUT_AMPL_WIDTH - 1),
		24295 => to_unsigned(23785, LUT_AMPL_WIDTH - 1),
		24296 => to_unsigned(23783, LUT_AMPL_WIDTH - 1),
		24297 => to_unsigned(23781, LUT_AMPL_WIDTH - 1),
		24298 => to_unsigned(23779, LUT_AMPL_WIDTH - 1),
		24299 => to_unsigned(23777, LUT_AMPL_WIDTH - 1),
		24300 => to_unsigned(23775, LUT_AMPL_WIDTH - 1),
		24301 => to_unsigned(23773, LUT_AMPL_WIDTH - 1),
		24302 => to_unsigned(23770, LUT_AMPL_WIDTH - 1),
		24303 => to_unsigned(23768, LUT_AMPL_WIDTH - 1),
		24304 => to_unsigned(23766, LUT_AMPL_WIDTH - 1),
		24305 => to_unsigned(23764, LUT_AMPL_WIDTH - 1),
		24306 => to_unsigned(23762, LUT_AMPL_WIDTH - 1),
		24307 => to_unsigned(23760, LUT_AMPL_WIDTH - 1),
		24308 => to_unsigned(23757, LUT_AMPL_WIDTH - 1),
		24309 => to_unsigned(23755, LUT_AMPL_WIDTH - 1),
		24310 => to_unsigned(23753, LUT_AMPL_WIDTH - 1),
		24311 => to_unsigned(23751, LUT_AMPL_WIDTH - 1),
		24312 => to_unsigned(23749, LUT_AMPL_WIDTH - 1),
		24313 => to_unsigned(23747, LUT_AMPL_WIDTH - 1),
		24314 => to_unsigned(23744, LUT_AMPL_WIDTH - 1),
		24315 => to_unsigned(23742, LUT_AMPL_WIDTH - 1),
		24316 => to_unsigned(23740, LUT_AMPL_WIDTH - 1),
		24317 => to_unsigned(23738, LUT_AMPL_WIDTH - 1),
		24318 => to_unsigned(23736, LUT_AMPL_WIDTH - 1),
		24319 => to_unsigned(23734, LUT_AMPL_WIDTH - 1),
		24320 => to_unsigned(23731, LUT_AMPL_WIDTH - 1),
		24321 => to_unsigned(23729, LUT_AMPL_WIDTH - 1),
		24322 => to_unsigned(23727, LUT_AMPL_WIDTH - 1),
		24323 => to_unsigned(23725, LUT_AMPL_WIDTH - 1),
		24324 => to_unsigned(23723, LUT_AMPL_WIDTH - 1),
		24325 => to_unsigned(23721, LUT_AMPL_WIDTH - 1),
		24326 => to_unsigned(23718, LUT_AMPL_WIDTH - 1),
		24327 => to_unsigned(23716, LUT_AMPL_WIDTH - 1),
		24328 => to_unsigned(23714, LUT_AMPL_WIDTH - 1),
		24329 => to_unsigned(23712, LUT_AMPL_WIDTH - 1),
		24330 => to_unsigned(23710, LUT_AMPL_WIDTH - 1),
		24331 => to_unsigned(23708, LUT_AMPL_WIDTH - 1),
		24332 => to_unsigned(23705, LUT_AMPL_WIDTH - 1),
		24333 => to_unsigned(23703, LUT_AMPL_WIDTH - 1),
		24334 => to_unsigned(23701, LUT_AMPL_WIDTH - 1),
		24335 => to_unsigned(23699, LUT_AMPL_WIDTH - 1),
		24336 => to_unsigned(23697, LUT_AMPL_WIDTH - 1),
		24337 => to_unsigned(23695, LUT_AMPL_WIDTH - 1),
		24338 => to_unsigned(23692, LUT_AMPL_WIDTH - 1),
		24339 => to_unsigned(23690, LUT_AMPL_WIDTH - 1),
		24340 => to_unsigned(23688, LUT_AMPL_WIDTH - 1),
		24341 => to_unsigned(23686, LUT_AMPL_WIDTH - 1),
		24342 => to_unsigned(23684, LUT_AMPL_WIDTH - 1),
		24343 => to_unsigned(23682, LUT_AMPL_WIDTH - 1),
		24344 => to_unsigned(23679, LUT_AMPL_WIDTH - 1),
		24345 => to_unsigned(23677, LUT_AMPL_WIDTH - 1),
		24346 => to_unsigned(23675, LUT_AMPL_WIDTH - 1),
		24347 => to_unsigned(23673, LUT_AMPL_WIDTH - 1),
		24348 => to_unsigned(23671, LUT_AMPL_WIDTH - 1),
		24349 => to_unsigned(23668, LUT_AMPL_WIDTH - 1),
		24350 => to_unsigned(23666, LUT_AMPL_WIDTH - 1),
		24351 => to_unsigned(23664, LUT_AMPL_WIDTH - 1),
		24352 => to_unsigned(23662, LUT_AMPL_WIDTH - 1),
		24353 => to_unsigned(23660, LUT_AMPL_WIDTH - 1),
		24354 => to_unsigned(23658, LUT_AMPL_WIDTH - 1),
		24355 => to_unsigned(23655, LUT_AMPL_WIDTH - 1),
		24356 => to_unsigned(23653, LUT_AMPL_WIDTH - 1),
		24357 => to_unsigned(23651, LUT_AMPL_WIDTH - 1),
		24358 => to_unsigned(23649, LUT_AMPL_WIDTH - 1),
		24359 => to_unsigned(23647, LUT_AMPL_WIDTH - 1),
		24360 => to_unsigned(23645, LUT_AMPL_WIDTH - 1),
		24361 => to_unsigned(23642, LUT_AMPL_WIDTH - 1),
		24362 => to_unsigned(23640, LUT_AMPL_WIDTH - 1),
		24363 => to_unsigned(23638, LUT_AMPL_WIDTH - 1),
		24364 => to_unsigned(23636, LUT_AMPL_WIDTH - 1),
		24365 => to_unsigned(23634, LUT_AMPL_WIDTH - 1),
		24366 => to_unsigned(23632, LUT_AMPL_WIDTH - 1),
		24367 => to_unsigned(23629, LUT_AMPL_WIDTH - 1),
		24368 => to_unsigned(23627, LUT_AMPL_WIDTH - 1),
		24369 => to_unsigned(23625, LUT_AMPL_WIDTH - 1),
		24370 => to_unsigned(23623, LUT_AMPL_WIDTH - 1),
		24371 => to_unsigned(23621, LUT_AMPL_WIDTH - 1),
		24372 => to_unsigned(23618, LUT_AMPL_WIDTH - 1),
		24373 => to_unsigned(23616, LUT_AMPL_WIDTH - 1),
		24374 => to_unsigned(23614, LUT_AMPL_WIDTH - 1),
		24375 => to_unsigned(23612, LUT_AMPL_WIDTH - 1),
		24376 => to_unsigned(23610, LUT_AMPL_WIDTH - 1),
		24377 => to_unsigned(23608, LUT_AMPL_WIDTH - 1),
		24378 => to_unsigned(23605, LUT_AMPL_WIDTH - 1),
		24379 => to_unsigned(23603, LUT_AMPL_WIDTH - 1),
		24380 => to_unsigned(23601, LUT_AMPL_WIDTH - 1),
		24381 => to_unsigned(23599, LUT_AMPL_WIDTH - 1),
		24382 => to_unsigned(23597, LUT_AMPL_WIDTH - 1),
		24383 => to_unsigned(23595, LUT_AMPL_WIDTH - 1),
		24384 => to_unsigned(23592, LUT_AMPL_WIDTH - 1),
		24385 => to_unsigned(23590, LUT_AMPL_WIDTH - 1),
		24386 => to_unsigned(23588, LUT_AMPL_WIDTH - 1),
		24387 => to_unsigned(23586, LUT_AMPL_WIDTH - 1),
		24388 => to_unsigned(23584, LUT_AMPL_WIDTH - 1),
		24389 => to_unsigned(23581, LUT_AMPL_WIDTH - 1),
		24390 => to_unsigned(23579, LUT_AMPL_WIDTH - 1),
		24391 => to_unsigned(23577, LUT_AMPL_WIDTH - 1),
		24392 => to_unsigned(23575, LUT_AMPL_WIDTH - 1),
		24393 => to_unsigned(23573, LUT_AMPL_WIDTH - 1),
		24394 => to_unsigned(23571, LUT_AMPL_WIDTH - 1),
		24395 => to_unsigned(23568, LUT_AMPL_WIDTH - 1),
		24396 => to_unsigned(23566, LUT_AMPL_WIDTH - 1),
		24397 => to_unsigned(23564, LUT_AMPL_WIDTH - 1),
		24398 => to_unsigned(23562, LUT_AMPL_WIDTH - 1),
		24399 => to_unsigned(23560, LUT_AMPL_WIDTH - 1),
		24400 => to_unsigned(23557, LUT_AMPL_WIDTH - 1),
		24401 => to_unsigned(23555, LUT_AMPL_WIDTH - 1),
		24402 => to_unsigned(23553, LUT_AMPL_WIDTH - 1),
		24403 => to_unsigned(23551, LUT_AMPL_WIDTH - 1),
		24404 => to_unsigned(23549, LUT_AMPL_WIDTH - 1),
		24405 => to_unsigned(23546, LUT_AMPL_WIDTH - 1),
		24406 => to_unsigned(23544, LUT_AMPL_WIDTH - 1),
		24407 => to_unsigned(23542, LUT_AMPL_WIDTH - 1),
		24408 => to_unsigned(23540, LUT_AMPL_WIDTH - 1),
		24409 => to_unsigned(23538, LUT_AMPL_WIDTH - 1),
		24410 => to_unsigned(23536, LUT_AMPL_WIDTH - 1),
		24411 => to_unsigned(23533, LUT_AMPL_WIDTH - 1),
		24412 => to_unsigned(23531, LUT_AMPL_WIDTH - 1),
		24413 => to_unsigned(23529, LUT_AMPL_WIDTH - 1),
		24414 => to_unsigned(23527, LUT_AMPL_WIDTH - 1),
		24415 => to_unsigned(23525, LUT_AMPL_WIDTH - 1),
		24416 => to_unsigned(23522, LUT_AMPL_WIDTH - 1),
		24417 => to_unsigned(23520, LUT_AMPL_WIDTH - 1),
		24418 => to_unsigned(23518, LUT_AMPL_WIDTH - 1),
		24419 => to_unsigned(23516, LUT_AMPL_WIDTH - 1),
		24420 => to_unsigned(23514, LUT_AMPL_WIDTH - 1),
		24421 => to_unsigned(23512, LUT_AMPL_WIDTH - 1),
		24422 => to_unsigned(23509, LUT_AMPL_WIDTH - 1),
		24423 => to_unsigned(23507, LUT_AMPL_WIDTH - 1),
		24424 => to_unsigned(23505, LUT_AMPL_WIDTH - 1),
		24425 => to_unsigned(23503, LUT_AMPL_WIDTH - 1),
		24426 => to_unsigned(23501, LUT_AMPL_WIDTH - 1),
		24427 => to_unsigned(23498, LUT_AMPL_WIDTH - 1),
		24428 => to_unsigned(23496, LUT_AMPL_WIDTH - 1),
		24429 => to_unsigned(23494, LUT_AMPL_WIDTH - 1),
		24430 => to_unsigned(23492, LUT_AMPL_WIDTH - 1),
		24431 => to_unsigned(23490, LUT_AMPL_WIDTH - 1),
		24432 => to_unsigned(23487, LUT_AMPL_WIDTH - 1),
		24433 => to_unsigned(23485, LUT_AMPL_WIDTH - 1),
		24434 => to_unsigned(23483, LUT_AMPL_WIDTH - 1),
		24435 => to_unsigned(23481, LUT_AMPL_WIDTH - 1),
		24436 => to_unsigned(23479, LUT_AMPL_WIDTH - 1),
		24437 => to_unsigned(23476, LUT_AMPL_WIDTH - 1),
		24438 => to_unsigned(23474, LUT_AMPL_WIDTH - 1),
		24439 => to_unsigned(23472, LUT_AMPL_WIDTH - 1),
		24440 => to_unsigned(23470, LUT_AMPL_WIDTH - 1),
		24441 => to_unsigned(23468, LUT_AMPL_WIDTH - 1),
		24442 => to_unsigned(23466, LUT_AMPL_WIDTH - 1),
		24443 => to_unsigned(23463, LUT_AMPL_WIDTH - 1),
		24444 => to_unsigned(23461, LUT_AMPL_WIDTH - 1),
		24445 => to_unsigned(23459, LUT_AMPL_WIDTH - 1),
		24446 => to_unsigned(23457, LUT_AMPL_WIDTH - 1),
		24447 => to_unsigned(23455, LUT_AMPL_WIDTH - 1),
		24448 => to_unsigned(23452, LUT_AMPL_WIDTH - 1),
		24449 => to_unsigned(23450, LUT_AMPL_WIDTH - 1),
		24450 => to_unsigned(23448, LUT_AMPL_WIDTH - 1),
		24451 => to_unsigned(23446, LUT_AMPL_WIDTH - 1),
		24452 => to_unsigned(23444, LUT_AMPL_WIDTH - 1),
		24453 => to_unsigned(23441, LUT_AMPL_WIDTH - 1),
		24454 => to_unsigned(23439, LUT_AMPL_WIDTH - 1),
		24455 => to_unsigned(23437, LUT_AMPL_WIDTH - 1),
		24456 => to_unsigned(23435, LUT_AMPL_WIDTH - 1),
		24457 => to_unsigned(23433, LUT_AMPL_WIDTH - 1),
		24458 => to_unsigned(23430, LUT_AMPL_WIDTH - 1),
		24459 => to_unsigned(23428, LUT_AMPL_WIDTH - 1),
		24460 => to_unsigned(23426, LUT_AMPL_WIDTH - 1),
		24461 => to_unsigned(23424, LUT_AMPL_WIDTH - 1),
		24462 => to_unsigned(23422, LUT_AMPL_WIDTH - 1),
		24463 => to_unsigned(23419, LUT_AMPL_WIDTH - 1),
		24464 => to_unsigned(23417, LUT_AMPL_WIDTH - 1),
		24465 => to_unsigned(23415, LUT_AMPL_WIDTH - 1),
		24466 => to_unsigned(23413, LUT_AMPL_WIDTH - 1),
		24467 => to_unsigned(23411, LUT_AMPL_WIDTH - 1),
		24468 => to_unsigned(23408, LUT_AMPL_WIDTH - 1),
		24469 => to_unsigned(23406, LUT_AMPL_WIDTH - 1),
		24470 => to_unsigned(23404, LUT_AMPL_WIDTH - 1),
		24471 => to_unsigned(23402, LUT_AMPL_WIDTH - 1),
		24472 => to_unsigned(23400, LUT_AMPL_WIDTH - 1),
		24473 => to_unsigned(23397, LUT_AMPL_WIDTH - 1),
		24474 => to_unsigned(23395, LUT_AMPL_WIDTH - 1),
		24475 => to_unsigned(23393, LUT_AMPL_WIDTH - 1),
		24476 => to_unsigned(23391, LUT_AMPL_WIDTH - 1),
		24477 => to_unsigned(23389, LUT_AMPL_WIDTH - 1),
		24478 => to_unsigned(23386, LUT_AMPL_WIDTH - 1),
		24479 => to_unsigned(23384, LUT_AMPL_WIDTH - 1),
		24480 => to_unsigned(23382, LUT_AMPL_WIDTH - 1),
		24481 => to_unsigned(23380, LUT_AMPL_WIDTH - 1),
		24482 => to_unsigned(23378, LUT_AMPL_WIDTH - 1),
		24483 => to_unsigned(23375, LUT_AMPL_WIDTH - 1),
		24484 => to_unsigned(23373, LUT_AMPL_WIDTH - 1),
		24485 => to_unsigned(23371, LUT_AMPL_WIDTH - 1),
		24486 => to_unsigned(23369, LUT_AMPL_WIDTH - 1),
		24487 => to_unsigned(23367, LUT_AMPL_WIDTH - 1),
		24488 => to_unsigned(23364, LUT_AMPL_WIDTH - 1),
		24489 => to_unsigned(23362, LUT_AMPL_WIDTH - 1),
		24490 => to_unsigned(23360, LUT_AMPL_WIDTH - 1),
		24491 => to_unsigned(23358, LUT_AMPL_WIDTH - 1),
		24492 => to_unsigned(23356, LUT_AMPL_WIDTH - 1),
		24493 => to_unsigned(23353, LUT_AMPL_WIDTH - 1),
		24494 => to_unsigned(23351, LUT_AMPL_WIDTH - 1),
		24495 => to_unsigned(23349, LUT_AMPL_WIDTH - 1),
		24496 => to_unsigned(23347, LUT_AMPL_WIDTH - 1),
		24497 => to_unsigned(23345, LUT_AMPL_WIDTH - 1),
		24498 => to_unsigned(23342, LUT_AMPL_WIDTH - 1),
		24499 => to_unsigned(23340, LUT_AMPL_WIDTH - 1),
		24500 => to_unsigned(23338, LUT_AMPL_WIDTH - 1),
		24501 => to_unsigned(23336, LUT_AMPL_WIDTH - 1),
		24502 => to_unsigned(23334, LUT_AMPL_WIDTH - 1),
		24503 => to_unsigned(23331, LUT_AMPL_WIDTH - 1),
		24504 => to_unsigned(23329, LUT_AMPL_WIDTH - 1),
		24505 => to_unsigned(23327, LUT_AMPL_WIDTH - 1),
		24506 => to_unsigned(23325, LUT_AMPL_WIDTH - 1),
		24507 => to_unsigned(23323, LUT_AMPL_WIDTH - 1),
		24508 => to_unsigned(23320, LUT_AMPL_WIDTH - 1),
		24509 => to_unsigned(23318, LUT_AMPL_WIDTH - 1),
		24510 => to_unsigned(23316, LUT_AMPL_WIDTH - 1),
		24511 => to_unsigned(23314, LUT_AMPL_WIDTH - 1),
		24512 => to_unsigned(23311, LUT_AMPL_WIDTH - 1),
		24513 => to_unsigned(23309, LUT_AMPL_WIDTH - 1),
		24514 => to_unsigned(23307, LUT_AMPL_WIDTH - 1),
		24515 => to_unsigned(23305, LUT_AMPL_WIDTH - 1),
		24516 => to_unsigned(23303, LUT_AMPL_WIDTH - 1),
		24517 => to_unsigned(23300, LUT_AMPL_WIDTH - 1),
		24518 => to_unsigned(23298, LUT_AMPL_WIDTH - 1),
		24519 => to_unsigned(23296, LUT_AMPL_WIDTH - 1),
		24520 => to_unsigned(23294, LUT_AMPL_WIDTH - 1),
		24521 => to_unsigned(23292, LUT_AMPL_WIDTH - 1),
		24522 => to_unsigned(23289, LUT_AMPL_WIDTH - 1),
		24523 => to_unsigned(23287, LUT_AMPL_WIDTH - 1),
		24524 => to_unsigned(23285, LUT_AMPL_WIDTH - 1),
		24525 => to_unsigned(23283, LUT_AMPL_WIDTH - 1),
		24526 => to_unsigned(23281, LUT_AMPL_WIDTH - 1),
		24527 => to_unsigned(23278, LUT_AMPL_WIDTH - 1),
		24528 => to_unsigned(23276, LUT_AMPL_WIDTH - 1),
		24529 => to_unsigned(23274, LUT_AMPL_WIDTH - 1),
		24530 => to_unsigned(23272, LUT_AMPL_WIDTH - 1),
		24531 => to_unsigned(23270, LUT_AMPL_WIDTH - 1),
		24532 => to_unsigned(23267, LUT_AMPL_WIDTH - 1),
		24533 => to_unsigned(23265, LUT_AMPL_WIDTH - 1),
		24534 => to_unsigned(23263, LUT_AMPL_WIDTH - 1),
		24535 => to_unsigned(23261, LUT_AMPL_WIDTH - 1),
		24536 => to_unsigned(23258, LUT_AMPL_WIDTH - 1),
		24537 => to_unsigned(23256, LUT_AMPL_WIDTH - 1),
		24538 => to_unsigned(23254, LUT_AMPL_WIDTH - 1),
		24539 => to_unsigned(23252, LUT_AMPL_WIDTH - 1),
		24540 => to_unsigned(23250, LUT_AMPL_WIDTH - 1),
		24541 => to_unsigned(23247, LUT_AMPL_WIDTH - 1),
		24542 => to_unsigned(23245, LUT_AMPL_WIDTH - 1),
		24543 => to_unsigned(23243, LUT_AMPL_WIDTH - 1),
		24544 => to_unsigned(23241, LUT_AMPL_WIDTH - 1),
		24545 => to_unsigned(23239, LUT_AMPL_WIDTH - 1),
		24546 => to_unsigned(23236, LUT_AMPL_WIDTH - 1),
		24547 => to_unsigned(23234, LUT_AMPL_WIDTH - 1),
		24548 => to_unsigned(23232, LUT_AMPL_WIDTH - 1),
		24549 => to_unsigned(23230, LUT_AMPL_WIDTH - 1),
		24550 => to_unsigned(23227, LUT_AMPL_WIDTH - 1),
		24551 => to_unsigned(23225, LUT_AMPL_WIDTH - 1),
		24552 => to_unsigned(23223, LUT_AMPL_WIDTH - 1),
		24553 => to_unsigned(23221, LUT_AMPL_WIDTH - 1),
		24554 => to_unsigned(23219, LUT_AMPL_WIDTH - 1),
		24555 => to_unsigned(23216, LUT_AMPL_WIDTH - 1),
		24556 => to_unsigned(23214, LUT_AMPL_WIDTH - 1),
		24557 => to_unsigned(23212, LUT_AMPL_WIDTH - 1),
		24558 => to_unsigned(23210, LUT_AMPL_WIDTH - 1),
		24559 => to_unsigned(23208, LUT_AMPL_WIDTH - 1),
		24560 => to_unsigned(23205, LUT_AMPL_WIDTH - 1),
		24561 => to_unsigned(23203, LUT_AMPL_WIDTH - 1),
		24562 => to_unsigned(23201, LUT_AMPL_WIDTH - 1),
		24563 => to_unsigned(23199, LUT_AMPL_WIDTH - 1),
		24564 => to_unsigned(23196, LUT_AMPL_WIDTH - 1),
		24565 => to_unsigned(23194, LUT_AMPL_WIDTH - 1),
		24566 => to_unsigned(23192, LUT_AMPL_WIDTH - 1),
		24567 => to_unsigned(23190, LUT_AMPL_WIDTH - 1),
		24568 => to_unsigned(23188, LUT_AMPL_WIDTH - 1),
		24569 => to_unsigned(23185, LUT_AMPL_WIDTH - 1),
		24570 => to_unsigned(23183, LUT_AMPL_WIDTH - 1),
		24571 => to_unsigned(23181, LUT_AMPL_WIDTH - 1),
		24572 => to_unsigned(23179, LUT_AMPL_WIDTH - 1),
		24573 => to_unsigned(23176, LUT_AMPL_WIDTH - 1),
		24574 => to_unsigned(23174, LUT_AMPL_WIDTH - 1),
		24575 => to_unsigned(23172, LUT_AMPL_WIDTH - 1),
		24576 => to_unsigned(23170, LUT_AMPL_WIDTH - 1),
		24577 => to_unsigned(23168, LUT_AMPL_WIDTH - 1),
		24578 => to_unsigned(23165, LUT_AMPL_WIDTH - 1),
		24579 => to_unsigned(23163, LUT_AMPL_WIDTH - 1),
		24580 => to_unsigned(23161, LUT_AMPL_WIDTH - 1),
		24581 => to_unsigned(23159, LUT_AMPL_WIDTH - 1),
		24582 => to_unsigned(23156, LUT_AMPL_WIDTH - 1),
		24583 => to_unsigned(23154, LUT_AMPL_WIDTH - 1),
		24584 => to_unsigned(23152, LUT_AMPL_WIDTH - 1),
		24585 => to_unsigned(23150, LUT_AMPL_WIDTH - 1),
		24586 => to_unsigned(23148, LUT_AMPL_WIDTH - 1),
		24587 => to_unsigned(23145, LUT_AMPL_WIDTH - 1),
		24588 => to_unsigned(23143, LUT_AMPL_WIDTH - 1),
		24589 => to_unsigned(23141, LUT_AMPL_WIDTH - 1),
		24590 => to_unsigned(23139, LUT_AMPL_WIDTH - 1),
		24591 => to_unsigned(23136, LUT_AMPL_WIDTH - 1),
		24592 => to_unsigned(23134, LUT_AMPL_WIDTH - 1),
		24593 => to_unsigned(23132, LUT_AMPL_WIDTH - 1),
		24594 => to_unsigned(23130, LUT_AMPL_WIDTH - 1),
		24595 => to_unsigned(23128, LUT_AMPL_WIDTH - 1),
		24596 => to_unsigned(23125, LUT_AMPL_WIDTH - 1),
		24597 => to_unsigned(23123, LUT_AMPL_WIDTH - 1),
		24598 => to_unsigned(23121, LUT_AMPL_WIDTH - 1),
		24599 => to_unsigned(23119, LUT_AMPL_WIDTH - 1),
		24600 => to_unsigned(23116, LUT_AMPL_WIDTH - 1),
		24601 => to_unsigned(23114, LUT_AMPL_WIDTH - 1),
		24602 => to_unsigned(23112, LUT_AMPL_WIDTH - 1),
		24603 => to_unsigned(23110, LUT_AMPL_WIDTH - 1),
		24604 => to_unsigned(23107, LUT_AMPL_WIDTH - 1),
		24605 => to_unsigned(23105, LUT_AMPL_WIDTH - 1),
		24606 => to_unsigned(23103, LUT_AMPL_WIDTH - 1),
		24607 => to_unsigned(23101, LUT_AMPL_WIDTH - 1),
		24608 => to_unsigned(23099, LUT_AMPL_WIDTH - 1),
		24609 => to_unsigned(23096, LUT_AMPL_WIDTH - 1),
		24610 => to_unsigned(23094, LUT_AMPL_WIDTH - 1),
		24611 => to_unsigned(23092, LUT_AMPL_WIDTH - 1),
		24612 => to_unsigned(23090, LUT_AMPL_WIDTH - 1),
		24613 => to_unsigned(23087, LUT_AMPL_WIDTH - 1),
		24614 => to_unsigned(23085, LUT_AMPL_WIDTH - 1),
		24615 => to_unsigned(23083, LUT_AMPL_WIDTH - 1),
		24616 => to_unsigned(23081, LUT_AMPL_WIDTH - 1),
		24617 => to_unsigned(23079, LUT_AMPL_WIDTH - 1),
		24618 => to_unsigned(23076, LUT_AMPL_WIDTH - 1),
		24619 => to_unsigned(23074, LUT_AMPL_WIDTH - 1),
		24620 => to_unsigned(23072, LUT_AMPL_WIDTH - 1),
		24621 => to_unsigned(23070, LUT_AMPL_WIDTH - 1),
		24622 => to_unsigned(23067, LUT_AMPL_WIDTH - 1),
		24623 => to_unsigned(23065, LUT_AMPL_WIDTH - 1),
		24624 => to_unsigned(23063, LUT_AMPL_WIDTH - 1),
		24625 => to_unsigned(23061, LUT_AMPL_WIDTH - 1),
		24626 => to_unsigned(23058, LUT_AMPL_WIDTH - 1),
		24627 => to_unsigned(23056, LUT_AMPL_WIDTH - 1),
		24628 => to_unsigned(23054, LUT_AMPL_WIDTH - 1),
		24629 => to_unsigned(23052, LUT_AMPL_WIDTH - 1),
		24630 => to_unsigned(23050, LUT_AMPL_WIDTH - 1),
		24631 => to_unsigned(23047, LUT_AMPL_WIDTH - 1),
		24632 => to_unsigned(23045, LUT_AMPL_WIDTH - 1),
		24633 => to_unsigned(23043, LUT_AMPL_WIDTH - 1),
		24634 => to_unsigned(23041, LUT_AMPL_WIDTH - 1),
		24635 => to_unsigned(23038, LUT_AMPL_WIDTH - 1),
		24636 => to_unsigned(23036, LUT_AMPL_WIDTH - 1),
		24637 => to_unsigned(23034, LUT_AMPL_WIDTH - 1),
		24638 => to_unsigned(23032, LUT_AMPL_WIDTH - 1),
		24639 => to_unsigned(23029, LUT_AMPL_WIDTH - 1),
		24640 => to_unsigned(23027, LUT_AMPL_WIDTH - 1),
		24641 => to_unsigned(23025, LUT_AMPL_WIDTH - 1),
		24642 => to_unsigned(23023, LUT_AMPL_WIDTH - 1),
		24643 => to_unsigned(23020, LUT_AMPL_WIDTH - 1),
		24644 => to_unsigned(23018, LUT_AMPL_WIDTH - 1),
		24645 => to_unsigned(23016, LUT_AMPL_WIDTH - 1),
		24646 => to_unsigned(23014, LUT_AMPL_WIDTH - 1),
		24647 => to_unsigned(23012, LUT_AMPL_WIDTH - 1),
		24648 => to_unsigned(23009, LUT_AMPL_WIDTH - 1),
		24649 => to_unsigned(23007, LUT_AMPL_WIDTH - 1),
		24650 => to_unsigned(23005, LUT_AMPL_WIDTH - 1),
		24651 => to_unsigned(23003, LUT_AMPL_WIDTH - 1),
		24652 => to_unsigned(23000, LUT_AMPL_WIDTH - 1),
		24653 => to_unsigned(22998, LUT_AMPL_WIDTH - 1),
		24654 => to_unsigned(22996, LUT_AMPL_WIDTH - 1),
		24655 => to_unsigned(22994, LUT_AMPL_WIDTH - 1),
		24656 => to_unsigned(22991, LUT_AMPL_WIDTH - 1),
		24657 => to_unsigned(22989, LUT_AMPL_WIDTH - 1),
		24658 => to_unsigned(22987, LUT_AMPL_WIDTH - 1),
		24659 => to_unsigned(22985, LUT_AMPL_WIDTH - 1),
		24660 => to_unsigned(22982, LUT_AMPL_WIDTH - 1),
		24661 => to_unsigned(22980, LUT_AMPL_WIDTH - 1),
		24662 => to_unsigned(22978, LUT_AMPL_WIDTH - 1),
		24663 => to_unsigned(22976, LUT_AMPL_WIDTH - 1),
		24664 => to_unsigned(22973, LUT_AMPL_WIDTH - 1),
		24665 => to_unsigned(22971, LUT_AMPL_WIDTH - 1),
		24666 => to_unsigned(22969, LUT_AMPL_WIDTH - 1),
		24667 => to_unsigned(22967, LUT_AMPL_WIDTH - 1),
		24668 => to_unsigned(22965, LUT_AMPL_WIDTH - 1),
		24669 => to_unsigned(22962, LUT_AMPL_WIDTH - 1),
		24670 => to_unsigned(22960, LUT_AMPL_WIDTH - 1),
		24671 => to_unsigned(22958, LUT_AMPL_WIDTH - 1),
		24672 => to_unsigned(22956, LUT_AMPL_WIDTH - 1),
		24673 => to_unsigned(22953, LUT_AMPL_WIDTH - 1),
		24674 => to_unsigned(22951, LUT_AMPL_WIDTH - 1),
		24675 => to_unsigned(22949, LUT_AMPL_WIDTH - 1),
		24676 => to_unsigned(22947, LUT_AMPL_WIDTH - 1),
		24677 => to_unsigned(22944, LUT_AMPL_WIDTH - 1),
		24678 => to_unsigned(22942, LUT_AMPL_WIDTH - 1),
		24679 => to_unsigned(22940, LUT_AMPL_WIDTH - 1),
		24680 => to_unsigned(22938, LUT_AMPL_WIDTH - 1),
		24681 => to_unsigned(22935, LUT_AMPL_WIDTH - 1),
		24682 => to_unsigned(22933, LUT_AMPL_WIDTH - 1),
		24683 => to_unsigned(22931, LUT_AMPL_WIDTH - 1),
		24684 => to_unsigned(22929, LUT_AMPL_WIDTH - 1),
		24685 => to_unsigned(22926, LUT_AMPL_WIDTH - 1),
		24686 => to_unsigned(22924, LUT_AMPL_WIDTH - 1),
		24687 => to_unsigned(22922, LUT_AMPL_WIDTH - 1),
		24688 => to_unsigned(22920, LUT_AMPL_WIDTH - 1),
		24689 => to_unsigned(22917, LUT_AMPL_WIDTH - 1),
		24690 => to_unsigned(22915, LUT_AMPL_WIDTH - 1),
		24691 => to_unsigned(22913, LUT_AMPL_WIDTH - 1),
		24692 => to_unsigned(22911, LUT_AMPL_WIDTH - 1),
		24693 => to_unsigned(22908, LUT_AMPL_WIDTH - 1),
		24694 => to_unsigned(22906, LUT_AMPL_WIDTH - 1),
		24695 => to_unsigned(22904, LUT_AMPL_WIDTH - 1),
		24696 => to_unsigned(22902, LUT_AMPL_WIDTH - 1),
		24697 => to_unsigned(22899, LUT_AMPL_WIDTH - 1),
		24698 => to_unsigned(22897, LUT_AMPL_WIDTH - 1),
		24699 => to_unsigned(22895, LUT_AMPL_WIDTH - 1),
		24700 => to_unsigned(22893, LUT_AMPL_WIDTH - 1),
		24701 => to_unsigned(22890, LUT_AMPL_WIDTH - 1),
		24702 => to_unsigned(22888, LUT_AMPL_WIDTH - 1),
		24703 => to_unsigned(22886, LUT_AMPL_WIDTH - 1),
		24704 => to_unsigned(22884, LUT_AMPL_WIDTH - 1),
		24705 => to_unsigned(22881, LUT_AMPL_WIDTH - 1),
		24706 => to_unsigned(22879, LUT_AMPL_WIDTH - 1),
		24707 => to_unsigned(22877, LUT_AMPL_WIDTH - 1),
		24708 => to_unsigned(22875, LUT_AMPL_WIDTH - 1),
		24709 => to_unsigned(22872, LUT_AMPL_WIDTH - 1),
		24710 => to_unsigned(22870, LUT_AMPL_WIDTH - 1),
		24711 => to_unsigned(22868, LUT_AMPL_WIDTH - 1),
		24712 => to_unsigned(22866, LUT_AMPL_WIDTH - 1),
		24713 => to_unsigned(22863, LUT_AMPL_WIDTH - 1),
		24714 => to_unsigned(22861, LUT_AMPL_WIDTH - 1),
		24715 => to_unsigned(22859, LUT_AMPL_WIDTH - 1),
		24716 => to_unsigned(22857, LUT_AMPL_WIDTH - 1),
		24717 => to_unsigned(22854, LUT_AMPL_WIDTH - 1),
		24718 => to_unsigned(22852, LUT_AMPL_WIDTH - 1),
		24719 => to_unsigned(22850, LUT_AMPL_WIDTH - 1),
		24720 => to_unsigned(22848, LUT_AMPL_WIDTH - 1),
		24721 => to_unsigned(22845, LUT_AMPL_WIDTH - 1),
		24722 => to_unsigned(22843, LUT_AMPL_WIDTH - 1),
		24723 => to_unsigned(22841, LUT_AMPL_WIDTH - 1),
		24724 => to_unsigned(22839, LUT_AMPL_WIDTH - 1),
		24725 => to_unsigned(22836, LUT_AMPL_WIDTH - 1),
		24726 => to_unsigned(22834, LUT_AMPL_WIDTH - 1),
		24727 => to_unsigned(22832, LUT_AMPL_WIDTH - 1),
		24728 => to_unsigned(22830, LUT_AMPL_WIDTH - 1),
		24729 => to_unsigned(22827, LUT_AMPL_WIDTH - 1),
		24730 => to_unsigned(22825, LUT_AMPL_WIDTH - 1),
		24731 => to_unsigned(22823, LUT_AMPL_WIDTH - 1),
		24732 => to_unsigned(22821, LUT_AMPL_WIDTH - 1),
		24733 => to_unsigned(22818, LUT_AMPL_WIDTH - 1),
		24734 => to_unsigned(22816, LUT_AMPL_WIDTH - 1),
		24735 => to_unsigned(22814, LUT_AMPL_WIDTH - 1),
		24736 => to_unsigned(22812, LUT_AMPL_WIDTH - 1),
		24737 => to_unsigned(22809, LUT_AMPL_WIDTH - 1),
		24738 => to_unsigned(22807, LUT_AMPL_WIDTH - 1),
		24739 => to_unsigned(22805, LUT_AMPL_WIDTH - 1),
		24740 => to_unsigned(22803, LUT_AMPL_WIDTH - 1),
		24741 => to_unsigned(22800, LUT_AMPL_WIDTH - 1),
		24742 => to_unsigned(22798, LUT_AMPL_WIDTH - 1),
		24743 => to_unsigned(22796, LUT_AMPL_WIDTH - 1),
		24744 => to_unsigned(22794, LUT_AMPL_WIDTH - 1),
		24745 => to_unsigned(22791, LUT_AMPL_WIDTH - 1),
		24746 => to_unsigned(22789, LUT_AMPL_WIDTH - 1),
		24747 => to_unsigned(22787, LUT_AMPL_WIDTH - 1),
		24748 => to_unsigned(22785, LUT_AMPL_WIDTH - 1),
		24749 => to_unsigned(22782, LUT_AMPL_WIDTH - 1),
		24750 => to_unsigned(22780, LUT_AMPL_WIDTH - 1),
		24751 => to_unsigned(22778, LUT_AMPL_WIDTH - 1),
		24752 => to_unsigned(22776, LUT_AMPL_WIDTH - 1),
		24753 => to_unsigned(22773, LUT_AMPL_WIDTH - 1),
		24754 => to_unsigned(22771, LUT_AMPL_WIDTH - 1),
		24755 => to_unsigned(22769, LUT_AMPL_WIDTH - 1),
		24756 => to_unsigned(22766, LUT_AMPL_WIDTH - 1),
		24757 => to_unsigned(22764, LUT_AMPL_WIDTH - 1),
		24758 => to_unsigned(22762, LUT_AMPL_WIDTH - 1),
		24759 => to_unsigned(22760, LUT_AMPL_WIDTH - 1),
		24760 => to_unsigned(22757, LUT_AMPL_WIDTH - 1),
		24761 => to_unsigned(22755, LUT_AMPL_WIDTH - 1),
		24762 => to_unsigned(22753, LUT_AMPL_WIDTH - 1),
		24763 => to_unsigned(22751, LUT_AMPL_WIDTH - 1),
		24764 => to_unsigned(22748, LUT_AMPL_WIDTH - 1),
		24765 => to_unsigned(22746, LUT_AMPL_WIDTH - 1),
		24766 => to_unsigned(22744, LUT_AMPL_WIDTH - 1),
		24767 => to_unsigned(22742, LUT_AMPL_WIDTH - 1),
		24768 => to_unsigned(22739, LUT_AMPL_WIDTH - 1),
		24769 => to_unsigned(22737, LUT_AMPL_WIDTH - 1),
		24770 => to_unsigned(22735, LUT_AMPL_WIDTH - 1),
		24771 => to_unsigned(22733, LUT_AMPL_WIDTH - 1),
		24772 => to_unsigned(22730, LUT_AMPL_WIDTH - 1),
		24773 => to_unsigned(22728, LUT_AMPL_WIDTH - 1),
		24774 => to_unsigned(22726, LUT_AMPL_WIDTH - 1),
		24775 => to_unsigned(22724, LUT_AMPL_WIDTH - 1),
		24776 => to_unsigned(22721, LUT_AMPL_WIDTH - 1),
		24777 => to_unsigned(22719, LUT_AMPL_WIDTH - 1),
		24778 => to_unsigned(22717, LUT_AMPL_WIDTH - 1),
		24779 => to_unsigned(22714, LUT_AMPL_WIDTH - 1),
		24780 => to_unsigned(22712, LUT_AMPL_WIDTH - 1),
		24781 => to_unsigned(22710, LUT_AMPL_WIDTH - 1),
		24782 => to_unsigned(22708, LUT_AMPL_WIDTH - 1),
		24783 => to_unsigned(22705, LUT_AMPL_WIDTH - 1),
		24784 => to_unsigned(22703, LUT_AMPL_WIDTH - 1),
		24785 => to_unsigned(22701, LUT_AMPL_WIDTH - 1),
		24786 => to_unsigned(22699, LUT_AMPL_WIDTH - 1),
		24787 => to_unsigned(22696, LUT_AMPL_WIDTH - 1),
		24788 => to_unsigned(22694, LUT_AMPL_WIDTH - 1),
		24789 => to_unsigned(22692, LUT_AMPL_WIDTH - 1),
		24790 => to_unsigned(22690, LUT_AMPL_WIDTH - 1),
		24791 => to_unsigned(22687, LUT_AMPL_WIDTH - 1),
		24792 => to_unsigned(22685, LUT_AMPL_WIDTH - 1),
		24793 => to_unsigned(22683, LUT_AMPL_WIDTH - 1),
		24794 => to_unsigned(22680, LUT_AMPL_WIDTH - 1),
		24795 => to_unsigned(22678, LUT_AMPL_WIDTH - 1),
		24796 => to_unsigned(22676, LUT_AMPL_WIDTH - 1),
		24797 => to_unsigned(22674, LUT_AMPL_WIDTH - 1),
		24798 => to_unsigned(22671, LUT_AMPL_WIDTH - 1),
		24799 => to_unsigned(22669, LUT_AMPL_WIDTH - 1),
		24800 => to_unsigned(22667, LUT_AMPL_WIDTH - 1),
		24801 => to_unsigned(22665, LUT_AMPL_WIDTH - 1),
		24802 => to_unsigned(22662, LUT_AMPL_WIDTH - 1),
		24803 => to_unsigned(22660, LUT_AMPL_WIDTH - 1),
		24804 => to_unsigned(22658, LUT_AMPL_WIDTH - 1),
		24805 => to_unsigned(22656, LUT_AMPL_WIDTH - 1),
		24806 => to_unsigned(22653, LUT_AMPL_WIDTH - 1),
		24807 => to_unsigned(22651, LUT_AMPL_WIDTH - 1),
		24808 => to_unsigned(22649, LUT_AMPL_WIDTH - 1),
		24809 => to_unsigned(22646, LUT_AMPL_WIDTH - 1),
		24810 => to_unsigned(22644, LUT_AMPL_WIDTH - 1),
		24811 => to_unsigned(22642, LUT_AMPL_WIDTH - 1),
		24812 => to_unsigned(22640, LUT_AMPL_WIDTH - 1),
		24813 => to_unsigned(22637, LUT_AMPL_WIDTH - 1),
		24814 => to_unsigned(22635, LUT_AMPL_WIDTH - 1),
		24815 => to_unsigned(22633, LUT_AMPL_WIDTH - 1),
		24816 => to_unsigned(22631, LUT_AMPL_WIDTH - 1),
		24817 => to_unsigned(22628, LUT_AMPL_WIDTH - 1),
		24818 => to_unsigned(22626, LUT_AMPL_WIDTH - 1),
		24819 => to_unsigned(22624, LUT_AMPL_WIDTH - 1),
		24820 => to_unsigned(22621, LUT_AMPL_WIDTH - 1),
		24821 => to_unsigned(22619, LUT_AMPL_WIDTH - 1),
		24822 => to_unsigned(22617, LUT_AMPL_WIDTH - 1),
		24823 => to_unsigned(22615, LUT_AMPL_WIDTH - 1),
		24824 => to_unsigned(22612, LUT_AMPL_WIDTH - 1),
		24825 => to_unsigned(22610, LUT_AMPL_WIDTH - 1),
		24826 => to_unsigned(22608, LUT_AMPL_WIDTH - 1),
		24827 => to_unsigned(22606, LUT_AMPL_WIDTH - 1),
		24828 => to_unsigned(22603, LUT_AMPL_WIDTH - 1),
		24829 => to_unsigned(22601, LUT_AMPL_WIDTH - 1),
		24830 => to_unsigned(22599, LUT_AMPL_WIDTH - 1),
		24831 => to_unsigned(22596, LUT_AMPL_WIDTH - 1),
		24832 => to_unsigned(22594, LUT_AMPL_WIDTH - 1),
		24833 => to_unsigned(22592, LUT_AMPL_WIDTH - 1),
		24834 => to_unsigned(22590, LUT_AMPL_WIDTH - 1),
		24835 => to_unsigned(22587, LUT_AMPL_WIDTH - 1),
		24836 => to_unsigned(22585, LUT_AMPL_WIDTH - 1),
		24837 => to_unsigned(22583, LUT_AMPL_WIDTH - 1),
		24838 => to_unsigned(22581, LUT_AMPL_WIDTH - 1),
		24839 => to_unsigned(22578, LUT_AMPL_WIDTH - 1),
		24840 => to_unsigned(22576, LUT_AMPL_WIDTH - 1),
		24841 => to_unsigned(22574, LUT_AMPL_WIDTH - 1),
		24842 => to_unsigned(22571, LUT_AMPL_WIDTH - 1),
		24843 => to_unsigned(22569, LUT_AMPL_WIDTH - 1),
		24844 => to_unsigned(22567, LUT_AMPL_WIDTH - 1),
		24845 => to_unsigned(22565, LUT_AMPL_WIDTH - 1),
		24846 => to_unsigned(22562, LUT_AMPL_WIDTH - 1),
		24847 => to_unsigned(22560, LUT_AMPL_WIDTH - 1),
		24848 => to_unsigned(22558, LUT_AMPL_WIDTH - 1),
		24849 => to_unsigned(22555, LUT_AMPL_WIDTH - 1),
		24850 => to_unsigned(22553, LUT_AMPL_WIDTH - 1),
		24851 => to_unsigned(22551, LUT_AMPL_WIDTH - 1),
		24852 => to_unsigned(22549, LUT_AMPL_WIDTH - 1),
		24853 => to_unsigned(22546, LUT_AMPL_WIDTH - 1),
		24854 => to_unsigned(22544, LUT_AMPL_WIDTH - 1),
		24855 => to_unsigned(22542, LUT_AMPL_WIDTH - 1),
		24856 => to_unsigned(22540, LUT_AMPL_WIDTH - 1),
		24857 => to_unsigned(22537, LUT_AMPL_WIDTH - 1),
		24858 => to_unsigned(22535, LUT_AMPL_WIDTH - 1),
		24859 => to_unsigned(22533, LUT_AMPL_WIDTH - 1),
		24860 => to_unsigned(22530, LUT_AMPL_WIDTH - 1),
		24861 => to_unsigned(22528, LUT_AMPL_WIDTH - 1),
		24862 => to_unsigned(22526, LUT_AMPL_WIDTH - 1),
		24863 => to_unsigned(22524, LUT_AMPL_WIDTH - 1),
		24864 => to_unsigned(22521, LUT_AMPL_WIDTH - 1),
		24865 => to_unsigned(22519, LUT_AMPL_WIDTH - 1),
		24866 => to_unsigned(22517, LUT_AMPL_WIDTH - 1),
		24867 => to_unsigned(22514, LUT_AMPL_WIDTH - 1),
		24868 => to_unsigned(22512, LUT_AMPL_WIDTH - 1),
		24869 => to_unsigned(22510, LUT_AMPL_WIDTH - 1),
		24870 => to_unsigned(22508, LUT_AMPL_WIDTH - 1),
		24871 => to_unsigned(22505, LUT_AMPL_WIDTH - 1),
		24872 => to_unsigned(22503, LUT_AMPL_WIDTH - 1),
		24873 => to_unsigned(22501, LUT_AMPL_WIDTH - 1),
		24874 => to_unsigned(22498, LUT_AMPL_WIDTH - 1),
		24875 => to_unsigned(22496, LUT_AMPL_WIDTH - 1),
		24876 => to_unsigned(22494, LUT_AMPL_WIDTH - 1),
		24877 => to_unsigned(22492, LUT_AMPL_WIDTH - 1),
		24878 => to_unsigned(22489, LUT_AMPL_WIDTH - 1),
		24879 => to_unsigned(22487, LUT_AMPL_WIDTH - 1),
		24880 => to_unsigned(22485, LUT_AMPL_WIDTH - 1),
		24881 => to_unsigned(22482, LUT_AMPL_WIDTH - 1),
		24882 => to_unsigned(22480, LUT_AMPL_WIDTH - 1),
		24883 => to_unsigned(22478, LUT_AMPL_WIDTH - 1),
		24884 => to_unsigned(22476, LUT_AMPL_WIDTH - 1),
		24885 => to_unsigned(22473, LUT_AMPL_WIDTH - 1),
		24886 => to_unsigned(22471, LUT_AMPL_WIDTH - 1),
		24887 => to_unsigned(22469, LUT_AMPL_WIDTH - 1),
		24888 => to_unsigned(22466, LUT_AMPL_WIDTH - 1),
		24889 => to_unsigned(22464, LUT_AMPL_WIDTH - 1),
		24890 => to_unsigned(22462, LUT_AMPL_WIDTH - 1),
		24891 => to_unsigned(22460, LUT_AMPL_WIDTH - 1),
		24892 => to_unsigned(22457, LUT_AMPL_WIDTH - 1),
		24893 => to_unsigned(22455, LUT_AMPL_WIDTH - 1),
		24894 => to_unsigned(22453, LUT_AMPL_WIDTH - 1),
		24895 => to_unsigned(22450, LUT_AMPL_WIDTH - 1),
		24896 => to_unsigned(22448, LUT_AMPL_WIDTH - 1),
		24897 => to_unsigned(22446, LUT_AMPL_WIDTH - 1),
		24898 => to_unsigned(22444, LUT_AMPL_WIDTH - 1),
		24899 => to_unsigned(22441, LUT_AMPL_WIDTH - 1),
		24900 => to_unsigned(22439, LUT_AMPL_WIDTH - 1),
		24901 => to_unsigned(22437, LUT_AMPL_WIDTH - 1),
		24902 => to_unsigned(22434, LUT_AMPL_WIDTH - 1),
		24903 => to_unsigned(22432, LUT_AMPL_WIDTH - 1),
		24904 => to_unsigned(22430, LUT_AMPL_WIDTH - 1),
		24905 => to_unsigned(22428, LUT_AMPL_WIDTH - 1),
		24906 => to_unsigned(22425, LUT_AMPL_WIDTH - 1),
		24907 => to_unsigned(22423, LUT_AMPL_WIDTH - 1),
		24908 => to_unsigned(22421, LUT_AMPL_WIDTH - 1),
		24909 => to_unsigned(22418, LUT_AMPL_WIDTH - 1),
		24910 => to_unsigned(22416, LUT_AMPL_WIDTH - 1),
		24911 => to_unsigned(22414, LUT_AMPL_WIDTH - 1),
		24912 => to_unsigned(22411, LUT_AMPL_WIDTH - 1),
		24913 => to_unsigned(22409, LUT_AMPL_WIDTH - 1),
		24914 => to_unsigned(22407, LUT_AMPL_WIDTH - 1),
		24915 => to_unsigned(22405, LUT_AMPL_WIDTH - 1),
		24916 => to_unsigned(22402, LUT_AMPL_WIDTH - 1),
		24917 => to_unsigned(22400, LUT_AMPL_WIDTH - 1),
		24918 => to_unsigned(22398, LUT_AMPL_WIDTH - 1),
		24919 => to_unsigned(22395, LUT_AMPL_WIDTH - 1),
		24920 => to_unsigned(22393, LUT_AMPL_WIDTH - 1),
		24921 => to_unsigned(22391, LUT_AMPL_WIDTH - 1),
		24922 => to_unsigned(22389, LUT_AMPL_WIDTH - 1),
		24923 => to_unsigned(22386, LUT_AMPL_WIDTH - 1),
		24924 => to_unsigned(22384, LUT_AMPL_WIDTH - 1),
		24925 => to_unsigned(22382, LUT_AMPL_WIDTH - 1),
		24926 => to_unsigned(22379, LUT_AMPL_WIDTH - 1),
		24927 => to_unsigned(22377, LUT_AMPL_WIDTH - 1),
		24928 => to_unsigned(22375, LUT_AMPL_WIDTH - 1),
		24929 => to_unsigned(22373, LUT_AMPL_WIDTH - 1),
		24930 => to_unsigned(22370, LUT_AMPL_WIDTH - 1),
		24931 => to_unsigned(22368, LUT_AMPL_WIDTH - 1),
		24932 => to_unsigned(22366, LUT_AMPL_WIDTH - 1),
		24933 => to_unsigned(22363, LUT_AMPL_WIDTH - 1),
		24934 => to_unsigned(22361, LUT_AMPL_WIDTH - 1),
		24935 => to_unsigned(22359, LUT_AMPL_WIDTH - 1),
		24936 => to_unsigned(22356, LUT_AMPL_WIDTH - 1),
		24937 => to_unsigned(22354, LUT_AMPL_WIDTH - 1),
		24938 => to_unsigned(22352, LUT_AMPL_WIDTH - 1),
		24939 => to_unsigned(22350, LUT_AMPL_WIDTH - 1),
		24940 => to_unsigned(22347, LUT_AMPL_WIDTH - 1),
		24941 => to_unsigned(22345, LUT_AMPL_WIDTH - 1),
		24942 => to_unsigned(22343, LUT_AMPL_WIDTH - 1),
		24943 => to_unsigned(22340, LUT_AMPL_WIDTH - 1),
		24944 => to_unsigned(22338, LUT_AMPL_WIDTH - 1),
		24945 => to_unsigned(22336, LUT_AMPL_WIDTH - 1),
		24946 => to_unsigned(22333, LUT_AMPL_WIDTH - 1),
		24947 => to_unsigned(22331, LUT_AMPL_WIDTH - 1),
		24948 => to_unsigned(22329, LUT_AMPL_WIDTH - 1),
		24949 => to_unsigned(22327, LUT_AMPL_WIDTH - 1),
		24950 => to_unsigned(22324, LUT_AMPL_WIDTH - 1),
		24951 => to_unsigned(22322, LUT_AMPL_WIDTH - 1),
		24952 => to_unsigned(22320, LUT_AMPL_WIDTH - 1),
		24953 => to_unsigned(22317, LUT_AMPL_WIDTH - 1),
		24954 => to_unsigned(22315, LUT_AMPL_WIDTH - 1),
		24955 => to_unsigned(22313, LUT_AMPL_WIDTH - 1),
		24956 => to_unsigned(22310, LUT_AMPL_WIDTH - 1),
		24957 => to_unsigned(22308, LUT_AMPL_WIDTH - 1),
		24958 => to_unsigned(22306, LUT_AMPL_WIDTH - 1),
		24959 => to_unsigned(22304, LUT_AMPL_WIDTH - 1),
		24960 => to_unsigned(22301, LUT_AMPL_WIDTH - 1),
		24961 => to_unsigned(22299, LUT_AMPL_WIDTH - 1),
		24962 => to_unsigned(22297, LUT_AMPL_WIDTH - 1),
		24963 => to_unsigned(22294, LUT_AMPL_WIDTH - 1),
		24964 => to_unsigned(22292, LUT_AMPL_WIDTH - 1),
		24965 => to_unsigned(22290, LUT_AMPL_WIDTH - 1),
		24966 => to_unsigned(22287, LUT_AMPL_WIDTH - 1),
		24967 => to_unsigned(22285, LUT_AMPL_WIDTH - 1),
		24968 => to_unsigned(22283, LUT_AMPL_WIDTH - 1),
		24969 => to_unsigned(22281, LUT_AMPL_WIDTH - 1),
		24970 => to_unsigned(22278, LUT_AMPL_WIDTH - 1),
		24971 => to_unsigned(22276, LUT_AMPL_WIDTH - 1),
		24972 => to_unsigned(22274, LUT_AMPL_WIDTH - 1),
		24973 => to_unsigned(22271, LUT_AMPL_WIDTH - 1),
		24974 => to_unsigned(22269, LUT_AMPL_WIDTH - 1),
		24975 => to_unsigned(22267, LUT_AMPL_WIDTH - 1),
		24976 => to_unsigned(22264, LUT_AMPL_WIDTH - 1),
		24977 => to_unsigned(22262, LUT_AMPL_WIDTH - 1),
		24978 => to_unsigned(22260, LUT_AMPL_WIDTH - 1),
		24979 => to_unsigned(22257, LUT_AMPL_WIDTH - 1),
		24980 => to_unsigned(22255, LUT_AMPL_WIDTH - 1),
		24981 => to_unsigned(22253, LUT_AMPL_WIDTH - 1),
		24982 => to_unsigned(22251, LUT_AMPL_WIDTH - 1),
		24983 => to_unsigned(22248, LUT_AMPL_WIDTH - 1),
		24984 => to_unsigned(22246, LUT_AMPL_WIDTH - 1),
		24985 => to_unsigned(22244, LUT_AMPL_WIDTH - 1),
		24986 => to_unsigned(22241, LUT_AMPL_WIDTH - 1),
		24987 => to_unsigned(22239, LUT_AMPL_WIDTH - 1),
		24988 => to_unsigned(22237, LUT_AMPL_WIDTH - 1),
		24989 => to_unsigned(22234, LUT_AMPL_WIDTH - 1),
		24990 => to_unsigned(22232, LUT_AMPL_WIDTH - 1),
		24991 => to_unsigned(22230, LUT_AMPL_WIDTH - 1),
		24992 => to_unsigned(22227, LUT_AMPL_WIDTH - 1),
		24993 => to_unsigned(22225, LUT_AMPL_WIDTH - 1),
		24994 => to_unsigned(22223, LUT_AMPL_WIDTH - 1),
		24995 => to_unsigned(22221, LUT_AMPL_WIDTH - 1),
		24996 => to_unsigned(22218, LUT_AMPL_WIDTH - 1),
		24997 => to_unsigned(22216, LUT_AMPL_WIDTH - 1),
		24998 => to_unsigned(22214, LUT_AMPL_WIDTH - 1),
		24999 => to_unsigned(22211, LUT_AMPL_WIDTH - 1),
		25000 => to_unsigned(22209, LUT_AMPL_WIDTH - 1),
		25001 => to_unsigned(22207, LUT_AMPL_WIDTH - 1),
		25002 => to_unsigned(22204, LUT_AMPL_WIDTH - 1),
		25003 => to_unsigned(22202, LUT_AMPL_WIDTH - 1),
		25004 => to_unsigned(22200, LUT_AMPL_WIDTH - 1),
		25005 => to_unsigned(22197, LUT_AMPL_WIDTH - 1),
		25006 => to_unsigned(22195, LUT_AMPL_WIDTH - 1),
		25007 => to_unsigned(22193, LUT_AMPL_WIDTH - 1),
		25008 => to_unsigned(22191, LUT_AMPL_WIDTH - 1),
		25009 => to_unsigned(22188, LUT_AMPL_WIDTH - 1),
		25010 => to_unsigned(22186, LUT_AMPL_WIDTH - 1),
		25011 => to_unsigned(22184, LUT_AMPL_WIDTH - 1),
		25012 => to_unsigned(22181, LUT_AMPL_WIDTH - 1),
		25013 => to_unsigned(22179, LUT_AMPL_WIDTH - 1),
		25014 => to_unsigned(22177, LUT_AMPL_WIDTH - 1),
		25015 => to_unsigned(22174, LUT_AMPL_WIDTH - 1),
		25016 => to_unsigned(22172, LUT_AMPL_WIDTH - 1),
		25017 => to_unsigned(22170, LUT_AMPL_WIDTH - 1),
		25018 => to_unsigned(22167, LUT_AMPL_WIDTH - 1),
		25019 => to_unsigned(22165, LUT_AMPL_WIDTH - 1),
		25020 => to_unsigned(22163, LUT_AMPL_WIDTH - 1),
		25021 => to_unsigned(22160, LUT_AMPL_WIDTH - 1),
		25022 => to_unsigned(22158, LUT_AMPL_WIDTH - 1),
		25023 => to_unsigned(22156, LUT_AMPL_WIDTH - 1),
		25024 => to_unsigned(22154, LUT_AMPL_WIDTH - 1),
		25025 => to_unsigned(22151, LUT_AMPL_WIDTH - 1),
		25026 => to_unsigned(22149, LUT_AMPL_WIDTH - 1),
		25027 => to_unsigned(22147, LUT_AMPL_WIDTH - 1),
		25028 => to_unsigned(22144, LUT_AMPL_WIDTH - 1),
		25029 => to_unsigned(22142, LUT_AMPL_WIDTH - 1),
		25030 => to_unsigned(22140, LUT_AMPL_WIDTH - 1),
		25031 => to_unsigned(22137, LUT_AMPL_WIDTH - 1),
		25032 => to_unsigned(22135, LUT_AMPL_WIDTH - 1),
		25033 => to_unsigned(22133, LUT_AMPL_WIDTH - 1),
		25034 => to_unsigned(22130, LUT_AMPL_WIDTH - 1),
		25035 => to_unsigned(22128, LUT_AMPL_WIDTH - 1),
		25036 => to_unsigned(22126, LUT_AMPL_WIDTH - 1),
		25037 => to_unsigned(22123, LUT_AMPL_WIDTH - 1),
		25038 => to_unsigned(22121, LUT_AMPL_WIDTH - 1),
		25039 => to_unsigned(22119, LUT_AMPL_WIDTH - 1),
		25040 => to_unsigned(22116, LUT_AMPL_WIDTH - 1),
		25041 => to_unsigned(22114, LUT_AMPL_WIDTH - 1),
		25042 => to_unsigned(22112, LUT_AMPL_WIDTH - 1),
		25043 => to_unsigned(22110, LUT_AMPL_WIDTH - 1),
		25044 => to_unsigned(22107, LUT_AMPL_WIDTH - 1),
		25045 => to_unsigned(22105, LUT_AMPL_WIDTH - 1),
		25046 => to_unsigned(22103, LUT_AMPL_WIDTH - 1),
		25047 => to_unsigned(22100, LUT_AMPL_WIDTH - 1),
		25048 => to_unsigned(22098, LUT_AMPL_WIDTH - 1),
		25049 => to_unsigned(22096, LUT_AMPL_WIDTH - 1),
		25050 => to_unsigned(22093, LUT_AMPL_WIDTH - 1),
		25051 => to_unsigned(22091, LUT_AMPL_WIDTH - 1),
		25052 => to_unsigned(22089, LUT_AMPL_WIDTH - 1),
		25053 => to_unsigned(22086, LUT_AMPL_WIDTH - 1),
		25054 => to_unsigned(22084, LUT_AMPL_WIDTH - 1),
		25055 => to_unsigned(22082, LUT_AMPL_WIDTH - 1),
		25056 => to_unsigned(22079, LUT_AMPL_WIDTH - 1),
		25057 => to_unsigned(22077, LUT_AMPL_WIDTH - 1),
		25058 => to_unsigned(22075, LUT_AMPL_WIDTH - 1),
		25059 => to_unsigned(22072, LUT_AMPL_WIDTH - 1),
		25060 => to_unsigned(22070, LUT_AMPL_WIDTH - 1),
		25061 => to_unsigned(22068, LUT_AMPL_WIDTH - 1),
		25062 => to_unsigned(22065, LUT_AMPL_WIDTH - 1),
		25063 => to_unsigned(22063, LUT_AMPL_WIDTH - 1),
		25064 => to_unsigned(22061, LUT_AMPL_WIDTH - 1),
		25065 => to_unsigned(22058, LUT_AMPL_WIDTH - 1),
		25066 => to_unsigned(22056, LUT_AMPL_WIDTH - 1),
		25067 => to_unsigned(22054, LUT_AMPL_WIDTH - 1),
		25068 => to_unsigned(22051, LUT_AMPL_WIDTH - 1),
		25069 => to_unsigned(22049, LUT_AMPL_WIDTH - 1),
		25070 => to_unsigned(22047, LUT_AMPL_WIDTH - 1),
		25071 => to_unsigned(22045, LUT_AMPL_WIDTH - 1),
		25072 => to_unsigned(22042, LUT_AMPL_WIDTH - 1),
		25073 => to_unsigned(22040, LUT_AMPL_WIDTH - 1),
		25074 => to_unsigned(22038, LUT_AMPL_WIDTH - 1),
		25075 => to_unsigned(22035, LUT_AMPL_WIDTH - 1),
		25076 => to_unsigned(22033, LUT_AMPL_WIDTH - 1),
		25077 => to_unsigned(22031, LUT_AMPL_WIDTH - 1),
		25078 => to_unsigned(22028, LUT_AMPL_WIDTH - 1),
		25079 => to_unsigned(22026, LUT_AMPL_WIDTH - 1),
		25080 => to_unsigned(22024, LUT_AMPL_WIDTH - 1),
		25081 => to_unsigned(22021, LUT_AMPL_WIDTH - 1),
		25082 => to_unsigned(22019, LUT_AMPL_WIDTH - 1),
		25083 => to_unsigned(22017, LUT_AMPL_WIDTH - 1),
		25084 => to_unsigned(22014, LUT_AMPL_WIDTH - 1),
		25085 => to_unsigned(22012, LUT_AMPL_WIDTH - 1),
		25086 => to_unsigned(22010, LUT_AMPL_WIDTH - 1),
		25087 => to_unsigned(22007, LUT_AMPL_WIDTH - 1),
		25088 => to_unsigned(22005, LUT_AMPL_WIDTH - 1),
		25089 => to_unsigned(22003, LUT_AMPL_WIDTH - 1),
		25090 => to_unsigned(22000, LUT_AMPL_WIDTH - 1),
		25091 => to_unsigned(21998, LUT_AMPL_WIDTH - 1),
		25092 => to_unsigned(21996, LUT_AMPL_WIDTH - 1),
		25093 => to_unsigned(21993, LUT_AMPL_WIDTH - 1),
		25094 => to_unsigned(21991, LUT_AMPL_WIDTH - 1),
		25095 => to_unsigned(21989, LUT_AMPL_WIDTH - 1),
		25096 => to_unsigned(21986, LUT_AMPL_WIDTH - 1),
		25097 => to_unsigned(21984, LUT_AMPL_WIDTH - 1),
		25098 => to_unsigned(21982, LUT_AMPL_WIDTH - 1),
		25099 => to_unsigned(21979, LUT_AMPL_WIDTH - 1),
		25100 => to_unsigned(21977, LUT_AMPL_WIDTH - 1),
		25101 => to_unsigned(21975, LUT_AMPL_WIDTH - 1),
		25102 => to_unsigned(21972, LUT_AMPL_WIDTH - 1),
		25103 => to_unsigned(21970, LUT_AMPL_WIDTH - 1),
		25104 => to_unsigned(21968, LUT_AMPL_WIDTH - 1),
		25105 => to_unsigned(21965, LUT_AMPL_WIDTH - 1),
		25106 => to_unsigned(21963, LUT_AMPL_WIDTH - 1),
		25107 => to_unsigned(21961, LUT_AMPL_WIDTH - 1),
		25108 => to_unsigned(21958, LUT_AMPL_WIDTH - 1),
		25109 => to_unsigned(21956, LUT_AMPL_WIDTH - 1),
		25110 => to_unsigned(21954, LUT_AMPL_WIDTH - 1),
		25111 => to_unsigned(21951, LUT_AMPL_WIDTH - 1),
		25112 => to_unsigned(21949, LUT_AMPL_WIDTH - 1),
		25113 => to_unsigned(21947, LUT_AMPL_WIDTH - 1),
		25114 => to_unsigned(21944, LUT_AMPL_WIDTH - 1),
		25115 => to_unsigned(21942, LUT_AMPL_WIDTH - 1),
		25116 => to_unsigned(21940, LUT_AMPL_WIDTH - 1),
		25117 => to_unsigned(21937, LUT_AMPL_WIDTH - 1),
		25118 => to_unsigned(21935, LUT_AMPL_WIDTH - 1),
		25119 => to_unsigned(21933, LUT_AMPL_WIDTH - 1),
		25120 => to_unsigned(21930, LUT_AMPL_WIDTH - 1),
		25121 => to_unsigned(21928, LUT_AMPL_WIDTH - 1),
		25122 => to_unsigned(21926, LUT_AMPL_WIDTH - 1),
		25123 => to_unsigned(21923, LUT_AMPL_WIDTH - 1),
		25124 => to_unsigned(21921, LUT_AMPL_WIDTH - 1),
		25125 => to_unsigned(21919, LUT_AMPL_WIDTH - 1),
		25126 => to_unsigned(21916, LUT_AMPL_WIDTH - 1),
		25127 => to_unsigned(21914, LUT_AMPL_WIDTH - 1),
		25128 => to_unsigned(21912, LUT_AMPL_WIDTH - 1),
		25129 => to_unsigned(21909, LUT_AMPL_WIDTH - 1),
		25130 => to_unsigned(21907, LUT_AMPL_WIDTH - 1),
		25131 => to_unsigned(21905, LUT_AMPL_WIDTH - 1),
		25132 => to_unsigned(21902, LUT_AMPL_WIDTH - 1),
		25133 => to_unsigned(21900, LUT_AMPL_WIDTH - 1),
		25134 => to_unsigned(21898, LUT_AMPL_WIDTH - 1),
		25135 => to_unsigned(21895, LUT_AMPL_WIDTH - 1),
		25136 => to_unsigned(21893, LUT_AMPL_WIDTH - 1),
		25137 => to_unsigned(21891, LUT_AMPL_WIDTH - 1),
		25138 => to_unsigned(21888, LUT_AMPL_WIDTH - 1),
		25139 => to_unsigned(21886, LUT_AMPL_WIDTH - 1),
		25140 => to_unsigned(21884, LUT_AMPL_WIDTH - 1),
		25141 => to_unsigned(21881, LUT_AMPL_WIDTH - 1),
		25142 => to_unsigned(21879, LUT_AMPL_WIDTH - 1),
		25143 => to_unsigned(21877, LUT_AMPL_WIDTH - 1),
		25144 => to_unsigned(21874, LUT_AMPL_WIDTH - 1),
		25145 => to_unsigned(21872, LUT_AMPL_WIDTH - 1),
		25146 => to_unsigned(21870, LUT_AMPL_WIDTH - 1),
		25147 => to_unsigned(21867, LUT_AMPL_WIDTH - 1),
		25148 => to_unsigned(21865, LUT_AMPL_WIDTH - 1),
		25149 => to_unsigned(21863, LUT_AMPL_WIDTH - 1),
		25150 => to_unsigned(21860, LUT_AMPL_WIDTH - 1),
		25151 => to_unsigned(21858, LUT_AMPL_WIDTH - 1),
		25152 => to_unsigned(21856, LUT_AMPL_WIDTH - 1),
		25153 => to_unsigned(21853, LUT_AMPL_WIDTH - 1),
		25154 => to_unsigned(21851, LUT_AMPL_WIDTH - 1),
		25155 => to_unsigned(21849, LUT_AMPL_WIDTH - 1),
		25156 => to_unsigned(21846, LUT_AMPL_WIDTH - 1),
		25157 => to_unsigned(21844, LUT_AMPL_WIDTH - 1),
		25158 => to_unsigned(21842, LUT_AMPL_WIDTH - 1),
		25159 => to_unsigned(21839, LUT_AMPL_WIDTH - 1),
		25160 => to_unsigned(21837, LUT_AMPL_WIDTH - 1),
		25161 => to_unsigned(21835, LUT_AMPL_WIDTH - 1),
		25162 => to_unsigned(21832, LUT_AMPL_WIDTH - 1),
		25163 => to_unsigned(21830, LUT_AMPL_WIDTH - 1),
		25164 => to_unsigned(21827, LUT_AMPL_WIDTH - 1),
		25165 => to_unsigned(21825, LUT_AMPL_WIDTH - 1),
		25166 => to_unsigned(21823, LUT_AMPL_WIDTH - 1),
		25167 => to_unsigned(21820, LUT_AMPL_WIDTH - 1),
		25168 => to_unsigned(21818, LUT_AMPL_WIDTH - 1),
		25169 => to_unsigned(21816, LUT_AMPL_WIDTH - 1),
		25170 => to_unsigned(21813, LUT_AMPL_WIDTH - 1),
		25171 => to_unsigned(21811, LUT_AMPL_WIDTH - 1),
		25172 => to_unsigned(21809, LUT_AMPL_WIDTH - 1),
		25173 => to_unsigned(21806, LUT_AMPL_WIDTH - 1),
		25174 => to_unsigned(21804, LUT_AMPL_WIDTH - 1),
		25175 => to_unsigned(21802, LUT_AMPL_WIDTH - 1),
		25176 => to_unsigned(21799, LUT_AMPL_WIDTH - 1),
		25177 => to_unsigned(21797, LUT_AMPL_WIDTH - 1),
		25178 => to_unsigned(21795, LUT_AMPL_WIDTH - 1),
		25179 => to_unsigned(21792, LUT_AMPL_WIDTH - 1),
		25180 => to_unsigned(21790, LUT_AMPL_WIDTH - 1),
		25181 => to_unsigned(21788, LUT_AMPL_WIDTH - 1),
		25182 => to_unsigned(21785, LUT_AMPL_WIDTH - 1),
		25183 => to_unsigned(21783, LUT_AMPL_WIDTH - 1),
		25184 => to_unsigned(21781, LUT_AMPL_WIDTH - 1),
		25185 => to_unsigned(21778, LUT_AMPL_WIDTH - 1),
		25186 => to_unsigned(21776, LUT_AMPL_WIDTH - 1),
		25187 => to_unsigned(21774, LUT_AMPL_WIDTH - 1),
		25188 => to_unsigned(21771, LUT_AMPL_WIDTH - 1),
		25189 => to_unsigned(21769, LUT_AMPL_WIDTH - 1),
		25190 => to_unsigned(21766, LUT_AMPL_WIDTH - 1),
		25191 => to_unsigned(21764, LUT_AMPL_WIDTH - 1),
		25192 => to_unsigned(21762, LUT_AMPL_WIDTH - 1),
		25193 => to_unsigned(21759, LUT_AMPL_WIDTH - 1),
		25194 => to_unsigned(21757, LUT_AMPL_WIDTH - 1),
		25195 => to_unsigned(21755, LUT_AMPL_WIDTH - 1),
		25196 => to_unsigned(21752, LUT_AMPL_WIDTH - 1),
		25197 => to_unsigned(21750, LUT_AMPL_WIDTH - 1),
		25198 => to_unsigned(21748, LUT_AMPL_WIDTH - 1),
		25199 => to_unsigned(21745, LUT_AMPL_WIDTH - 1),
		25200 => to_unsigned(21743, LUT_AMPL_WIDTH - 1),
		25201 => to_unsigned(21741, LUT_AMPL_WIDTH - 1),
		25202 => to_unsigned(21738, LUT_AMPL_WIDTH - 1),
		25203 => to_unsigned(21736, LUT_AMPL_WIDTH - 1),
		25204 => to_unsigned(21734, LUT_AMPL_WIDTH - 1),
		25205 => to_unsigned(21731, LUT_AMPL_WIDTH - 1),
		25206 => to_unsigned(21729, LUT_AMPL_WIDTH - 1),
		25207 => to_unsigned(21727, LUT_AMPL_WIDTH - 1),
		25208 => to_unsigned(21724, LUT_AMPL_WIDTH - 1),
		25209 => to_unsigned(21722, LUT_AMPL_WIDTH - 1),
		25210 => to_unsigned(21719, LUT_AMPL_WIDTH - 1),
		25211 => to_unsigned(21717, LUT_AMPL_WIDTH - 1),
		25212 => to_unsigned(21715, LUT_AMPL_WIDTH - 1),
		25213 => to_unsigned(21712, LUT_AMPL_WIDTH - 1),
		25214 => to_unsigned(21710, LUT_AMPL_WIDTH - 1),
		25215 => to_unsigned(21708, LUT_AMPL_WIDTH - 1),
		25216 => to_unsigned(21705, LUT_AMPL_WIDTH - 1),
		25217 => to_unsigned(21703, LUT_AMPL_WIDTH - 1),
		25218 => to_unsigned(21701, LUT_AMPL_WIDTH - 1),
		25219 => to_unsigned(21698, LUT_AMPL_WIDTH - 1),
		25220 => to_unsigned(21696, LUT_AMPL_WIDTH - 1),
		25221 => to_unsigned(21694, LUT_AMPL_WIDTH - 1),
		25222 => to_unsigned(21691, LUT_AMPL_WIDTH - 1),
		25223 => to_unsigned(21689, LUT_AMPL_WIDTH - 1),
		25224 => to_unsigned(21687, LUT_AMPL_WIDTH - 1),
		25225 => to_unsigned(21684, LUT_AMPL_WIDTH - 1),
		25226 => to_unsigned(21682, LUT_AMPL_WIDTH - 1),
		25227 => to_unsigned(21679, LUT_AMPL_WIDTH - 1),
		25228 => to_unsigned(21677, LUT_AMPL_WIDTH - 1),
		25229 => to_unsigned(21675, LUT_AMPL_WIDTH - 1),
		25230 => to_unsigned(21672, LUT_AMPL_WIDTH - 1),
		25231 => to_unsigned(21670, LUT_AMPL_WIDTH - 1),
		25232 => to_unsigned(21668, LUT_AMPL_WIDTH - 1),
		25233 => to_unsigned(21665, LUT_AMPL_WIDTH - 1),
		25234 => to_unsigned(21663, LUT_AMPL_WIDTH - 1),
		25235 => to_unsigned(21661, LUT_AMPL_WIDTH - 1),
		25236 => to_unsigned(21658, LUT_AMPL_WIDTH - 1),
		25237 => to_unsigned(21656, LUT_AMPL_WIDTH - 1),
		25238 => to_unsigned(21654, LUT_AMPL_WIDTH - 1),
		25239 => to_unsigned(21651, LUT_AMPL_WIDTH - 1),
		25240 => to_unsigned(21649, LUT_AMPL_WIDTH - 1),
		25241 => to_unsigned(21646, LUT_AMPL_WIDTH - 1),
		25242 => to_unsigned(21644, LUT_AMPL_WIDTH - 1),
		25243 => to_unsigned(21642, LUT_AMPL_WIDTH - 1),
		25244 => to_unsigned(21639, LUT_AMPL_WIDTH - 1),
		25245 => to_unsigned(21637, LUT_AMPL_WIDTH - 1),
		25246 => to_unsigned(21635, LUT_AMPL_WIDTH - 1),
		25247 => to_unsigned(21632, LUT_AMPL_WIDTH - 1),
		25248 => to_unsigned(21630, LUT_AMPL_WIDTH - 1),
		25249 => to_unsigned(21628, LUT_AMPL_WIDTH - 1),
		25250 => to_unsigned(21625, LUT_AMPL_WIDTH - 1),
		25251 => to_unsigned(21623, LUT_AMPL_WIDTH - 1),
		25252 => to_unsigned(21621, LUT_AMPL_WIDTH - 1),
		25253 => to_unsigned(21618, LUT_AMPL_WIDTH - 1),
		25254 => to_unsigned(21616, LUT_AMPL_WIDTH - 1),
		25255 => to_unsigned(21613, LUT_AMPL_WIDTH - 1),
		25256 => to_unsigned(21611, LUT_AMPL_WIDTH - 1),
		25257 => to_unsigned(21609, LUT_AMPL_WIDTH - 1),
		25258 => to_unsigned(21606, LUT_AMPL_WIDTH - 1),
		25259 => to_unsigned(21604, LUT_AMPL_WIDTH - 1),
		25260 => to_unsigned(21602, LUT_AMPL_WIDTH - 1),
		25261 => to_unsigned(21599, LUT_AMPL_WIDTH - 1),
		25262 => to_unsigned(21597, LUT_AMPL_WIDTH - 1),
		25263 => to_unsigned(21595, LUT_AMPL_WIDTH - 1),
		25264 => to_unsigned(21592, LUT_AMPL_WIDTH - 1),
		25265 => to_unsigned(21590, LUT_AMPL_WIDTH - 1),
		25266 => to_unsigned(21587, LUT_AMPL_WIDTH - 1),
		25267 => to_unsigned(21585, LUT_AMPL_WIDTH - 1),
		25268 => to_unsigned(21583, LUT_AMPL_WIDTH - 1),
		25269 => to_unsigned(21580, LUT_AMPL_WIDTH - 1),
		25270 => to_unsigned(21578, LUT_AMPL_WIDTH - 1),
		25271 => to_unsigned(21576, LUT_AMPL_WIDTH - 1),
		25272 => to_unsigned(21573, LUT_AMPL_WIDTH - 1),
		25273 => to_unsigned(21571, LUT_AMPL_WIDTH - 1),
		25274 => to_unsigned(21569, LUT_AMPL_WIDTH - 1),
		25275 => to_unsigned(21566, LUT_AMPL_WIDTH - 1),
		25276 => to_unsigned(21564, LUT_AMPL_WIDTH - 1),
		25277 => to_unsigned(21561, LUT_AMPL_WIDTH - 1),
		25278 => to_unsigned(21559, LUT_AMPL_WIDTH - 1),
		25279 => to_unsigned(21557, LUT_AMPL_WIDTH - 1),
		25280 => to_unsigned(21554, LUT_AMPL_WIDTH - 1),
		25281 => to_unsigned(21552, LUT_AMPL_WIDTH - 1),
		25282 => to_unsigned(21550, LUT_AMPL_WIDTH - 1),
		25283 => to_unsigned(21547, LUT_AMPL_WIDTH - 1),
		25284 => to_unsigned(21545, LUT_AMPL_WIDTH - 1),
		25285 => to_unsigned(21543, LUT_AMPL_WIDTH - 1),
		25286 => to_unsigned(21540, LUT_AMPL_WIDTH - 1),
		25287 => to_unsigned(21538, LUT_AMPL_WIDTH - 1),
		25288 => to_unsigned(21535, LUT_AMPL_WIDTH - 1),
		25289 => to_unsigned(21533, LUT_AMPL_WIDTH - 1),
		25290 => to_unsigned(21531, LUT_AMPL_WIDTH - 1),
		25291 => to_unsigned(21528, LUT_AMPL_WIDTH - 1),
		25292 => to_unsigned(21526, LUT_AMPL_WIDTH - 1),
		25293 => to_unsigned(21524, LUT_AMPL_WIDTH - 1),
		25294 => to_unsigned(21521, LUT_AMPL_WIDTH - 1),
		25295 => to_unsigned(21519, LUT_AMPL_WIDTH - 1),
		25296 => to_unsigned(21516, LUT_AMPL_WIDTH - 1),
		25297 => to_unsigned(21514, LUT_AMPL_WIDTH - 1),
		25298 => to_unsigned(21512, LUT_AMPL_WIDTH - 1),
		25299 => to_unsigned(21509, LUT_AMPL_WIDTH - 1),
		25300 => to_unsigned(21507, LUT_AMPL_WIDTH - 1),
		25301 => to_unsigned(21505, LUT_AMPL_WIDTH - 1),
		25302 => to_unsigned(21502, LUT_AMPL_WIDTH - 1),
		25303 => to_unsigned(21500, LUT_AMPL_WIDTH - 1),
		25304 => to_unsigned(21498, LUT_AMPL_WIDTH - 1),
		25305 => to_unsigned(21495, LUT_AMPL_WIDTH - 1),
		25306 => to_unsigned(21493, LUT_AMPL_WIDTH - 1),
		25307 => to_unsigned(21490, LUT_AMPL_WIDTH - 1),
		25308 => to_unsigned(21488, LUT_AMPL_WIDTH - 1),
		25309 => to_unsigned(21486, LUT_AMPL_WIDTH - 1),
		25310 => to_unsigned(21483, LUT_AMPL_WIDTH - 1),
		25311 => to_unsigned(21481, LUT_AMPL_WIDTH - 1),
		25312 => to_unsigned(21479, LUT_AMPL_WIDTH - 1),
		25313 => to_unsigned(21476, LUT_AMPL_WIDTH - 1),
		25314 => to_unsigned(21474, LUT_AMPL_WIDTH - 1),
		25315 => to_unsigned(21471, LUT_AMPL_WIDTH - 1),
		25316 => to_unsigned(21469, LUT_AMPL_WIDTH - 1),
		25317 => to_unsigned(21467, LUT_AMPL_WIDTH - 1),
		25318 => to_unsigned(21464, LUT_AMPL_WIDTH - 1),
		25319 => to_unsigned(21462, LUT_AMPL_WIDTH - 1),
		25320 => to_unsigned(21460, LUT_AMPL_WIDTH - 1),
		25321 => to_unsigned(21457, LUT_AMPL_WIDTH - 1),
		25322 => to_unsigned(21455, LUT_AMPL_WIDTH - 1),
		25323 => to_unsigned(21452, LUT_AMPL_WIDTH - 1),
		25324 => to_unsigned(21450, LUT_AMPL_WIDTH - 1),
		25325 => to_unsigned(21448, LUT_AMPL_WIDTH - 1),
		25326 => to_unsigned(21445, LUT_AMPL_WIDTH - 1),
		25327 => to_unsigned(21443, LUT_AMPL_WIDTH - 1),
		25328 => to_unsigned(21441, LUT_AMPL_WIDTH - 1),
		25329 => to_unsigned(21438, LUT_AMPL_WIDTH - 1),
		25330 => to_unsigned(21436, LUT_AMPL_WIDTH - 1),
		25331 => to_unsigned(21433, LUT_AMPL_WIDTH - 1),
		25332 => to_unsigned(21431, LUT_AMPL_WIDTH - 1),
		25333 => to_unsigned(21429, LUT_AMPL_WIDTH - 1),
		25334 => to_unsigned(21426, LUT_AMPL_WIDTH - 1),
		25335 => to_unsigned(21424, LUT_AMPL_WIDTH - 1),
		25336 => to_unsigned(21422, LUT_AMPL_WIDTH - 1),
		25337 => to_unsigned(21419, LUT_AMPL_WIDTH - 1),
		25338 => to_unsigned(21417, LUT_AMPL_WIDTH - 1),
		25339 => to_unsigned(21414, LUT_AMPL_WIDTH - 1),
		25340 => to_unsigned(21412, LUT_AMPL_WIDTH - 1),
		25341 => to_unsigned(21410, LUT_AMPL_WIDTH - 1),
		25342 => to_unsigned(21407, LUT_AMPL_WIDTH - 1),
		25343 => to_unsigned(21405, LUT_AMPL_WIDTH - 1),
		25344 => to_unsigned(21403, LUT_AMPL_WIDTH - 1),
		25345 => to_unsigned(21400, LUT_AMPL_WIDTH - 1),
		25346 => to_unsigned(21398, LUT_AMPL_WIDTH - 1),
		25347 => to_unsigned(21395, LUT_AMPL_WIDTH - 1),
		25348 => to_unsigned(21393, LUT_AMPL_WIDTH - 1),
		25349 => to_unsigned(21391, LUT_AMPL_WIDTH - 1),
		25350 => to_unsigned(21388, LUT_AMPL_WIDTH - 1),
		25351 => to_unsigned(21386, LUT_AMPL_WIDTH - 1),
		25352 => to_unsigned(21383, LUT_AMPL_WIDTH - 1),
		25353 => to_unsigned(21381, LUT_AMPL_WIDTH - 1),
		25354 => to_unsigned(21379, LUT_AMPL_WIDTH - 1),
		25355 => to_unsigned(21376, LUT_AMPL_WIDTH - 1),
		25356 => to_unsigned(21374, LUT_AMPL_WIDTH - 1),
		25357 => to_unsigned(21372, LUT_AMPL_WIDTH - 1),
		25358 => to_unsigned(21369, LUT_AMPL_WIDTH - 1),
		25359 => to_unsigned(21367, LUT_AMPL_WIDTH - 1),
		25360 => to_unsigned(21364, LUT_AMPL_WIDTH - 1),
		25361 => to_unsigned(21362, LUT_AMPL_WIDTH - 1),
		25362 => to_unsigned(21360, LUT_AMPL_WIDTH - 1),
		25363 => to_unsigned(21357, LUT_AMPL_WIDTH - 1),
		25364 => to_unsigned(21355, LUT_AMPL_WIDTH - 1),
		25365 => to_unsigned(21353, LUT_AMPL_WIDTH - 1),
		25366 => to_unsigned(21350, LUT_AMPL_WIDTH - 1),
		25367 => to_unsigned(21348, LUT_AMPL_WIDTH - 1),
		25368 => to_unsigned(21345, LUT_AMPL_WIDTH - 1),
		25369 => to_unsigned(21343, LUT_AMPL_WIDTH - 1),
		25370 => to_unsigned(21341, LUT_AMPL_WIDTH - 1),
		25371 => to_unsigned(21338, LUT_AMPL_WIDTH - 1),
		25372 => to_unsigned(21336, LUT_AMPL_WIDTH - 1),
		25373 => to_unsigned(21333, LUT_AMPL_WIDTH - 1),
		25374 => to_unsigned(21331, LUT_AMPL_WIDTH - 1),
		25375 => to_unsigned(21329, LUT_AMPL_WIDTH - 1),
		25376 => to_unsigned(21326, LUT_AMPL_WIDTH - 1),
		25377 => to_unsigned(21324, LUT_AMPL_WIDTH - 1),
		25378 => to_unsigned(21322, LUT_AMPL_WIDTH - 1),
		25379 => to_unsigned(21319, LUT_AMPL_WIDTH - 1),
		25380 => to_unsigned(21317, LUT_AMPL_WIDTH - 1),
		25381 => to_unsigned(21314, LUT_AMPL_WIDTH - 1),
		25382 => to_unsigned(21312, LUT_AMPL_WIDTH - 1),
		25383 => to_unsigned(21310, LUT_AMPL_WIDTH - 1),
		25384 => to_unsigned(21307, LUT_AMPL_WIDTH - 1),
		25385 => to_unsigned(21305, LUT_AMPL_WIDTH - 1),
		25386 => to_unsigned(21302, LUT_AMPL_WIDTH - 1),
		25387 => to_unsigned(21300, LUT_AMPL_WIDTH - 1),
		25388 => to_unsigned(21298, LUT_AMPL_WIDTH - 1),
		25389 => to_unsigned(21295, LUT_AMPL_WIDTH - 1),
		25390 => to_unsigned(21293, LUT_AMPL_WIDTH - 1),
		25391 => to_unsigned(21290, LUT_AMPL_WIDTH - 1),
		25392 => to_unsigned(21288, LUT_AMPL_WIDTH - 1),
		25393 => to_unsigned(21286, LUT_AMPL_WIDTH - 1),
		25394 => to_unsigned(21283, LUT_AMPL_WIDTH - 1),
		25395 => to_unsigned(21281, LUT_AMPL_WIDTH - 1),
		25396 => to_unsigned(21279, LUT_AMPL_WIDTH - 1),
		25397 => to_unsigned(21276, LUT_AMPL_WIDTH - 1),
		25398 => to_unsigned(21274, LUT_AMPL_WIDTH - 1),
		25399 => to_unsigned(21271, LUT_AMPL_WIDTH - 1),
		25400 => to_unsigned(21269, LUT_AMPL_WIDTH - 1),
		25401 => to_unsigned(21267, LUT_AMPL_WIDTH - 1),
		25402 => to_unsigned(21264, LUT_AMPL_WIDTH - 1),
		25403 => to_unsigned(21262, LUT_AMPL_WIDTH - 1),
		25404 => to_unsigned(21259, LUT_AMPL_WIDTH - 1),
		25405 => to_unsigned(21257, LUT_AMPL_WIDTH - 1),
		25406 => to_unsigned(21255, LUT_AMPL_WIDTH - 1),
		25407 => to_unsigned(21252, LUT_AMPL_WIDTH - 1),
		25408 => to_unsigned(21250, LUT_AMPL_WIDTH - 1),
		25409 => to_unsigned(21247, LUT_AMPL_WIDTH - 1),
		25410 => to_unsigned(21245, LUT_AMPL_WIDTH - 1),
		25411 => to_unsigned(21243, LUT_AMPL_WIDTH - 1),
		25412 => to_unsigned(21240, LUT_AMPL_WIDTH - 1),
		25413 => to_unsigned(21238, LUT_AMPL_WIDTH - 1),
		25414 => to_unsigned(21236, LUT_AMPL_WIDTH - 1),
		25415 => to_unsigned(21233, LUT_AMPL_WIDTH - 1),
		25416 => to_unsigned(21231, LUT_AMPL_WIDTH - 1),
		25417 => to_unsigned(21228, LUT_AMPL_WIDTH - 1),
		25418 => to_unsigned(21226, LUT_AMPL_WIDTH - 1),
		25419 => to_unsigned(21224, LUT_AMPL_WIDTH - 1),
		25420 => to_unsigned(21221, LUT_AMPL_WIDTH - 1),
		25421 => to_unsigned(21219, LUT_AMPL_WIDTH - 1),
		25422 => to_unsigned(21216, LUT_AMPL_WIDTH - 1),
		25423 => to_unsigned(21214, LUT_AMPL_WIDTH - 1),
		25424 => to_unsigned(21212, LUT_AMPL_WIDTH - 1),
		25425 => to_unsigned(21209, LUT_AMPL_WIDTH - 1),
		25426 => to_unsigned(21207, LUT_AMPL_WIDTH - 1),
		25427 => to_unsigned(21204, LUT_AMPL_WIDTH - 1),
		25428 => to_unsigned(21202, LUT_AMPL_WIDTH - 1),
		25429 => to_unsigned(21200, LUT_AMPL_WIDTH - 1),
		25430 => to_unsigned(21197, LUT_AMPL_WIDTH - 1),
		25431 => to_unsigned(21195, LUT_AMPL_WIDTH - 1),
		25432 => to_unsigned(21192, LUT_AMPL_WIDTH - 1),
		25433 => to_unsigned(21190, LUT_AMPL_WIDTH - 1),
		25434 => to_unsigned(21188, LUT_AMPL_WIDTH - 1),
		25435 => to_unsigned(21185, LUT_AMPL_WIDTH - 1),
		25436 => to_unsigned(21183, LUT_AMPL_WIDTH - 1),
		25437 => to_unsigned(21180, LUT_AMPL_WIDTH - 1),
		25438 => to_unsigned(21178, LUT_AMPL_WIDTH - 1),
		25439 => to_unsigned(21176, LUT_AMPL_WIDTH - 1),
		25440 => to_unsigned(21173, LUT_AMPL_WIDTH - 1),
		25441 => to_unsigned(21171, LUT_AMPL_WIDTH - 1),
		25442 => to_unsigned(21168, LUT_AMPL_WIDTH - 1),
		25443 => to_unsigned(21166, LUT_AMPL_WIDTH - 1),
		25444 => to_unsigned(21164, LUT_AMPL_WIDTH - 1),
		25445 => to_unsigned(21161, LUT_AMPL_WIDTH - 1),
		25446 => to_unsigned(21159, LUT_AMPL_WIDTH - 1),
		25447 => to_unsigned(21156, LUT_AMPL_WIDTH - 1),
		25448 => to_unsigned(21154, LUT_AMPL_WIDTH - 1),
		25449 => to_unsigned(21152, LUT_AMPL_WIDTH - 1),
		25450 => to_unsigned(21149, LUT_AMPL_WIDTH - 1),
		25451 => to_unsigned(21147, LUT_AMPL_WIDTH - 1),
		25452 => to_unsigned(21144, LUT_AMPL_WIDTH - 1),
		25453 => to_unsigned(21142, LUT_AMPL_WIDTH - 1),
		25454 => to_unsigned(21140, LUT_AMPL_WIDTH - 1),
		25455 => to_unsigned(21137, LUT_AMPL_WIDTH - 1),
		25456 => to_unsigned(21135, LUT_AMPL_WIDTH - 1),
		25457 => to_unsigned(21132, LUT_AMPL_WIDTH - 1),
		25458 => to_unsigned(21130, LUT_AMPL_WIDTH - 1),
		25459 => to_unsigned(21128, LUT_AMPL_WIDTH - 1),
		25460 => to_unsigned(21125, LUT_AMPL_WIDTH - 1),
		25461 => to_unsigned(21123, LUT_AMPL_WIDTH - 1),
		25462 => to_unsigned(21120, LUT_AMPL_WIDTH - 1),
		25463 => to_unsigned(21118, LUT_AMPL_WIDTH - 1),
		25464 => to_unsigned(21116, LUT_AMPL_WIDTH - 1),
		25465 => to_unsigned(21113, LUT_AMPL_WIDTH - 1),
		25466 => to_unsigned(21111, LUT_AMPL_WIDTH - 1),
		25467 => to_unsigned(21108, LUT_AMPL_WIDTH - 1),
		25468 => to_unsigned(21106, LUT_AMPL_WIDTH - 1),
		25469 => to_unsigned(21104, LUT_AMPL_WIDTH - 1),
		25470 => to_unsigned(21101, LUT_AMPL_WIDTH - 1),
		25471 => to_unsigned(21099, LUT_AMPL_WIDTH - 1),
		25472 => to_unsigned(21096, LUT_AMPL_WIDTH - 1),
		25473 => to_unsigned(21094, LUT_AMPL_WIDTH - 1),
		25474 => to_unsigned(21092, LUT_AMPL_WIDTH - 1),
		25475 => to_unsigned(21089, LUT_AMPL_WIDTH - 1),
		25476 => to_unsigned(21087, LUT_AMPL_WIDTH - 1),
		25477 => to_unsigned(21084, LUT_AMPL_WIDTH - 1),
		25478 => to_unsigned(21082, LUT_AMPL_WIDTH - 1),
		25479 => to_unsigned(21080, LUT_AMPL_WIDTH - 1),
		25480 => to_unsigned(21077, LUT_AMPL_WIDTH - 1),
		25481 => to_unsigned(21075, LUT_AMPL_WIDTH - 1),
		25482 => to_unsigned(21072, LUT_AMPL_WIDTH - 1),
		25483 => to_unsigned(21070, LUT_AMPL_WIDTH - 1),
		25484 => to_unsigned(21068, LUT_AMPL_WIDTH - 1),
		25485 => to_unsigned(21065, LUT_AMPL_WIDTH - 1),
		25486 => to_unsigned(21063, LUT_AMPL_WIDTH - 1),
		25487 => to_unsigned(21060, LUT_AMPL_WIDTH - 1),
		25488 => to_unsigned(21058, LUT_AMPL_WIDTH - 1),
		25489 => to_unsigned(21056, LUT_AMPL_WIDTH - 1),
		25490 => to_unsigned(21053, LUT_AMPL_WIDTH - 1),
		25491 => to_unsigned(21051, LUT_AMPL_WIDTH - 1),
		25492 => to_unsigned(21048, LUT_AMPL_WIDTH - 1),
		25493 => to_unsigned(21046, LUT_AMPL_WIDTH - 1),
		25494 => to_unsigned(21043, LUT_AMPL_WIDTH - 1),
		25495 => to_unsigned(21041, LUT_AMPL_WIDTH - 1),
		25496 => to_unsigned(21039, LUT_AMPL_WIDTH - 1),
		25497 => to_unsigned(21036, LUT_AMPL_WIDTH - 1),
		25498 => to_unsigned(21034, LUT_AMPL_WIDTH - 1),
		25499 => to_unsigned(21031, LUT_AMPL_WIDTH - 1),
		25500 => to_unsigned(21029, LUT_AMPL_WIDTH - 1),
		25501 => to_unsigned(21027, LUT_AMPL_WIDTH - 1),
		25502 => to_unsigned(21024, LUT_AMPL_WIDTH - 1),
		25503 => to_unsigned(21022, LUT_AMPL_WIDTH - 1),
		25504 => to_unsigned(21019, LUT_AMPL_WIDTH - 1),
		25505 => to_unsigned(21017, LUT_AMPL_WIDTH - 1),
		25506 => to_unsigned(21015, LUT_AMPL_WIDTH - 1),
		25507 => to_unsigned(21012, LUT_AMPL_WIDTH - 1),
		25508 => to_unsigned(21010, LUT_AMPL_WIDTH - 1),
		25509 => to_unsigned(21007, LUT_AMPL_WIDTH - 1),
		25510 => to_unsigned(21005, LUT_AMPL_WIDTH - 1),
		25511 => to_unsigned(21003, LUT_AMPL_WIDTH - 1),
		25512 => to_unsigned(21000, LUT_AMPL_WIDTH - 1),
		25513 => to_unsigned(20998, LUT_AMPL_WIDTH - 1),
		25514 => to_unsigned(20995, LUT_AMPL_WIDTH - 1),
		25515 => to_unsigned(20993, LUT_AMPL_WIDTH - 1),
		25516 => to_unsigned(20990, LUT_AMPL_WIDTH - 1),
		25517 => to_unsigned(20988, LUT_AMPL_WIDTH - 1),
		25518 => to_unsigned(20986, LUT_AMPL_WIDTH - 1),
		25519 => to_unsigned(20983, LUT_AMPL_WIDTH - 1),
		25520 => to_unsigned(20981, LUT_AMPL_WIDTH - 1),
		25521 => to_unsigned(20978, LUT_AMPL_WIDTH - 1),
		25522 => to_unsigned(20976, LUT_AMPL_WIDTH - 1),
		25523 => to_unsigned(20974, LUT_AMPL_WIDTH - 1),
		25524 => to_unsigned(20971, LUT_AMPL_WIDTH - 1),
		25525 => to_unsigned(20969, LUT_AMPL_WIDTH - 1),
		25526 => to_unsigned(20966, LUT_AMPL_WIDTH - 1),
		25527 => to_unsigned(20964, LUT_AMPL_WIDTH - 1),
		25528 => to_unsigned(20962, LUT_AMPL_WIDTH - 1),
		25529 => to_unsigned(20959, LUT_AMPL_WIDTH - 1),
		25530 => to_unsigned(20957, LUT_AMPL_WIDTH - 1),
		25531 => to_unsigned(20954, LUT_AMPL_WIDTH - 1),
		25532 => to_unsigned(20952, LUT_AMPL_WIDTH - 1),
		25533 => to_unsigned(20949, LUT_AMPL_WIDTH - 1),
		25534 => to_unsigned(20947, LUT_AMPL_WIDTH - 1),
		25535 => to_unsigned(20945, LUT_AMPL_WIDTH - 1),
		25536 => to_unsigned(20942, LUT_AMPL_WIDTH - 1),
		25537 => to_unsigned(20940, LUT_AMPL_WIDTH - 1),
		25538 => to_unsigned(20937, LUT_AMPL_WIDTH - 1),
		25539 => to_unsigned(20935, LUT_AMPL_WIDTH - 1),
		25540 => to_unsigned(20933, LUT_AMPL_WIDTH - 1),
		25541 => to_unsigned(20930, LUT_AMPL_WIDTH - 1),
		25542 => to_unsigned(20928, LUT_AMPL_WIDTH - 1),
		25543 => to_unsigned(20925, LUT_AMPL_WIDTH - 1),
		25544 => to_unsigned(20923, LUT_AMPL_WIDTH - 1),
		25545 => to_unsigned(20920, LUT_AMPL_WIDTH - 1),
		25546 => to_unsigned(20918, LUT_AMPL_WIDTH - 1),
		25547 => to_unsigned(20916, LUT_AMPL_WIDTH - 1),
		25548 => to_unsigned(20913, LUT_AMPL_WIDTH - 1),
		25549 => to_unsigned(20911, LUT_AMPL_WIDTH - 1),
		25550 => to_unsigned(20908, LUT_AMPL_WIDTH - 1),
		25551 => to_unsigned(20906, LUT_AMPL_WIDTH - 1),
		25552 => to_unsigned(20904, LUT_AMPL_WIDTH - 1),
		25553 => to_unsigned(20901, LUT_AMPL_WIDTH - 1),
		25554 => to_unsigned(20899, LUT_AMPL_WIDTH - 1),
		25555 => to_unsigned(20896, LUT_AMPL_WIDTH - 1),
		25556 => to_unsigned(20894, LUT_AMPL_WIDTH - 1),
		25557 => to_unsigned(20891, LUT_AMPL_WIDTH - 1),
		25558 => to_unsigned(20889, LUT_AMPL_WIDTH - 1),
		25559 => to_unsigned(20887, LUT_AMPL_WIDTH - 1),
		25560 => to_unsigned(20884, LUT_AMPL_WIDTH - 1),
		25561 => to_unsigned(20882, LUT_AMPL_WIDTH - 1),
		25562 => to_unsigned(20879, LUT_AMPL_WIDTH - 1),
		25563 => to_unsigned(20877, LUT_AMPL_WIDTH - 1),
		25564 => to_unsigned(20874, LUT_AMPL_WIDTH - 1),
		25565 => to_unsigned(20872, LUT_AMPL_WIDTH - 1),
		25566 => to_unsigned(20870, LUT_AMPL_WIDTH - 1),
		25567 => to_unsigned(20867, LUT_AMPL_WIDTH - 1),
		25568 => to_unsigned(20865, LUT_AMPL_WIDTH - 1),
		25569 => to_unsigned(20862, LUT_AMPL_WIDTH - 1),
		25570 => to_unsigned(20860, LUT_AMPL_WIDTH - 1),
		25571 => to_unsigned(20858, LUT_AMPL_WIDTH - 1),
		25572 => to_unsigned(20855, LUT_AMPL_WIDTH - 1),
		25573 => to_unsigned(20853, LUT_AMPL_WIDTH - 1),
		25574 => to_unsigned(20850, LUT_AMPL_WIDTH - 1),
		25575 => to_unsigned(20848, LUT_AMPL_WIDTH - 1),
		25576 => to_unsigned(20845, LUT_AMPL_WIDTH - 1),
		25577 => to_unsigned(20843, LUT_AMPL_WIDTH - 1),
		25578 => to_unsigned(20841, LUT_AMPL_WIDTH - 1),
		25579 => to_unsigned(20838, LUT_AMPL_WIDTH - 1),
		25580 => to_unsigned(20836, LUT_AMPL_WIDTH - 1),
		25581 => to_unsigned(20833, LUT_AMPL_WIDTH - 1),
		25582 => to_unsigned(20831, LUT_AMPL_WIDTH - 1),
		25583 => to_unsigned(20828, LUT_AMPL_WIDTH - 1),
		25584 => to_unsigned(20826, LUT_AMPL_WIDTH - 1),
		25585 => to_unsigned(20824, LUT_AMPL_WIDTH - 1),
		25586 => to_unsigned(20821, LUT_AMPL_WIDTH - 1),
		25587 => to_unsigned(20819, LUT_AMPL_WIDTH - 1),
		25588 => to_unsigned(20816, LUT_AMPL_WIDTH - 1),
		25589 => to_unsigned(20814, LUT_AMPL_WIDTH - 1),
		25590 => to_unsigned(20811, LUT_AMPL_WIDTH - 1),
		25591 => to_unsigned(20809, LUT_AMPL_WIDTH - 1),
		25592 => to_unsigned(20807, LUT_AMPL_WIDTH - 1),
		25593 => to_unsigned(20804, LUT_AMPL_WIDTH - 1),
		25594 => to_unsigned(20802, LUT_AMPL_WIDTH - 1),
		25595 => to_unsigned(20799, LUT_AMPL_WIDTH - 1),
		25596 => to_unsigned(20797, LUT_AMPL_WIDTH - 1),
		25597 => to_unsigned(20794, LUT_AMPL_WIDTH - 1),
		25598 => to_unsigned(20792, LUT_AMPL_WIDTH - 1),
		25599 => to_unsigned(20790, LUT_AMPL_WIDTH - 1),
		25600 => to_unsigned(20787, LUT_AMPL_WIDTH - 1),
		25601 => to_unsigned(20785, LUT_AMPL_WIDTH - 1),
		25602 => to_unsigned(20782, LUT_AMPL_WIDTH - 1),
		25603 => to_unsigned(20780, LUT_AMPL_WIDTH - 1),
		25604 => to_unsigned(20777, LUT_AMPL_WIDTH - 1),
		25605 => to_unsigned(20775, LUT_AMPL_WIDTH - 1),
		25606 => to_unsigned(20773, LUT_AMPL_WIDTH - 1),
		25607 => to_unsigned(20770, LUT_AMPL_WIDTH - 1),
		25608 => to_unsigned(20768, LUT_AMPL_WIDTH - 1),
		25609 => to_unsigned(20765, LUT_AMPL_WIDTH - 1),
		25610 => to_unsigned(20763, LUT_AMPL_WIDTH - 1),
		25611 => to_unsigned(20760, LUT_AMPL_WIDTH - 1),
		25612 => to_unsigned(20758, LUT_AMPL_WIDTH - 1),
		25613 => to_unsigned(20756, LUT_AMPL_WIDTH - 1),
		25614 => to_unsigned(20753, LUT_AMPL_WIDTH - 1),
		25615 => to_unsigned(20751, LUT_AMPL_WIDTH - 1),
		25616 => to_unsigned(20748, LUT_AMPL_WIDTH - 1),
		25617 => to_unsigned(20746, LUT_AMPL_WIDTH - 1),
		25618 => to_unsigned(20743, LUT_AMPL_WIDTH - 1),
		25619 => to_unsigned(20741, LUT_AMPL_WIDTH - 1),
		25620 => to_unsigned(20739, LUT_AMPL_WIDTH - 1),
		25621 => to_unsigned(20736, LUT_AMPL_WIDTH - 1),
		25622 => to_unsigned(20734, LUT_AMPL_WIDTH - 1),
		25623 => to_unsigned(20731, LUT_AMPL_WIDTH - 1),
		25624 => to_unsigned(20729, LUT_AMPL_WIDTH - 1),
		25625 => to_unsigned(20726, LUT_AMPL_WIDTH - 1),
		25626 => to_unsigned(20724, LUT_AMPL_WIDTH - 1),
		25627 => to_unsigned(20722, LUT_AMPL_WIDTH - 1),
		25628 => to_unsigned(20719, LUT_AMPL_WIDTH - 1),
		25629 => to_unsigned(20717, LUT_AMPL_WIDTH - 1),
		25630 => to_unsigned(20714, LUT_AMPL_WIDTH - 1),
		25631 => to_unsigned(20712, LUT_AMPL_WIDTH - 1),
		25632 => to_unsigned(20709, LUT_AMPL_WIDTH - 1),
		25633 => to_unsigned(20707, LUT_AMPL_WIDTH - 1),
		25634 => to_unsigned(20704, LUT_AMPL_WIDTH - 1),
		25635 => to_unsigned(20702, LUT_AMPL_WIDTH - 1),
		25636 => to_unsigned(20700, LUT_AMPL_WIDTH - 1),
		25637 => to_unsigned(20697, LUT_AMPL_WIDTH - 1),
		25638 => to_unsigned(20695, LUT_AMPL_WIDTH - 1),
		25639 => to_unsigned(20692, LUT_AMPL_WIDTH - 1),
		25640 => to_unsigned(20690, LUT_AMPL_WIDTH - 1),
		25641 => to_unsigned(20687, LUT_AMPL_WIDTH - 1),
		25642 => to_unsigned(20685, LUT_AMPL_WIDTH - 1),
		25643 => to_unsigned(20683, LUT_AMPL_WIDTH - 1),
		25644 => to_unsigned(20680, LUT_AMPL_WIDTH - 1),
		25645 => to_unsigned(20678, LUT_AMPL_WIDTH - 1),
		25646 => to_unsigned(20675, LUT_AMPL_WIDTH - 1),
		25647 => to_unsigned(20673, LUT_AMPL_WIDTH - 1),
		25648 => to_unsigned(20670, LUT_AMPL_WIDTH - 1),
		25649 => to_unsigned(20668, LUT_AMPL_WIDTH - 1),
		25650 => to_unsigned(20666, LUT_AMPL_WIDTH - 1),
		25651 => to_unsigned(20663, LUT_AMPL_WIDTH - 1),
		25652 => to_unsigned(20661, LUT_AMPL_WIDTH - 1),
		25653 => to_unsigned(20658, LUT_AMPL_WIDTH - 1),
		25654 => to_unsigned(20656, LUT_AMPL_WIDTH - 1),
		25655 => to_unsigned(20653, LUT_AMPL_WIDTH - 1),
		25656 => to_unsigned(20651, LUT_AMPL_WIDTH - 1),
		25657 => to_unsigned(20648, LUT_AMPL_WIDTH - 1),
		25658 => to_unsigned(20646, LUT_AMPL_WIDTH - 1),
		25659 => to_unsigned(20644, LUT_AMPL_WIDTH - 1),
		25660 => to_unsigned(20641, LUT_AMPL_WIDTH - 1),
		25661 => to_unsigned(20639, LUT_AMPL_WIDTH - 1),
		25662 => to_unsigned(20636, LUT_AMPL_WIDTH - 1),
		25663 => to_unsigned(20634, LUT_AMPL_WIDTH - 1),
		25664 => to_unsigned(20631, LUT_AMPL_WIDTH - 1),
		25665 => to_unsigned(20629, LUT_AMPL_WIDTH - 1),
		25666 => to_unsigned(20626, LUT_AMPL_WIDTH - 1),
		25667 => to_unsigned(20624, LUT_AMPL_WIDTH - 1),
		25668 => to_unsigned(20622, LUT_AMPL_WIDTH - 1),
		25669 => to_unsigned(20619, LUT_AMPL_WIDTH - 1),
		25670 => to_unsigned(20617, LUT_AMPL_WIDTH - 1),
		25671 => to_unsigned(20614, LUT_AMPL_WIDTH - 1),
		25672 => to_unsigned(20612, LUT_AMPL_WIDTH - 1),
		25673 => to_unsigned(20609, LUT_AMPL_WIDTH - 1),
		25674 => to_unsigned(20607, LUT_AMPL_WIDTH - 1),
		25675 => to_unsigned(20604, LUT_AMPL_WIDTH - 1),
		25676 => to_unsigned(20602, LUT_AMPL_WIDTH - 1),
		25677 => to_unsigned(20600, LUT_AMPL_WIDTH - 1),
		25678 => to_unsigned(20597, LUT_AMPL_WIDTH - 1),
		25679 => to_unsigned(20595, LUT_AMPL_WIDTH - 1),
		25680 => to_unsigned(20592, LUT_AMPL_WIDTH - 1),
		25681 => to_unsigned(20590, LUT_AMPL_WIDTH - 1),
		25682 => to_unsigned(20587, LUT_AMPL_WIDTH - 1),
		25683 => to_unsigned(20585, LUT_AMPL_WIDTH - 1),
		25684 => to_unsigned(20583, LUT_AMPL_WIDTH - 1),
		25685 => to_unsigned(20580, LUT_AMPL_WIDTH - 1),
		25686 => to_unsigned(20578, LUT_AMPL_WIDTH - 1),
		25687 => to_unsigned(20575, LUT_AMPL_WIDTH - 1),
		25688 => to_unsigned(20573, LUT_AMPL_WIDTH - 1),
		25689 => to_unsigned(20570, LUT_AMPL_WIDTH - 1),
		25690 => to_unsigned(20568, LUT_AMPL_WIDTH - 1),
		25691 => to_unsigned(20565, LUT_AMPL_WIDTH - 1),
		25692 => to_unsigned(20563, LUT_AMPL_WIDTH - 1),
		25693 => to_unsigned(20560, LUT_AMPL_WIDTH - 1),
		25694 => to_unsigned(20558, LUT_AMPL_WIDTH - 1),
		25695 => to_unsigned(20556, LUT_AMPL_WIDTH - 1),
		25696 => to_unsigned(20553, LUT_AMPL_WIDTH - 1),
		25697 => to_unsigned(20551, LUT_AMPL_WIDTH - 1),
		25698 => to_unsigned(20548, LUT_AMPL_WIDTH - 1),
		25699 => to_unsigned(20546, LUT_AMPL_WIDTH - 1),
		25700 => to_unsigned(20543, LUT_AMPL_WIDTH - 1),
		25701 => to_unsigned(20541, LUT_AMPL_WIDTH - 1),
		25702 => to_unsigned(20538, LUT_AMPL_WIDTH - 1),
		25703 => to_unsigned(20536, LUT_AMPL_WIDTH - 1),
		25704 => to_unsigned(20534, LUT_AMPL_WIDTH - 1),
		25705 => to_unsigned(20531, LUT_AMPL_WIDTH - 1),
		25706 => to_unsigned(20529, LUT_AMPL_WIDTH - 1),
		25707 => to_unsigned(20526, LUT_AMPL_WIDTH - 1),
		25708 => to_unsigned(20524, LUT_AMPL_WIDTH - 1),
		25709 => to_unsigned(20521, LUT_AMPL_WIDTH - 1),
		25710 => to_unsigned(20519, LUT_AMPL_WIDTH - 1),
		25711 => to_unsigned(20516, LUT_AMPL_WIDTH - 1),
		25712 => to_unsigned(20514, LUT_AMPL_WIDTH - 1),
		25713 => to_unsigned(20512, LUT_AMPL_WIDTH - 1),
		25714 => to_unsigned(20509, LUT_AMPL_WIDTH - 1),
		25715 => to_unsigned(20507, LUT_AMPL_WIDTH - 1),
		25716 => to_unsigned(20504, LUT_AMPL_WIDTH - 1),
		25717 => to_unsigned(20502, LUT_AMPL_WIDTH - 1),
		25718 => to_unsigned(20499, LUT_AMPL_WIDTH - 1),
		25719 => to_unsigned(20497, LUT_AMPL_WIDTH - 1),
		25720 => to_unsigned(20494, LUT_AMPL_WIDTH - 1),
		25721 => to_unsigned(20492, LUT_AMPL_WIDTH - 1),
		25722 => to_unsigned(20489, LUT_AMPL_WIDTH - 1),
		25723 => to_unsigned(20487, LUT_AMPL_WIDTH - 1),
		25724 => to_unsigned(20485, LUT_AMPL_WIDTH - 1),
		25725 => to_unsigned(20482, LUT_AMPL_WIDTH - 1),
		25726 => to_unsigned(20480, LUT_AMPL_WIDTH - 1),
		25727 => to_unsigned(20477, LUT_AMPL_WIDTH - 1),
		25728 => to_unsigned(20475, LUT_AMPL_WIDTH - 1),
		25729 => to_unsigned(20472, LUT_AMPL_WIDTH - 1),
		25730 => to_unsigned(20470, LUT_AMPL_WIDTH - 1),
		25731 => to_unsigned(20467, LUT_AMPL_WIDTH - 1),
		25732 => to_unsigned(20465, LUT_AMPL_WIDTH - 1),
		25733 => to_unsigned(20463, LUT_AMPL_WIDTH - 1),
		25734 => to_unsigned(20460, LUT_AMPL_WIDTH - 1),
		25735 => to_unsigned(20458, LUT_AMPL_WIDTH - 1),
		25736 => to_unsigned(20455, LUT_AMPL_WIDTH - 1),
		25737 => to_unsigned(20453, LUT_AMPL_WIDTH - 1),
		25738 => to_unsigned(20450, LUT_AMPL_WIDTH - 1),
		25739 => to_unsigned(20448, LUT_AMPL_WIDTH - 1),
		25740 => to_unsigned(20445, LUT_AMPL_WIDTH - 1),
		25741 => to_unsigned(20443, LUT_AMPL_WIDTH - 1),
		25742 => to_unsigned(20440, LUT_AMPL_WIDTH - 1),
		25743 => to_unsigned(20438, LUT_AMPL_WIDTH - 1),
		25744 => to_unsigned(20436, LUT_AMPL_WIDTH - 1),
		25745 => to_unsigned(20433, LUT_AMPL_WIDTH - 1),
		25746 => to_unsigned(20431, LUT_AMPL_WIDTH - 1),
		25747 => to_unsigned(20428, LUT_AMPL_WIDTH - 1),
		25748 => to_unsigned(20426, LUT_AMPL_WIDTH - 1),
		25749 => to_unsigned(20423, LUT_AMPL_WIDTH - 1),
		25750 => to_unsigned(20421, LUT_AMPL_WIDTH - 1),
		25751 => to_unsigned(20418, LUT_AMPL_WIDTH - 1),
		25752 => to_unsigned(20416, LUT_AMPL_WIDTH - 1),
		25753 => to_unsigned(20413, LUT_AMPL_WIDTH - 1),
		25754 => to_unsigned(20411, LUT_AMPL_WIDTH - 1),
		25755 => to_unsigned(20408, LUT_AMPL_WIDTH - 1),
		25756 => to_unsigned(20406, LUT_AMPL_WIDTH - 1),
		25757 => to_unsigned(20404, LUT_AMPL_WIDTH - 1),
		25758 => to_unsigned(20401, LUT_AMPL_WIDTH - 1),
		25759 => to_unsigned(20399, LUT_AMPL_WIDTH - 1),
		25760 => to_unsigned(20396, LUT_AMPL_WIDTH - 1),
		25761 => to_unsigned(20394, LUT_AMPL_WIDTH - 1),
		25762 => to_unsigned(20391, LUT_AMPL_WIDTH - 1),
		25763 => to_unsigned(20389, LUT_AMPL_WIDTH - 1),
		25764 => to_unsigned(20386, LUT_AMPL_WIDTH - 1),
		25765 => to_unsigned(20384, LUT_AMPL_WIDTH - 1),
		25766 => to_unsigned(20381, LUT_AMPL_WIDTH - 1),
		25767 => to_unsigned(20379, LUT_AMPL_WIDTH - 1),
		25768 => to_unsigned(20377, LUT_AMPL_WIDTH - 1),
		25769 => to_unsigned(20374, LUT_AMPL_WIDTH - 1),
		25770 => to_unsigned(20372, LUT_AMPL_WIDTH - 1),
		25771 => to_unsigned(20369, LUT_AMPL_WIDTH - 1),
		25772 => to_unsigned(20367, LUT_AMPL_WIDTH - 1),
		25773 => to_unsigned(20364, LUT_AMPL_WIDTH - 1),
		25774 => to_unsigned(20362, LUT_AMPL_WIDTH - 1),
		25775 => to_unsigned(20359, LUT_AMPL_WIDTH - 1),
		25776 => to_unsigned(20357, LUT_AMPL_WIDTH - 1),
		25777 => to_unsigned(20354, LUT_AMPL_WIDTH - 1),
		25778 => to_unsigned(20352, LUT_AMPL_WIDTH - 1),
		25779 => to_unsigned(20349, LUT_AMPL_WIDTH - 1),
		25780 => to_unsigned(20347, LUT_AMPL_WIDTH - 1),
		25781 => to_unsigned(20345, LUT_AMPL_WIDTH - 1),
		25782 => to_unsigned(20342, LUT_AMPL_WIDTH - 1),
		25783 => to_unsigned(20340, LUT_AMPL_WIDTH - 1),
		25784 => to_unsigned(20337, LUT_AMPL_WIDTH - 1),
		25785 => to_unsigned(20335, LUT_AMPL_WIDTH - 1),
		25786 => to_unsigned(20332, LUT_AMPL_WIDTH - 1),
		25787 => to_unsigned(20330, LUT_AMPL_WIDTH - 1),
		25788 => to_unsigned(20327, LUT_AMPL_WIDTH - 1),
		25789 => to_unsigned(20325, LUT_AMPL_WIDTH - 1),
		25790 => to_unsigned(20322, LUT_AMPL_WIDTH - 1),
		25791 => to_unsigned(20320, LUT_AMPL_WIDTH - 1),
		25792 => to_unsigned(20317, LUT_AMPL_WIDTH - 1),
		25793 => to_unsigned(20315, LUT_AMPL_WIDTH - 1),
		25794 => to_unsigned(20312, LUT_AMPL_WIDTH - 1),
		25795 => to_unsigned(20310, LUT_AMPL_WIDTH - 1),
		25796 => to_unsigned(20308, LUT_AMPL_WIDTH - 1),
		25797 => to_unsigned(20305, LUT_AMPL_WIDTH - 1),
		25798 => to_unsigned(20303, LUT_AMPL_WIDTH - 1),
		25799 => to_unsigned(20300, LUT_AMPL_WIDTH - 1),
		25800 => to_unsigned(20298, LUT_AMPL_WIDTH - 1),
		25801 => to_unsigned(20295, LUT_AMPL_WIDTH - 1),
		25802 => to_unsigned(20293, LUT_AMPL_WIDTH - 1),
		25803 => to_unsigned(20290, LUT_AMPL_WIDTH - 1),
		25804 => to_unsigned(20288, LUT_AMPL_WIDTH - 1),
		25805 => to_unsigned(20285, LUT_AMPL_WIDTH - 1),
		25806 => to_unsigned(20283, LUT_AMPL_WIDTH - 1),
		25807 => to_unsigned(20280, LUT_AMPL_WIDTH - 1),
		25808 => to_unsigned(20278, LUT_AMPL_WIDTH - 1),
		25809 => to_unsigned(20275, LUT_AMPL_WIDTH - 1),
		25810 => to_unsigned(20273, LUT_AMPL_WIDTH - 1),
		25811 => to_unsigned(20271, LUT_AMPL_WIDTH - 1),
		25812 => to_unsigned(20268, LUT_AMPL_WIDTH - 1),
		25813 => to_unsigned(20266, LUT_AMPL_WIDTH - 1),
		25814 => to_unsigned(20263, LUT_AMPL_WIDTH - 1),
		25815 => to_unsigned(20261, LUT_AMPL_WIDTH - 1),
		25816 => to_unsigned(20258, LUT_AMPL_WIDTH - 1),
		25817 => to_unsigned(20256, LUT_AMPL_WIDTH - 1),
		25818 => to_unsigned(20253, LUT_AMPL_WIDTH - 1),
		25819 => to_unsigned(20251, LUT_AMPL_WIDTH - 1),
		25820 => to_unsigned(20248, LUT_AMPL_WIDTH - 1),
		25821 => to_unsigned(20246, LUT_AMPL_WIDTH - 1),
		25822 => to_unsigned(20243, LUT_AMPL_WIDTH - 1),
		25823 => to_unsigned(20241, LUT_AMPL_WIDTH - 1),
		25824 => to_unsigned(20238, LUT_AMPL_WIDTH - 1),
		25825 => to_unsigned(20236, LUT_AMPL_WIDTH - 1),
		25826 => to_unsigned(20234, LUT_AMPL_WIDTH - 1),
		25827 => to_unsigned(20231, LUT_AMPL_WIDTH - 1),
		25828 => to_unsigned(20229, LUT_AMPL_WIDTH - 1),
		25829 => to_unsigned(20226, LUT_AMPL_WIDTH - 1),
		25830 => to_unsigned(20224, LUT_AMPL_WIDTH - 1),
		25831 => to_unsigned(20221, LUT_AMPL_WIDTH - 1),
		25832 => to_unsigned(20219, LUT_AMPL_WIDTH - 1),
		25833 => to_unsigned(20216, LUT_AMPL_WIDTH - 1),
		25834 => to_unsigned(20214, LUT_AMPL_WIDTH - 1),
		25835 => to_unsigned(20211, LUT_AMPL_WIDTH - 1),
		25836 => to_unsigned(20209, LUT_AMPL_WIDTH - 1),
		25837 => to_unsigned(20206, LUT_AMPL_WIDTH - 1),
		25838 => to_unsigned(20204, LUT_AMPL_WIDTH - 1),
		25839 => to_unsigned(20201, LUT_AMPL_WIDTH - 1),
		25840 => to_unsigned(20199, LUT_AMPL_WIDTH - 1),
		25841 => to_unsigned(20196, LUT_AMPL_WIDTH - 1),
		25842 => to_unsigned(20194, LUT_AMPL_WIDTH - 1),
		25843 => to_unsigned(20191, LUT_AMPL_WIDTH - 1),
		25844 => to_unsigned(20189, LUT_AMPL_WIDTH - 1),
		25845 => to_unsigned(20187, LUT_AMPL_WIDTH - 1),
		25846 => to_unsigned(20184, LUT_AMPL_WIDTH - 1),
		25847 => to_unsigned(20182, LUT_AMPL_WIDTH - 1),
		25848 => to_unsigned(20179, LUT_AMPL_WIDTH - 1),
		25849 => to_unsigned(20177, LUT_AMPL_WIDTH - 1),
		25850 => to_unsigned(20174, LUT_AMPL_WIDTH - 1),
		25851 => to_unsigned(20172, LUT_AMPL_WIDTH - 1),
		25852 => to_unsigned(20169, LUT_AMPL_WIDTH - 1),
		25853 => to_unsigned(20167, LUT_AMPL_WIDTH - 1),
		25854 => to_unsigned(20164, LUT_AMPL_WIDTH - 1),
		25855 => to_unsigned(20162, LUT_AMPL_WIDTH - 1),
		25856 => to_unsigned(20159, LUT_AMPL_WIDTH - 1),
		25857 => to_unsigned(20157, LUT_AMPL_WIDTH - 1),
		25858 => to_unsigned(20154, LUT_AMPL_WIDTH - 1),
		25859 => to_unsigned(20152, LUT_AMPL_WIDTH - 1),
		25860 => to_unsigned(20149, LUT_AMPL_WIDTH - 1),
		25861 => to_unsigned(20147, LUT_AMPL_WIDTH - 1),
		25862 => to_unsigned(20144, LUT_AMPL_WIDTH - 1),
		25863 => to_unsigned(20142, LUT_AMPL_WIDTH - 1),
		25864 => to_unsigned(20139, LUT_AMPL_WIDTH - 1),
		25865 => to_unsigned(20137, LUT_AMPL_WIDTH - 1),
		25866 => to_unsigned(20135, LUT_AMPL_WIDTH - 1),
		25867 => to_unsigned(20132, LUT_AMPL_WIDTH - 1),
		25868 => to_unsigned(20130, LUT_AMPL_WIDTH - 1),
		25869 => to_unsigned(20127, LUT_AMPL_WIDTH - 1),
		25870 => to_unsigned(20125, LUT_AMPL_WIDTH - 1),
		25871 => to_unsigned(20122, LUT_AMPL_WIDTH - 1),
		25872 => to_unsigned(20120, LUT_AMPL_WIDTH - 1),
		25873 => to_unsigned(20117, LUT_AMPL_WIDTH - 1),
		25874 => to_unsigned(20115, LUT_AMPL_WIDTH - 1),
		25875 => to_unsigned(20112, LUT_AMPL_WIDTH - 1),
		25876 => to_unsigned(20110, LUT_AMPL_WIDTH - 1),
		25877 => to_unsigned(20107, LUT_AMPL_WIDTH - 1),
		25878 => to_unsigned(20105, LUT_AMPL_WIDTH - 1),
		25879 => to_unsigned(20102, LUT_AMPL_WIDTH - 1),
		25880 => to_unsigned(20100, LUT_AMPL_WIDTH - 1),
		25881 => to_unsigned(20097, LUT_AMPL_WIDTH - 1),
		25882 => to_unsigned(20095, LUT_AMPL_WIDTH - 1),
		25883 => to_unsigned(20092, LUT_AMPL_WIDTH - 1),
		25884 => to_unsigned(20090, LUT_AMPL_WIDTH - 1),
		25885 => to_unsigned(20087, LUT_AMPL_WIDTH - 1),
		25886 => to_unsigned(20085, LUT_AMPL_WIDTH - 1),
		25887 => to_unsigned(20082, LUT_AMPL_WIDTH - 1),
		25888 => to_unsigned(20080, LUT_AMPL_WIDTH - 1),
		25889 => to_unsigned(20077, LUT_AMPL_WIDTH - 1),
		25890 => to_unsigned(20075, LUT_AMPL_WIDTH - 1),
		25891 => to_unsigned(20072, LUT_AMPL_WIDTH - 1),
		25892 => to_unsigned(20070, LUT_AMPL_WIDTH - 1),
		25893 => to_unsigned(20068, LUT_AMPL_WIDTH - 1),
		25894 => to_unsigned(20065, LUT_AMPL_WIDTH - 1),
		25895 => to_unsigned(20063, LUT_AMPL_WIDTH - 1),
		25896 => to_unsigned(20060, LUT_AMPL_WIDTH - 1),
		25897 => to_unsigned(20058, LUT_AMPL_WIDTH - 1),
		25898 => to_unsigned(20055, LUT_AMPL_WIDTH - 1),
		25899 => to_unsigned(20053, LUT_AMPL_WIDTH - 1),
		25900 => to_unsigned(20050, LUT_AMPL_WIDTH - 1),
		25901 => to_unsigned(20048, LUT_AMPL_WIDTH - 1),
		25902 => to_unsigned(20045, LUT_AMPL_WIDTH - 1),
		25903 => to_unsigned(20043, LUT_AMPL_WIDTH - 1),
		25904 => to_unsigned(20040, LUT_AMPL_WIDTH - 1),
		25905 => to_unsigned(20038, LUT_AMPL_WIDTH - 1),
		25906 => to_unsigned(20035, LUT_AMPL_WIDTH - 1),
		25907 => to_unsigned(20033, LUT_AMPL_WIDTH - 1),
		25908 => to_unsigned(20030, LUT_AMPL_WIDTH - 1),
		25909 => to_unsigned(20028, LUT_AMPL_WIDTH - 1),
		25910 => to_unsigned(20025, LUT_AMPL_WIDTH - 1),
		25911 => to_unsigned(20023, LUT_AMPL_WIDTH - 1),
		25912 => to_unsigned(20020, LUT_AMPL_WIDTH - 1),
		25913 => to_unsigned(20018, LUT_AMPL_WIDTH - 1),
		25914 => to_unsigned(20015, LUT_AMPL_WIDTH - 1),
		25915 => to_unsigned(20013, LUT_AMPL_WIDTH - 1),
		25916 => to_unsigned(20010, LUT_AMPL_WIDTH - 1),
		25917 => to_unsigned(20008, LUT_AMPL_WIDTH - 1),
		25918 => to_unsigned(20005, LUT_AMPL_WIDTH - 1),
		25919 => to_unsigned(20003, LUT_AMPL_WIDTH - 1),
		25920 => to_unsigned(20000, LUT_AMPL_WIDTH - 1),
		25921 => to_unsigned(19998, LUT_AMPL_WIDTH - 1),
		25922 => to_unsigned(19995, LUT_AMPL_WIDTH - 1),
		25923 => to_unsigned(19993, LUT_AMPL_WIDTH - 1),
		25924 => to_unsigned(19990, LUT_AMPL_WIDTH - 1),
		25925 => to_unsigned(19988, LUT_AMPL_WIDTH - 1),
		25926 => to_unsigned(19985, LUT_AMPL_WIDTH - 1),
		25927 => to_unsigned(19983, LUT_AMPL_WIDTH - 1),
		25928 => to_unsigned(19981, LUT_AMPL_WIDTH - 1),
		25929 => to_unsigned(19978, LUT_AMPL_WIDTH - 1),
		25930 => to_unsigned(19976, LUT_AMPL_WIDTH - 1),
		25931 => to_unsigned(19973, LUT_AMPL_WIDTH - 1),
		25932 => to_unsigned(19971, LUT_AMPL_WIDTH - 1),
		25933 => to_unsigned(19968, LUT_AMPL_WIDTH - 1),
		25934 => to_unsigned(19966, LUT_AMPL_WIDTH - 1),
		25935 => to_unsigned(19963, LUT_AMPL_WIDTH - 1),
		25936 => to_unsigned(19961, LUT_AMPL_WIDTH - 1),
		25937 => to_unsigned(19958, LUT_AMPL_WIDTH - 1),
		25938 => to_unsigned(19956, LUT_AMPL_WIDTH - 1),
		25939 => to_unsigned(19953, LUT_AMPL_WIDTH - 1),
		25940 => to_unsigned(19951, LUT_AMPL_WIDTH - 1),
		25941 => to_unsigned(19948, LUT_AMPL_WIDTH - 1),
		25942 => to_unsigned(19946, LUT_AMPL_WIDTH - 1),
		25943 => to_unsigned(19943, LUT_AMPL_WIDTH - 1),
		25944 => to_unsigned(19941, LUT_AMPL_WIDTH - 1),
		25945 => to_unsigned(19938, LUT_AMPL_WIDTH - 1),
		25946 => to_unsigned(19936, LUT_AMPL_WIDTH - 1),
		25947 => to_unsigned(19933, LUT_AMPL_WIDTH - 1),
		25948 => to_unsigned(19931, LUT_AMPL_WIDTH - 1),
		25949 => to_unsigned(19928, LUT_AMPL_WIDTH - 1),
		25950 => to_unsigned(19926, LUT_AMPL_WIDTH - 1),
		25951 => to_unsigned(19923, LUT_AMPL_WIDTH - 1),
		25952 => to_unsigned(19921, LUT_AMPL_WIDTH - 1),
		25953 => to_unsigned(19918, LUT_AMPL_WIDTH - 1),
		25954 => to_unsigned(19916, LUT_AMPL_WIDTH - 1),
		25955 => to_unsigned(19913, LUT_AMPL_WIDTH - 1),
		25956 => to_unsigned(19911, LUT_AMPL_WIDTH - 1),
		25957 => to_unsigned(19908, LUT_AMPL_WIDTH - 1),
		25958 => to_unsigned(19906, LUT_AMPL_WIDTH - 1),
		25959 => to_unsigned(19903, LUT_AMPL_WIDTH - 1),
		25960 => to_unsigned(19901, LUT_AMPL_WIDTH - 1),
		25961 => to_unsigned(19898, LUT_AMPL_WIDTH - 1),
		25962 => to_unsigned(19896, LUT_AMPL_WIDTH - 1),
		25963 => to_unsigned(19893, LUT_AMPL_WIDTH - 1),
		25964 => to_unsigned(19891, LUT_AMPL_WIDTH - 1),
		25965 => to_unsigned(19888, LUT_AMPL_WIDTH - 1),
		25966 => to_unsigned(19886, LUT_AMPL_WIDTH - 1),
		25967 => to_unsigned(19883, LUT_AMPL_WIDTH - 1),
		25968 => to_unsigned(19881, LUT_AMPL_WIDTH - 1),
		25969 => to_unsigned(19878, LUT_AMPL_WIDTH - 1),
		25970 => to_unsigned(19876, LUT_AMPL_WIDTH - 1),
		25971 => to_unsigned(19873, LUT_AMPL_WIDTH - 1),
		25972 => to_unsigned(19871, LUT_AMPL_WIDTH - 1),
		25973 => to_unsigned(19868, LUT_AMPL_WIDTH - 1),
		25974 => to_unsigned(19866, LUT_AMPL_WIDTH - 1),
		25975 => to_unsigned(19863, LUT_AMPL_WIDTH - 1),
		25976 => to_unsigned(19861, LUT_AMPL_WIDTH - 1),
		25977 => to_unsigned(19858, LUT_AMPL_WIDTH - 1),
		25978 => to_unsigned(19856, LUT_AMPL_WIDTH - 1),
		25979 => to_unsigned(19853, LUT_AMPL_WIDTH - 1),
		25980 => to_unsigned(19851, LUT_AMPL_WIDTH - 1),
		25981 => to_unsigned(19848, LUT_AMPL_WIDTH - 1),
		25982 => to_unsigned(19846, LUT_AMPL_WIDTH - 1),
		25983 => to_unsigned(19843, LUT_AMPL_WIDTH - 1),
		25984 => to_unsigned(19841, LUT_AMPL_WIDTH - 1),
		25985 => to_unsigned(19838, LUT_AMPL_WIDTH - 1),
		25986 => to_unsigned(19836, LUT_AMPL_WIDTH - 1),
		25987 => to_unsigned(19833, LUT_AMPL_WIDTH - 1),
		25988 => to_unsigned(19831, LUT_AMPL_WIDTH - 1),
		25989 => to_unsigned(19828, LUT_AMPL_WIDTH - 1),
		25990 => to_unsigned(19826, LUT_AMPL_WIDTH - 1),
		25991 => to_unsigned(19823, LUT_AMPL_WIDTH - 1),
		25992 => to_unsigned(19821, LUT_AMPL_WIDTH - 1),
		25993 => to_unsigned(19818, LUT_AMPL_WIDTH - 1),
		25994 => to_unsigned(19816, LUT_AMPL_WIDTH - 1),
		25995 => to_unsigned(19813, LUT_AMPL_WIDTH - 1),
		25996 => to_unsigned(19811, LUT_AMPL_WIDTH - 1),
		25997 => to_unsigned(19808, LUT_AMPL_WIDTH - 1),
		25998 => to_unsigned(19806, LUT_AMPL_WIDTH - 1),
		25999 => to_unsigned(19803, LUT_AMPL_WIDTH - 1),
		26000 => to_unsigned(19801, LUT_AMPL_WIDTH - 1),
		26001 => to_unsigned(19798, LUT_AMPL_WIDTH - 1),
		26002 => to_unsigned(19796, LUT_AMPL_WIDTH - 1),
		26003 => to_unsigned(19793, LUT_AMPL_WIDTH - 1),
		26004 => to_unsigned(19791, LUT_AMPL_WIDTH - 1),
		26005 => to_unsigned(19788, LUT_AMPL_WIDTH - 1),
		26006 => to_unsigned(19786, LUT_AMPL_WIDTH - 1),
		26007 => to_unsigned(19783, LUT_AMPL_WIDTH - 1),
		26008 => to_unsigned(19781, LUT_AMPL_WIDTH - 1),
		26009 => to_unsigned(19778, LUT_AMPL_WIDTH - 1),
		26010 => to_unsigned(19776, LUT_AMPL_WIDTH - 1),
		26011 => to_unsigned(19773, LUT_AMPL_WIDTH - 1),
		26012 => to_unsigned(19771, LUT_AMPL_WIDTH - 1),
		26013 => to_unsigned(19768, LUT_AMPL_WIDTH - 1),
		26014 => to_unsigned(19766, LUT_AMPL_WIDTH - 1),
		26015 => to_unsigned(19763, LUT_AMPL_WIDTH - 1),
		26016 => to_unsigned(19761, LUT_AMPL_WIDTH - 1),
		26017 => to_unsigned(19758, LUT_AMPL_WIDTH - 1),
		26018 => to_unsigned(19756, LUT_AMPL_WIDTH - 1),
		26019 => to_unsigned(19753, LUT_AMPL_WIDTH - 1),
		26020 => to_unsigned(19751, LUT_AMPL_WIDTH - 1),
		26021 => to_unsigned(19748, LUT_AMPL_WIDTH - 1),
		26022 => to_unsigned(19746, LUT_AMPL_WIDTH - 1),
		26023 => to_unsigned(19743, LUT_AMPL_WIDTH - 1),
		26024 => to_unsigned(19741, LUT_AMPL_WIDTH - 1),
		26025 => to_unsigned(19738, LUT_AMPL_WIDTH - 1),
		26026 => to_unsigned(19736, LUT_AMPL_WIDTH - 1),
		26027 => to_unsigned(19733, LUT_AMPL_WIDTH - 1),
		26028 => to_unsigned(19731, LUT_AMPL_WIDTH - 1),
		26029 => to_unsigned(19728, LUT_AMPL_WIDTH - 1),
		26030 => to_unsigned(19726, LUT_AMPL_WIDTH - 1),
		26031 => to_unsigned(19723, LUT_AMPL_WIDTH - 1),
		26032 => to_unsigned(19721, LUT_AMPL_WIDTH - 1),
		26033 => to_unsigned(19718, LUT_AMPL_WIDTH - 1),
		26034 => to_unsigned(19716, LUT_AMPL_WIDTH - 1),
		26035 => to_unsigned(19713, LUT_AMPL_WIDTH - 1),
		26036 => to_unsigned(19711, LUT_AMPL_WIDTH - 1),
		26037 => to_unsigned(19708, LUT_AMPL_WIDTH - 1),
		26038 => to_unsigned(19706, LUT_AMPL_WIDTH - 1),
		26039 => to_unsigned(19703, LUT_AMPL_WIDTH - 1),
		26040 => to_unsigned(19700, LUT_AMPL_WIDTH - 1),
		26041 => to_unsigned(19698, LUT_AMPL_WIDTH - 1),
		26042 => to_unsigned(19695, LUT_AMPL_WIDTH - 1),
		26043 => to_unsigned(19693, LUT_AMPL_WIDTH - 1),
		26044 => to_unsigned(19690, LUT_AMPL_WIDTH - 1),
		26045 => to_unsigned(19688, LUT_AMPL_WIDTH - 1),
		26046 => to_unsigned(19685, LUT_AMPL_WIDTH - 1),
		26047 => to_unsigned(19683, LUT_AMPL_WIDTH - 1),
		26048 => to_unsigned(19680, LUT_AMPL_WIDTH - 1),
		26049 => to_unsigned(19678, LUT_AMPL_WIDTH - 1),
		26050 => to_unsigned(19675, LUT_AMPL_WIDTH - 1),
		26051 => to_unsigned(19673, LUT_AMPL_WIDTH - 1),
		26052 => to_unsigned(19670, LUT_AMPL_WIDTH - 1),
		26053 => to_unsigned(19668, LUT_AMPL_WIDTH - 1),
		26054 => to_unsigned(19665, LUT_AMPL_WIDTH - 1),
		26055 => to_unsigned(19663, LUT_AMPL_WIDTH - 1),
		26056 => to_unsigned(19660, LUT_AMPL_WIDTH - 1),
		26057 => to_unsigned(19658, LUT_AMPL_WIDTH - 1),
		26058 => to_unsigned(19655, LUT_AMPL_WIDTH - 1),
		26059 => to_unsigned(19653, LUT_AMPL_WIDTH - 1),
		26060 => to_unsigned(19650, LUT_AMPL_WIDTH - 1),
		26061 => to_unsigned(19648, LUT_AMPL_WIDTH - 1),
		26062 => to_unsigned(19645, LUT_AMPL_WIDTH - 1),
		26063 => to_unsigned(19643, LUT_AMPL_WIDTH - 1),
		26064 => to_unsigned(19640, LUT_AMPL_WIDTH - 1),
		26065 => to_unsigned(19638, LUT_AMPL_WIDTH - 1),
		26066 => to_unsigned(19635, LUT_AMPL_WIDTH - 1),
		26067 => to_unsigned(19633, LUT_AMPL_WIDTH - 1),
		26068 => to_unsigned(19630, LUT_AMPL_WIDTH - 1),
		26069 => to_unsigned(19628, LUT_AMPL_WIDTH - 1),
		26070 => to_unsigned(19625, LUT_AMPL_WIDTH - 1),
		26071 => to_unsigned(19623, LUT_AMPL_WIDTH - 1),
		26072 => to_unsigned(19620, LUT_AMPL_WIDTH - 1),
		26073 => to_unsigned(19618, LUT_AMPL_WIDTH - 1),
		26074 => to_unsigned(19615, LUT_AMPL_WIDTH - 1),
		26075 => to_unsigned(19613, LUT_AMPL_WIDTH - 1),
		26076 => to_unsigned(19610, LUT_AMPL_WIDTH - 1),
		26077 => to_unsigned(19607, LUT_AMPL_WIDTH - 1),
		26078 => to_unsigned(19605, LUT_AMPL_WIDTH - 1),
		26079 => to_unsigned(19602, LUT_AMPL_WIDTH - 1),
		26080 => to_unsigned(19600, LUT_AMPL_WIDTH - 1),
		26081 => to_unsigned(19597, LUT_AMPL_WIDTH - 1),
		26082 => to_unsigned(19595, LUT_AMPL_WIDTH - 1),
		26083 => to_unsigned(19592, LUT_AMPL_WIDTH - 1),
		26084 => to_unsigned(19590, LUT_AMPL_WIDTH - 1),
		26085 => to_unsigned(19587, LUT_AMPL_WIDTH - 1),
		26086 => to_unsigned(19585, LUT_AMPL_WIDTH - 1),
		26087 => to_unsigned(19582, LUT_AMPL_WIDTH - 1),
		26088 => to_unsigned(19580, LUT_AMPL_WIDTH - 1),
		26089 => to_unsigned(19577, LUT_AMPL_WIDTH - 1),
		26090 => to_unsigned(19575, LUT_AMPL_WIDTH - 1),
		26091 => to_unsigned(19572, LUT_AMPL_WIDTH - 1),
		26092 => to_unsigned(19570, LUT_AMPL_WIDTH - 1),
		26093 => to_unsigned(19567, LUT_AMPL_WIDTH - 1),
		26094 => to_unsigned(19565, LUT_AMPL_WIDTH - 1),
		26095 => to_unsigned(19562, LUT_AMPL_WIDTH - 1),
		26096 => to_unsigned(19560, LUT_AMPL_WIDTH - 1),
		26097 => to_unsigned(19557, LUT_AMPL_WIDTH - 1),
		26098 => to_unsigned(19555, LUT_AMPL_WIDTH - 1),
		26099 => to_unsigned(19552, LUT_AMPL_WIDTH - 1),
		26100 => to_unsigned(19550, LUT_AMPL_WIDTH - 1),
		26101 => to_unsigned(19547, LUT_AMPL_WIDTH - 1),
		26102 => to_unsigned(19545, LUT_AMPL_WIDTH - 1),
		26103 => to_unsigned(19542, LUT_AMPL_WIDTH - 1),
		26104 => to_unsigned(19539, LUT_AMPL_WIDTH - 1),
		26105 => to_unsigned(19537, LUT_AMPL_WIDTH - 1),
		26106 => to_unsigned(19534, LUT_AMPL_WIDTH - 1),
		26107 => to_unsigned(19532, LUT_AMPL_WIDTH - 1),
		26108 => to_unsigned(19529, LUT_AMPL_WIDTH - 1),
		26109 => to_unsigned(19527, LUT_AMPL_WIDTH - 1),
		26110 => to_unsigned(19524, LUT_AMPL_WIDTH - 1),
		26111 => to_unsigned(19522, LUT_AMPL_WIDTH - 1),
		26112 => to_unsigned(19519, LUT_AMPL_WIDTH - 1),
		26113 => to_unsigned(19517, LUT_AMPL_WIDTH - 1),
		26114 => to_unsigned(19514, LUT_AMPL_WIDTH - 1),
		26115 => to_unsigned(19512, LUT_AMPL_WIDTH - 1),
		26116 => to_unsigned(19509, LUT_AMPL_WIDTH - 1),
		26117 => to_unsigned(19507, LUT_AMPL_WIDTH - 1),
		26118 => to_unsigned(19504, LUT_AMPL_WIDTH - 1),
		26119 => to_unsigned(19502, LUT_AMPL_WIDTH - 1),
		26120 => to_unsigned(19499, LUT_AMPL_WIDTH - 1),
		26121 => to_unsigned(19497, LUT_AMPL_WIDTH - 1),
		26122 => to_unsigned(19494, LUT_AMPL_WIDTH - 1),
		26123 => to_unsigned(19492, LUT_AMPL_WIDTH - 1),
		26124 => to_unsigned(19489, LUT_AMPL_WIDTH - 1),
		26125 => to_unsigned(19486, LUT_AMPL_WIDTH - 1),
		26126 => to_unsigned(19484, LUT_AMPL_WIDTH - 1),
		26127 => to_unsigned(19481, LUT_AMPL_WIDTH - 1),
		26128 => to_unsigned(19479, LUT_AMPL_WIDTH - 1),
		26129 => to_unsigned(19476, LUT_AMPL_WIDTH - 1),
		26130 => to_unsigned(19474, LUT_AMPL_WIDTH - 1),
		26131 => to_unsigned(19471, LUT_AMPL_WIDTH - 1),
		26132 => to_unsigned(19469, LUT_AMPL_WIDTH - 1),
		26133 => to_unsigned(19466, LUT_AMPL_WIDTH - 1),
		26134 => to_unsigned(19464, LUT_AMPL_WIDTH - 1),
		26135 => to_unsigned(19461, LUT_AMPL_WIDTH - 1),
		26136 => to_unsigned(19459, LUT_AMPL_WIDTH - 1),
		26137 => to_unsigned(19456, LUT_AMPL_WIDTH - 1),
		26138 => to_unsigned(19454, LUT_AMPL_WIDTH - 1),
		26139 => to_unsigned(19451, LUT_AMPL_WIDTH - 1),
		26140 => to_unsigned(19449, LUT_AMPL_WIDTH - 1),
		26141 => to_unsigned(19446, LUT_AMPL_WIDTH - 1),
		26142 => to_unsigned(19444, LUT_AMPL_WIDTH - 1),
		26143 => to_unsigned(19441, LUT_AMPL_WIDTH - 1),
		26144 => to_unsigned(19438, LUT_AMPL_WIDTH - 1),
		26145 => to_unsigned(19436, LUT_AMPL_WIDTH - 1),
		26146 => to_unsigned(19433, LUT_AMPL_WIDTH - 1),
		26147 => to_unsigned(19431, LUT_AMPL_WIDTH - 1),
		26148 => to_unsigned(19428, LUT_AMPL_WIDTH - 1),
		26149 => to_unsigned(19426, LUT_AMPL_WIDTH - 1),
		26150 => to_unsigned(19423, LUT_AMPL_WIDTH - 1),
		26151 => to_unsigned(19421, LUT_AMPL_WIDTH - 1),
		26152 => to_unsigned(19418, LUT_AMPL_WIDTH - 1),
		26153 => to_unsigned(19416, LUT_AMPL_WIDTH - 1),
		26154 => to_unsigned(19413, LUT_AMPL_WIDTH - 1),
		26155 => to_unsigned(19411, LUT_AMPL_WIDTH - 1),
		26156 => to_unsigned(19408, LUT_AMPL_WIDTH - 1),
		26157 => to_unsigned(19406, LUT_AMPL_WIDTH - 1),
		26158 => to_unsigned(19403, LUT_AMPL_WIDTH - 1),
		26159 => to_unsigned(19400, LUT_AMPL_WIDTH - 1),
		26160 => to_unsigned(19398, LUT_AMPL_WIDTH - 1),
		26161 => to_unsigned(19395, LUT_AMPL_WIDTH - 1),
		26162 => to_unsigned(19393, LUT_AMPL_WIDTH - 1),
		26163 => to_unsigned(19390, LUT_AMPL_WIDTH - 1),
		26164 => to_unsigned(19388, LUT_AMPL_WIDTH - 1),
		26165 => to_unsigned(19385, LUT_AMPL_WIDTH - 1),
		26166 => to_unsigned(19383, LUT_AMPL_WIDTH - 1),
		26167 => to_unsigned(19380, LUT_AMPL_WIDTH - 1),
		26168 => to_unsigned(19378, LUT_AMPL_WIDTH - 1),
		26169 => to_unsigned(19375, LUT_AMPL_WIDTH - 1),
		26170 => to_unsigned(19373, LUT_AMPL_WIDTH - 1),
		26171 => to_unsigned(19370, LUT_AMPL_WIDTH - 1),
		26172 => to_unsigned(19368, LUT_AMPL_WIDTH - 1),
		26173 => to_unsigned(19365, LUT_AMPL_WIDTH - 1),
		26174 => to_unsigned(19362, LUT_AMPL_WIDTH - 1),
		26175 => to_unsigned(19360, LUT_AMPL_WIDTH - 1),
		26176 => to_unsigned(19357, LUT_AMPL_WIDTH - 1),
		26177 => to_unsigned(19355, LUT_AMPL_WIDTH - 1),
		26178 => to_unsigned(19352, LUT_AMPL_WIDTH - 1),
		26179 => to_unsigned(19350, LUT_AMPL_WIDTH - 1),
		26180 => to_unsigned(19347, LUT_AMPL_WIDTH - 1),
		26181 => to_unsigned(19345, LUT_AMPL_WIDTH - 1),
		26182 => to_unsigned(19342, LUT_AMPL_WIDTH - 1),
		26183 => to_unsigned(19340, LUT_AMPL_WIDTH - 1),
		26184 => to_unsigned(19337, LUT_AMPL_WIDTH - 1),
		26185 => to_unsigned(19335, LUT_AMPL_WIDTH - 1),
		26186 => to_unsigned(19332, LUT_AMPL_WIDTH - 1),
		26187 => to_unsigned(19330, LUT_AMPL_WIDTH - 1),
		26188 => to_unsigned(19327, LUT_AMPL_WIDTH - 1),
		26189 => to_unsigned(19324, LUT_AMPL_WIDTH - 1),
		26190 => to_unsigned(19322, LUT_AMPL_WIDTH - 1),
		26191 => to_unsigned(19319, LUT_AMPL_WIDTH - 1),
		26192 => to_unsigned(19317, LUT_AMPL_WIDTH - 1),
		26193 => to_unsigned(19314, LUT_AMPL_WIDTH - 1),
		26194 => to_unsigned(19312, LUT_AMPL_WIDTH - 1),
		26195 => to_unsigned(19309, LUT_AMPL_WIDTH - 1),
		26196 => to_unsigned(19307, LUT_AMPL_WIDTH - 1),
		26197 => to_unsigned(19304, LUT_AMPL_WIDTH - 1),
		26198 => to_unsigned(19302, LUT_AMPL_WIDTH - 1),
		26199 => to_unsigned(19299, LUT_AMPL_WIDTH - 1),
		26200 => to_unsigned(19297, LUT_AMPL_WIDTH - 1),
		26201 => to_unsigned(19294, LUT_AMPL_WIDTH - 1),
		26202 => to_unsigned(19291, LUT_AMPL_WIDTH - 1),
		26203 => to_unsigned(19289, LUT_AMPL_WIDTH - 1),
		26204 => to_unsigned(19286, LUT_AMPL_WIDTH - 1),
		26205 => to_unsigned(19284, LUT_AMPL_WIDTH - 1),
		26206 => to_unsigned(19281, LUT_AMPL_WIDTH - 1),
		26207 => to_unsigned(19279, LUT_AMPL_WIDTH - 1),
		26208 => to_unsigned(19276, LUT_AMPL_WIDTH - 1),
		26209 => to_unsigned(19274, LUT_AMPL_WIDTH - 1),
		26210 => to_unsigned(19271, LUT_AMPL_WIDTH - 1),
		26211 => to_unsigned(19269, LUT_AMPL_WIDTH - 1),
		26212 => to_unsigned(19266, LUT_AMPL_WIDTH - 1),
		26213 => to_unsigned(19264, LUT_AMPL_WIDTH - 1),
		26214 => to_unsigned(19261, LUT_AMPL_WIDTH - 1),
		26215 => to_unsigned(19258, LUT_AMPL_WIDTH - 1),
		26216 => to_unsigned(19256, LUT_AMPL_WIDTH - 1),
		26217 => to_unsigned(19253, LUT_AMPL_WIDTH - 1),
		26218 => to_unsigned(19251, LUT_AMPL_WIDTH - 1),
		26219 => to_unsigned(19248, LUT_AMPL_WIDTH - 1),
		26220 => to_unsigned(19246, LUT_AMPL_WIDTH - 1),
		26221 => to_unsigned(19243, LUT_AMPL_WIDTH - 1),
		26222 => to_unsigned(19241, LUT_AMPL_WIDTH - 1),
		26223 => to_unsigned(19238, LUT_AMPL_WIDTH - 1),
		26224 => to_unsigned(19236, LUT_AMPL_WIDTH - 1),
		26225 => to_unsigned(19233, LUT_AMPL_WIDTH - 1),
		26226 => to_unsigned(19230, LUT_AMPL_WIDTH - 1),
		26227 => to_unsigned(19228, LUT_AMPL_WIDTH - 1),
		26228 => to_unsigned(19225, LUT_AMPL_WIDTH - 1),
		26229 => to_unsigned(19223, LUT_AMPL_WIDTH - 1),
		26230 => to_unsigned(19220, LUT_AMPL_WIDTH - 1),
		26231 => to_unsigned(19218, LUT_AMPL_WIDTH - 1),
		26232 => to_unsigned(19215, LUT_AMPL_WIDTH - 1),
		26233 => to_unsigned(19213, LUT_AMPL_WIDTH - 1),
		26234 => to_unsigned(19210, LUT_AMPL_WIDTH - 1),
		26235 => to_unsigned(19208, LUT_AMPL_WIDTH - 1),
		26236 => to_unsigned(19205, LUT_AMPL_WIDTH - 1),
		26237 => to_unsigned(19202, LUT_AMPL_WIDTH - 1),
		26238 => to_unsigned(19200, LUT_AMPL_WIDTH - 1),
		26239 => to_unsigned(19197, LUT_AMPL_WIDTH - 1),
		26240 => to_unsigned(19195, LUT_AMPL_WIDTH - 1),
		26241 => to_unsigned(19192, LUT_AMPL_WIDTH - 1),
		26242 => to_unsigned(19190, LUT_AMPL_WIDTH - 1),
		26243 => to_unsigned(19187, LUT_AMPL_WIDTH - 1),
		26244 => to_unsigned(19185, LUT_AMPL_WIDTH - 1),
		26245 => to_unsigned(19182, LUT_AMPL_WIDTH - 1),
		26246 => to_unsigned(19180, LUT_AMPL_WIDTH - 1),
		26247 => to_unsigned(19177, LUT_AMPL_WIDTH - 1),
		26248 => to_unsigned(19174, LUT_AMPL_WIDTH - 1),
		26249 => to_unsigned(19172, LUT_AMPL_WIDTH - 1),
		26250 => to_unsigned(19169, LUT_AMPL_WIDTH - 1),
		26251 => to_unsigned(19167, LUT_AMPL_WIDTH - 1),
		26252 => to_unsigned(19164, LUT_AMPL_WIDTH - 1),
		26253 => to_unsigned(19162, LUT_AMPL_WIDTH - 1),
		26254 => to_unsigned(19159, LUT_AMPL_WIDTH - 1),
		26255 => to_unsigned(19157, LUT_AMPL_WIDTH - 1),
		26256 => to_unsigned(19154, LUT_AMPL_WIDTH - 1),
		26257 => to_unsigned(19152, LUT_AMPL_WIDTH - 1),
		26258 => to_unsigned(19149, LUT_AMPL_WIDTH - 1),
		26259 => to_unsigned(19146, LUT_AMPL_WIDTH - 1),
		26260 => to_unsigned(19144, LUT_AMPL_WIDTH - 1),
		26261 => to_unsigned(19141, LUT_AMPL_WIDTH - 1),
		26262 => to_unsigned(19139, LUT_AMPL_WIDTH - 1),
		26263 => to_unsigned(19136, LUT_AMPL_WIDTH - 1),
		26264 => to_unsigned(19134, LUT_AMPL_WIDTH - 1),
		26265 => to_unsigned(19131, LUT_AMPL_WIDTH - 1),
		26266 => to_unsigned(19129, LUT_AMPL_WIDTH - 1),
		26267 => to_unsigned(19126, LUT_AMPL_WIDTH - 1),
		26268 => to_unsigned(19123, LUT_AMPL_WIDTH - 1),
		26269 => to_unsigned(19121, LUT_AMPL_WIDTH - 1),
		26270 => to_unsigned(19118, LUT_AMPL_WIDTH - 1),
		26271 => to_unsigned(19116, LUT_AMPL_WIDTH - 1),
		26272 => to_unsigned(19113, LUT_AMPL_WIDTH - 1),
		26273 => to_unsigned(19111, LUT_AMPL_WIDTH - 1),
		26274 => to_unsigned(19108, LUT_AMPL_WIDTH - 1),
		26275 => to_unsigned(19106, LUT_AMPL_WIDTH - 1),
		26276 => to_unsigned(19103, LUT_AMPL_WIDTH - 1),
		26277 => to_unsigned(19101, LUT_AMPL_WIDTH - 1),
		26278 => to_unsigned(19098, LUT_AMPL_WIDTH - 1),
		26279 => to_unsigned(19095, LUT_AMPL_WIDTH - 1),
		26280 => to_unsigned(19093, LUT_AMPL_WIDTH - 1),
		26281 => to_unsigned(19090, LUT_AMPL_WIDTH - 1),
		26282 => to_unsigned(19088, LUT_AMPL_WIDTH - 1),
		26283 => to_unsigned(19085, LUT_AMPL_WIDTH - 1),
		26284 => to_unsigned(19083, LUT_AMPL_WIDTH - 1),
		26285 => to_unsigned(19080, LUT_AMPL_WIDTH - 1),
		26286 => to_unsigned(19078, LUT_AMPL_WIDTH - 1),
		26287 => to_unsigned(19075, LUT_AMPL_WIDTH - 1),
		26288 => to_unsigned(19072, LUT_AMPL_WIDTH - 1),
		26289 => to_unsigned(19070, LUT_AMPL_WIDTH - 1),
		26290 => to_unsigned(19067, LUT_AMPL_WIDTH - 1),
		26291 => to_unsigned(19065, LUT_AMPL_WIDTH - 1),
		26292 => to_unsigned(19062, LUT_AMPL_WIDTH - 1),
		26293 => to_unsigned(19060, LUT_AMPL_WIDTH - 1),
		26294 => to_unsigned(19057, LUT_AMPL_WIDTH - 1),
		26295 => to_unsigned(19055, LUT_AMPL_WIDTH - 1),
		26296 => to_unsigned(19052, LUT_AMPL_WIDTH - 1),
		26297 => to_unsigned(19049, LUT_AMPL_WIDTH - 1),
		26298 => to_unsigned(19047, LUT_AMPL_WIDTH - 1),
		26299 => to_unsigned(19044, LUT_AMPL_WIDTH - 1),
		26300 => to_unsigned(19042, LUT_AMPL_WIDTH - 1),
		26301 => to_unsigned(19039, LUT_AMPL_WIDTH - 1),
		26302 => to_unsigned(19037, LUT_AMPL_WIDTH - 1),
		26303 => to_unsigned(19034, LUT_AMPL_WIDTH - 1),
		26304 => to_unsigned(19032, LUT_AMPL_WIDTH - 1),
		26305 => to_unsigned(19029, LUT_AMPL_WIDTH - 1),
		26306 => to_unsigned(19026, LUT_AMPL_WIDTH - 1),
		26307 => to_unsigned(19024, LUT_AMPL_WIDTH - 1),
		26308 => to_unsigned(19021, LUT_AMPL_WIDTH - 1),
		26309 => to_unsigned(19019, LUT_AMPL_WIDTH - 1),
		26310 => to_unsigned(19016, LUT_AMPL_WIDTH - 1),
		26311 => to_unsigned(19014, LUT_AMPL_WIDTH - 1),
		26312 => to_unsigned(19011, LUT_AMPL_WIDTH - 1),
		26313 => to_unsigned(19009, LUT_AMPL_WIDTH - 1),
		26314 => to_unsigned(19006, LUT_AMPL_WIDTH - 1),
		26315 => to_unsigned(19003, LUT_AMPL_WIDTH - 1),
		26316 => to_unsigned(19001, LUT_AMPL_WIDTH - 1),
		26317 => to_unsigned(18998, LUT_AMPL_WIDTH - 1),
		26318 => to_unsigned(18996, LUT_AMPL_WIDTH - 1),
		26319 => to_unsigned(18993, LUT_AMPL_WIDTH - 1),
		26320 => to_unsigned(18991, LUT_AMPL_WIDTH - 1),
		26321 => to_unsigned(18988, LUT_AMPL_WIDTH - 1),
		26322 => to_unsigned(18985, LUT_AMPL_WIDTH - 1),
		26323 => to_unsigned(18983, LUT_AMPL_WIDTH - 1),
		26324 => to_unsigned(18980, LUT_AMPL_WIDTH - 1),
		26325 => to_unsigned(18978, LUT_AMPL_WIDTH - 1),
		26326 => to_unsigned(18975, LUT_AMPL_WIDTH - 1),
		26327 => to_unsigned(18973, LUT_AMPL_WIDTH - 1),
		26328 => to_unsigned(18970, LUT_AMPL_WIDTH - 1),
		26329 => to_unsigned(18968, LUT_AMPL_WIDTH - 1),
		26330 => to_unsigned(18965, LUT_AMPL_WIDTH - 1),
		26331 => to_unsigned(18962, LUT_AMPL_WIDTH - 1),
		26332 => to_unsigned(18960, LUT_AMPL_WIDTH - 1),
		26333 => to_unsigned(18957, LUT_AMPL_WIDTH - 1),
		26334 => to_unsigned(18955, LUT_AMPL_WIDTH - 1),
		26335 => to_unsigned(18952, LUT_AMPL_WIDTH - 1),
		26336 => to_unsigned(18950, LUT_AMPL_WIDTH - 1),
		26337 => to_unsigned(18947, LUT_AMPL_WIDTH - 1),
		26338 => to_unsigned(18944, LUT_AMPL_WIDTH - 1),
		26339 => to_unsigned(18942, LUT_AMPL_WIDTH - 1),
		26340 => to_unsigned(18939, LUT_AMPL_WIDTH - 1),
		26341 => to_unsigned(18937, LUT_AMPL_WIDTH - 1),
		26342 => to_unsigned(18934, LUT_AMPL_WIDTH - 1),
		26343 => to_unsigned(18932, LUT_AMPL_WIDTH - 1),
		26344 => to_unsigned(18929, LUT_AMPL_WIDTH - 1),
		26345 => to_unsigned(18927, LUT_AMPL_WIDTH - 1),
		26346 => to_unsigned(18924, LUT_AMPL_WIDTH - 1),
		26347 => to_unsigned(18921, LUT_AMPL_WIDTH - 1),
		26348 => to_unsigned(18919, LUT_AMPL_WIDTH - 1),
		26349 => to_unsigned(18916, LUT_AMPL_WIDTH - 1),
		26350 => to_unsigned(18914, LUT_AMPL_WIDTH - 1),
		26351 => to_unsigned(18911, LUT_AMPL_WIDTH - 1),
		26352 => to_unsigned(18909, LUT_AMPL_WIDTH - 1),
		26353 => to_unsigned(18906, LUT_AMPL_WIDTH - 1),
		26354 => to_unsigned(18903, LUT_AMPL_WIDTH - 1),
		26355 => to_unsigned(18901, LUT_AMPL_WIDTH - 1),
		26356 => to_unsigned(18898, LUT_AMPL_WIDTH - 1),
		26357 => to_unsigned(18896, LUT_AMPL_WIDTH - 1),
		26358 => to_unsigned(18893, LUT_AMPL_WIDTH - 1),
		26359 => to_unsigned(18891, LUT_AMPL_WIDTH - 1),
		26360 => to_unsigned(18888, LUT_AMPL_WIDTH - 1),
		26361 => to_unsigned(18885, LUT_AMPL_WIDTH - 1),
		26362 => to_unsigned(18883, LUT_AMPL_WIDTH - 1),
		26363 => to_unsigned(18880, LUT_AMPL_WIDTH - 1),
		26364 => to_unsigned(18878, LUT_AMPL_WIDTH - 1),
		26365 => to_unsigned(18875, LUT_AMPL_WIDTH - 1),
		26366 => to_unsigned(18873, LUT_AMPL_WIDTH - 1),
		26367 => to_unsigned(18870, LUT_AMPL_WIDTH - 1),
		26368 => to_unsigned(18868, LUT_AMPL_WIDTH - 1),
		26369 => to_unsigned(18865, LUT_AMPL_WIDTH - 1),
		26370 => to_unsigned(18862, LUT_AMPL_WIDTH - 1),
		26371 => to_unsigned(18860, LUT_AMPL_WIDTH - 1),
		26372 => to_unsigned(18857, LUT_AMPL_WIDTH - 1),
		26373 => to_unsigned(18855, LUT_AMPL_WIDTH - 1),
		26374 => to_unsigned(18852, LUT_AMPL_WIDTH - 1),
		26375 => to_unsigned(18850, LUT_AMPL_WIDTH - 1),
		26376 => to_unsigned(18847, LUT_AMPL_WIDTH - 1),
		26377 => to_unsigned(18844, LUT_AMPL_WIDTH - 1),
		26378 => to_unsigned(18842, LUT_AMPL_WIDTH - 1),
		26379 => to_unsigned(18839, LUT_AMPL_WIDTH - 1),
		26380 => to_unsigned(18837, LUT_AMPL_WIDTH - 1),
		26381 => to_unsigned(18834, LUT_AMPL_WIDTH - 1),
		26382 => to_unsigned(18832, LUT_AMPL_WIDTH - 1),
		26383 => to_unsigned(18829, LUT_AMPL_WIDTH - 1),
		26384 => to_unsigned(18826, LUT_AMPL_WIDTH - 1),
		26385 => to_unsigned(18824, LUT_AMPL_WIDTH - 1),
		26386 => to_unsigned(18821, LUT_AMPL_WIDTH - 1),
		26387 => to_unsigned(18819, LUT_AMPL_WIDTH - 1),
		26388 => to_unsigned(18816, LUT_AMPL_WIDTH - 1),
		26389 => to_unsigned(18814, LUT_AMPL_WIDTH - 1),
		26390 => to_unsigned(18811, LUT_AMPL_WIDTH - 1),
		26391 => to_unsigned(18808, LUT_AMPL_WIDTH - 1),
		26392 => to_unsigned(18806, LUT_AMPL_WIDTH - 1),
		26393 => to_unsigned(18803, LUT_AMPL_WIDTH - 1),
		26394 => to_unsigned(18801, LUT_AMPL_WIDTH - 1),
		26395 => to_unsigned(18798, LUT_AMPL_WIDTH - 1),
		26396 => to_unsigned(18796, LUT_AMPL_WIDTH - 1),
		26397 => to_unsigned(18793, LUT_AMPL_WIDTH - 1),
		26398 => to_unsigned(18790, LUT_AMPL_WIDTH - 1),
		26399 => to_unsigned(18788, LUT_AMPL_WIDTH - 1),
		26400 => to_unsigned(18785, LUT_AMPL_WIDTH - 1),
		26401 => to_unsigned(18783, LUT_AMPL_WIDTH - 1),
		26402 => to_unsigned(18780, LUT_AMPL_WIDTH - 1),
		26403 => to_unsigned(18778, LUT_AMPL_WIDTH - 1),
		26404 => to_unsigned(18775, LUT_AMPL_WIDTH - 1),
		26405 => to_unsigned(18772, LUT_AMPL_WIDTH - 1),
		26406 => to_unsigned(18770, LUT_AMPL_WIDTH - 1),
		26407 => to_unsigned(18767, LUT_AMPL_WIDTH - 1),
		26408 => to_unsigned(18765, LUT_AMPL_WIDTH - 1),
		26409 => to_unsigned(18762, LUT_AMPL_WIDTH - 1),
		26410 => to_unsigned(18759, LUT_AMPL_WIDTH - 1),
		26411 => to_unsigned(18757, LUT_AMPL_WIDTH - 1),
		26412 => to_unsigned(18754, LUT_AMPL_WIDTH - 1),
		26413 => to_unsigned(18752, LUT_AMPL_WIDTH - 1),
		26414 => to_unsigned(18749, LUT_AMPL_WIDTH - 1),
		26415 => to_unsigned(18747, LUT_AMPL_WIDTH - 1),
		26416 => to_unsigned(18744, LUT_AMPL_WIDTH - 1),
		26417 => to_unsigned(18741, LUT_AMPL_WIDTH - 1),
		26418 => to_unsigned(18739, LUT_AMPL_WIDTH - 1),
		26419 => to_unsigned(18736, LUT_AMPL_WIDTH - 1),
		26420 => to_unsigned(18734, LUT_AMPL_WIDTH - 1),
		26421 => to_unsigned(18731, LUT_AMPL_WIDTH - 1),
		26422 => to_unsigned(18729, LUT_AMPL_WIDTH - 1),
		26423 => to_unsigned(18726, LUT_AMPL_WIDTH - 1),
		26424 => to_unsigned(18723, LUT_AMPL_WIDTH - 1),
		26425 => to_unsigned(18721, LUT_AMPL_WIDTH - 1),
		26426 => to_unsigned(18718, LUT_AMPL_WIDTH - 1),
		26427 => to_unsigned(18716, LUT_AMPL_WIDTH - 1),
		26428 => to_unsigned(18713, LUT_AMPL_WIDTH - 1),
		26429 => to_unsigned(18711, LUT_AMPL_WIDTH - 1),
		26430 => to_unsigned(18708, LUT_AMPL_WIDTH - 1),
		26431 => to_unsigned(18705, LUT_AMPL_WIDTH - 1),
		26432 => to_unsigned(18703, LUT_AMPL_WIDTH - 1),
		26433 => to_unsigned(18700, LUT_AMPL_WIDTH - 1),
		26434 => to_unsigned(18698, LUT_AMPL_WIDTH - 1),
		26435 => to_unsigned(18695, LUT_AMPL_WIDTH - 1),
		26436 => to_unsigned(18692, LUT_AMPL_WIDTH - 1),
		26437 => to_unsigned(18690, LUT_AMPL_WIDTH - 1),
		26438 => to_unsigned(18687, LUT_AMPL_WIDTH - 1),
		26439 => to_unsigned(18685, LUT_AMPL_WIDTH - 1),
		26440 => to_unsigned(18682, LUT_AMPL_WIDTH - 1),
		26441 => to_unsigned(18680, LUT_AMPL_WIDTH - 1),
		26442 => to_unsigned(18677, LUT_AMPL_WIDTH - 1),
		26443 => to_unsigned(18674, LUT_AMPL_WIDTH - 1),
		26444 => to_unsigned(18672, LUT_AMPL_WIDTH - 1),
		26445 => to_unsigned(18669, LUT_AMPL_WIDTH - 1),
		26446 => to_unsigned(18667, LUT_AMPL_WIDTH - 1),
		26447 => to_unsigned(18664, LUT_AMPL_WIDTH - 1),
		26448 => to_unsigned(18661, LUT_AMPL_WIDTH - 1),
		26449 => to_unsigned(18659, LUT_AMPL_WIDTH - 1),
		26450 => to_unsigned(18656, LUT_AMPL_WIDTH - 1),
		26451 => to_unsigned(18654, LUT_AMPL_WIDTH - 1),
		26452 => to_unsigned(18651, LUT_AMPL_WIDTH - 1),
		26453 => to_unsigned(18649, LUT_AMPL_WIDTH - 1),
		26454 => to_unsigned(18646, LUT_AMPL_WIDTH - 1),
		26455 => to_unsigned(18643, LUT_AMPL_WIDTH - 1),
		26456 => to_unsigned(18641, LUT_AMPL_WIDTH - 1),
		26457 => to_unsigned(18638, LUT_AMPL_WIDTH - 1),
		26458 => to_unsigned(18636, LUT_AMPL_WIDTH - 1),
		26459 => to_unsigned(18633, LUT_AMPL_WIDTH - 1),
		26460 => to_unsigned(18630, LUT_AMPL_WIDTH - 1),
		26461 => to_unsigned(18628, LUT_AMPL_WIDTH - 1),
		26462 => to_unsigned(18625, LUT_AMPL_WIDTH - 1),
		26463 => to_unsigned(18623, LUT_AMPL_WIDTH - 1),
		26464 => to_unsigned(18620, LUT_AMPL_WIDTH - 1),
		26465 => to_unsigned(18618, LUT_AMPL_WIDTH - 1),
		26466 => to_unsigned(18615, LUT_AMPL_WIDTH - 1),
		26467 => to_unsigned(18612, LUT_AMPL_WIDTH - 1),
		26468 => to_unsigned(18610, LUT_AMPL_WIDTH - 1),
		26469 => to_unsigned(18607, LUT_AMPL_WIDTH - 1),
		26470 => to_unsigned(18605, LUT_AMPL_WIDTH - 1),
		26471 => to_unsigned(18602, LUT_AMPL_WIDTH - 1),
		26472 => to_unsigned(18599, LUT_AMPL_WIDTH - 1),
		26473 => to_unsigned(18597, LUT_AMPL_WIDTH - 1),
		26474 => to_unsigned(18594, LUT_AMPL_WIDTH - 1),
		26475 => to_unsigned(18592, LUT_AMPL_WIDTH - 1),
		26476 => to_unsigned(18589, LUT_AMPL_WIDTH - 1),
		26477 => to_unsigned(18587, LUT_AMPL_WIDTH - 1),
		26478 => to_unsigned(18584, LUT_AMPL_WIDTH - 1),
		26479 => to_unsigned(18581, LUT_AMPL_WIDTH - 1),
		26480 => to_unsigned(18579, LUT_AMPL_WIDTH - 1),
		26481 => to_unsigned(18576, LUT_AMPL_WIDTH - 1),
		26482 => to_unsigned(18574, LUT_AMPL_WIDTH - 1),
		26483 => to_unsigned(18571, LUT_AMPL_WIDTH - 1),
		26484 => to_unsigned(18568, LUT_AMPL_WIDTH - 1),
		26485 => to_unsigned(18566, LUT_AMPL_WIDTH - 1),
		26486 => to_unsigned(18563, LUT_AMPL_WIDTH - 1),
		26487 => to_unsigned(18561, LUT_AMPL_WIDTH - 1),
		26488 => to_unsigned(18558, LUT_AMPL_WIDTH - 1),
		26489 => to_unsigned(18555, LUT_AMPL_WIDTH - 1),
		26490 => to_unsigned(18553, LUT_AMPL_WIDTH - 1),
		26491 => to_unsigned(18550, LUT_AMPL_WIDTH - 1),
		26492 => to_unsigned(18548, LUT_AMPL_WIDTH - 1),
		26493 => to_unsigned(18545, LUT_AMPL_WIDTH - 1),
		26494 => to_unsigned(18543, LUT_AMPL_WIDTH - 1),
		26495 => to_unsigned(18540, LUT_AMPL_WIDTH - 1),
		26496 => to_unsigned(18537, LUT_AMPL_WIDTH - 1),
		26497 => to_unsigned(18535, LUT_AMPL_WIDTH - 1),
		26498 => to_unsigned(18532, LUT_AMPL_WIDTH - 1),
		26499 => to_unsigned(18530, LUT_AMPL_WIDTH - 1),
		26500 => to_unsigned(18527, LUT_AMPL_WIDTH - 1),
		26501 => to_unsigned(18524, LUT_AMPL_WIDTH - 1),
		26502 => to_unsigned(18522, LUT_AMPL_WIDTH - 1),
		26503 => to_unsigned(18519, LUT_AMPL_WIDTH - 1),
		26504 => to_unsigned(18517, LUT_AMPL_WIDTH - 1),
		26505 => to_unsigned(18514, LUT_AMPL_WIDTH - 1),
		26506 => to_unsigned(18511, LUT_AMPL_WIDTH - 1),
		26507 => to_unsigned(18509, LUT_AMPL_WIDTH - 1),
		26508 => to_unsigned(18506, LUT_AMPL_WIDTH - 1),
		26509 => to_unsigned(18504, LUT_AMPL_WIDTH - 1),
		26510 => to_unsigned(18501, LUT_AMPL_WIDTH - 1),
		26511 => to_unsigned(18498, LUT_AMPL_WIDTH - 1),
		26512 => to_unsigned(18496, LUT_AMPL_WIDTH - 1),
		26513 => to_unsigned(18493, LUT_AMPL_WIDTH - 1),
		26514 => to_unsigned(18491, LUT_AMPL_WIDTH - 1),
		26515 => to_unsigned(18488, LUT_AMPL_WIDTH - 1),
		26516 => to_unsigned(18485, LUT_AMPL_WIDTH - 1),
		26517 => to_unsigned(18483, LUT_AMPL_WIDTH - 1),
		26518 => to_unsigned(18480, LUT_AMPL_WIDTH - 1),
		26519 => to_unsigned(18478, LUT_AMPL_WIDTH - 1),
		26520 => to_unsigned(18475, LUT_AMPL_WIDTH - 1),
		26521 => to_unsigned(18473, LUT_AMPL_WIDTH - 1),
		26522 => to_unsigned(18470, LUT_AMPL_WIDTH - 1),
		26523 => to_unsigned(18467, LUT_AMPL_WIDTH - 1),
		26524 => to_unsigned(18465, LUT_AMPL_WIDTH - 1),
		26525 => to_unsigned(18462, LUT_AMPL_WIDTH - 1),
		26526 => to_unsigned(18460, LUT_AMPL_WIDTH - 1),
		26527 => to_unsigned(18457, LUT_AMPL_WIDTH - 1),
		26528 => to_unsigned(18454, LUT_AMPL_WIDTH - 1),
		26529 => to_unsigned(18452, LUT_AMPL_WIDTH - 1),
		26530 => to_unsigned(18449, LUT_AMPL_WIDTH - 1),
		26531 => to_unsigned(18447, LUT_AMPL_WIDTH - 1),
		26532 => to_unsigned(18444, LUT_AMPL_WIDTH - 1),
		26533 => to_unsigned(18441, LUT_AMPL_WIDTH - 1),
		26534 => to_unsigned(18439, LUT_AMPL_WIDTH - 1),
		26535 => to_unsigned(18436, LUT_AMPL_WIDTH - 1),
		26536 => to_unsigned(18434, LUT_AMPL_WIDTH - 1),
		26537 => to_unsigned(18431, LUT_AMPL_WIDTH - 1),
		26538 => to_unsigned(18428, LUT_AMPL_WIDTH - 1),
		26539 => to_unsigned(18426, LUT_AMPL_WIDTH - 1),
		26540 => to_unsigned(18423, LUT_AMPL_WIDTH - 1),
		26541 => to_unsigned(18421, LUT_AMPL_WIDTH - 1),
		26542 => to_unsigned(18418, LUT_AMPL_WIDTH - 1),
		26543 => to_unsigned(18415, LUT_AMPL_WIDTH - 1),
		26544 => to_unsigned(18413, LUT_AMPL_WIDTH - 1),
		26545 => to_unsigned(18410, LUT_AMPL_WIDTH - 1),
		26546 => to_unsigned(18408, LUT_AMPL_WIDTH - 1),
		26547 => to_unsigned(18405, LUT_AMPL_WIDTH - 1),
		26548 => to_unsigned(18402, LUT_AMPL_WIDTH - 1),
		26549 => to_unsigned(18400, LUT_AMPL_WIDTH - 1),
		26550 => to_unsigned(18397, LUT_AMPL_WIDTH - 1),
		26551 => to_unsigned(18395, LUT_AMPL_WIDTH - 1),
		26552 => to_unsigned(18392, LUT_AMPL_WIDTH - 1),
		26553 => to_unsigned(18389, LUT_AMPL_WIDTH - 1),
		26554 => to_unsigned(18387, LUT_AMPL_WIDTH - 1),
		26555 => to_unsigned(18384, LUT_AMPL_WIDTH - 1),
		26556 => to_unsigned(18382, LUT_AMPL_WIDTH - 1),
		26557 => to_unsigned(18379, LUT_AMPL_WIDTH - 1),
		26558 => to_unsigned(18376, LUT_AMPL_WIDTH - 1),
		26559 => to_unsigned(18374, LUT_AMPL_WIDTH - 1),
		26560 => to_unsigned(18371, LUT_AMPL_WIDTH - 1),
		26561 => to_unsigned(18369, LUT_AMPL_WIDTH - 1),
		26562 => to_unsigned(18366, LUT_AMPL_WIDTH - 1),
		26563 => to_unsigned(18363, LUT_AMPL_WIDTH - 1),
		26564 => to_unsigned(18361, LUT_AMPL_WIDTH - 1),
		26565 => to_unsigned(18358, LUT_AMPL_WIDTH - 1),
		26566 => to_unsigned(18356, LUT_AMPL_WIDTH - 1),
		26567 => to_unsigned(18353, LUT_AMPL_WIDTH - 1),
		26568 => to_unsigned(18350, LUT_AMPL_WIDTH - 1),
		26569 => to_unsigned(18348, LUT_AMPL_WIDTH - 1),
		26570 => to_unsigned(18345, LUT_AMPL_WIDTH - 1),
		26571 => to_unsigned(18343, LUT_AMPL_WIDTH - 1),
		26572 => to_unsigned(18340, LUT_AMPL_WIDTH - 1),
		26573 => to_unsigned(18337, LUT_AMPL_WIDTH - 1),
		26574 => to_unsigned(18335, LUT_AMPL_WIDTH - 1),
		26575 => to_unsigned(18332, LUT_AMPL_WIDTH - 1),
		26576 => to_unsigned(18330, LUT_AMPL_WIDTH - 1),
		26577 => to_unsigned(18327, LUT_AMPL_WIDTH - 1),
		26578 => to_unsigned(18324, LUT_AMPL_WIDTH - 1),
		26579 => to_unsigned(18322, LUT_AMPL_WIDTH - 1),
		26580 => to_unsigned(18319, LUT_AMPL_WIDTH - 1),
		26581 => to_unsigned(18317, LUT_AMPL_WIDTH - 1),
		26582 => to_unsigned(18314, LUT_AMPL_WIDTH - 1),
		26583 => to_unsigned(18311, LUT_AMPL_WIDTH - 1),
		26584 => to_unsigned(18309, LUT_AMPL_WIDTH - 1),
		26585 => to_unsigned(18306, LUT_AMPL_WIDTH - 1),
		26586 => to_unsigned(18304, LUT_AMPL_WIDTH - 1),
		26587 => to_unsigned(18301, LUT_AMPL_WIDTH - 1),
		26588 => to_unsigned(18298, LUT_AMPL_WIDTH - 1),
		26589 => to_unsigned(18296, LUT_AMPL_WIDTH - 1),
		26590 => to_unsigned(18293, LUT_AMPL_WIDTH - 1),
		26591 => to_unsigned(18290, LUT_AMPL_WIDTH - 1),
		26592 => to_unsigned(18288, LUT_AMPL_WIDTH - 1),
		26593 => to_unsigned(18285, LUT_AMPL_WIDTH - 1),
		26594 => to_unsigned(18283, LUT_AMPL_WIDTH - 1),
		26595 => to_unsigned(18280, LUT_AMPL_WIDTH - 1),
		26596 => to_unsigned(18277, LUT_AMPL_WIDTH - 1),
		26597 => to_unsigned(18275, LUT_AMPL_WIDTH - 1),
		26598 => to_unsigned(18272, LUT_AMPL_WIDTH - 1),
		26599 => to_unsigned(18270, LUT_AMPL_WIDTH - 1),
		26600 => to_unsigned(18267, LUT_AMPL_WIDTH - 1),
		26601 => to_unsigned(18264, LUT_AMPL_WIDTH - 1),
		26602 => to_unsigned(18262, LUT_AMPL_WIDTH - 1),
		26603 => to_unsigned(18259, LUT_AMPL_WIDTH - 1),
		26604 => to_unsigned(18257, LUT_AMPL_WIDTH - 1),
		26605 => to_unsigned(18254, LUT_AMPL_WIDTH - 1),
		26606 => to_unsigned(18251, LUT_AMPL_WIDTH - 1),
		26607 => to_unsigned(18249, LUT_AMPL_WIDTH - 1),
		26608 => to_unsigned(18246, LUT_AMPL_WIDTH - 1),
		26609 => to_unsigned(18244, LUT_AMPL_WIDTH - 1),
		26610 => to_unsigned(18241, LUT_AMPL_WIDTH - 1),
		26611 => to_unsigned(18238, LUT_AMPL_WIDTH - 1),
		26612 => to_unsigned(18236, LUT_AMPL_WIDTH - 1),
		26613 => to_unsigned(18233, LUT_AMPL_WIDTH - 1),
		26614 => to_unsigned(18230, LUT_AMPL_WIDTH - 1),
		26615 => to_unsigned(18228, LUT_AMPL_WIDTH - 1),
		26616 => to_unsigned(18225, LUT_AMPL_WIDTH - 1),
		26617 => to_unsigned(18223, LUT_AMPL_WIDTH - 1),
		26618 => to_unsigned(18220, LUT_AMPL_WIDTH - 1),
		26619 => to_unsigned(18217, LUT_AMPL_WIDTH - 1),
		26620 => to_unsigned(18215, LUT_AMPL_WIDTH - 1),
		26621 => to_unsigned(18212, LUT_AMPL_WIDTH - 1),
		26622 => to_unsigned(18210, LUT_AMPL_WIDTH - 1),
		26623 => to_unsigned(18207, LUT_AMPL_WIDTH - 1),
		26624 => to_unsigned(18204, LUT_AMPL_WIDTH - 1),
		26625 => to_unsigned(18202, LUT_AMPL_WIDTH - 1),
		26626 => to_unsigned(18199, LUT_AMPL_WIDTH - 1),
		26627 => to_unsigned(18197, LUT_AMPL_WIDTH - 1),
		26628 => to_unsigned(18194, LUT_AMPL_WIDTH - 1),
		26629 => to_unsigned(18191, LUT_AMPL_WIDTH - 1),
		26630 => to_unsigned(18189, LUT_AMPL_WIDTH - 1),
		26631 => to_unsigned(18186, LUT_AMPL_WIDTH - 1),
		26632 => to_unsigned(18183, LUT_AMPL_WIDTH - 1),
		26633 => to_unsigned(18181, LUT_AMPL_WIDTH - 1),
		26634 => to_unsigned(18178, LUT_AMPL_WIDTH - 1),
		26635 => to_unsigned(18176, LUT_AMPL_WIDTH - 1),
		26636 => to_unsigned(18173, LUT_AMPL_WIDTH - 1),
		26637 => to_unsigned(18170, LUT_AMPL_WIDTH - 1),
		26638 => to_unsigned(18168, LUT_AMPL_WIDTH - 1),
		26639 => to_unsigned(18165, LUT_AMPL_WIDTH - 1),
		26640 => to_unsigned(18163, LUT_AMPL_WIDTH - 1),
		26641 => to_unsigned(18160, LUT_AMPL_WIDTH - 1),
		26642 => to_unsigned(18157, LUT_AMPL_WIDTH - 1),
		26643 => to_unsigned(18155, LUT_AMPL_WIDTH - 1),
		26644 => to_unsigned(18152, LUT_AMPL_WIDTH - 1),
		26645 => to_unsigned(18149, LUT_AMPL_WIDTH - 1),
		26646 => to_unsigned(18147, LUT_AMPL_WIDTH - 1),
		26647 => to_unsigned(18144, LUT_AMPL_WIDTH - 1),
		26648 => to_unsigned(18142, LUT_AMPL_WIDTH - 1),
		26649 => to_unsigned(18139, LUT_AMPL_WIDTH - 1),
		26650 => to_unsigned(18136, LUT_AMPL_WIDTH - 1),
		26651 => to_unsigned(18134, LUT_AMPL_WIDTH - 1),
		26652 => to_unsigned(18131, LUT_AMPL_WIDTH - 1),
		26653 => to_unsigned(18129, LUT_AMPL_WIDTH - 1),
		26654 => to_unsigned(18126, LUT_AMPL_WIDTH - 1),
		26655 => to_unsigned(18123, LUT_AMPL_WIDTH - 1),
		26656 => to_unsigned(18121, LUT_AMPL_WIDTH - 1),
		26657 => to_unsigned(18118, LUT_AMPL_WIDTH - 1),
		26658 => to_unsigned(18115, LUT_AMPL_WIDTH - 1),
		26659 => to_unsigned(18113, LUT_AMPL_WIDTH - 1),
		26660 => to_unsigned(18110, LUT_AMPL_WIDTH - 1),
		26661 => to_unsigned(18108, LUT_AMPL_WIDTH - 1),
		26662 => to_unsigned(18105, LUT_AMPL_WIDTH - 1),
		26663 => to_unsigned(18102, LUT_AMPL_WIDTH - 1),
		26664 => to_unsigned(18100, LUT_AMPL_WIDTH - 1),
		26665 => to_unsigned(18097, LUT_AMPL_WIDTH - 1),
		26666 => to_unsigned(18095, LUT_AMPL_WIDTH - 1),
		26667 => to_unsigned(18092, LUT_AMPL_WIDTH - 1),
		26668 => to_unsigned(18089, LUT_AMPL_WIDTH - 1),
		26669 => to_unsigned(18087, LUT_AMPL_WIDTH - 1),
		26670 => to_unsigned(18084, LUT_AMPL_WIDTH - 1),
		26671 => to_unsigned(18081, LUT_AMPL_WIDTH - 1),
		26672 => to_unsigned(18079, LUT_AMPL_WIDTH - 1),
		26673 => to_unsigned(18076, LUT_AMPL_WIDTH - 1),
		26674 => to_unsigned(18074, LUT_AMPL_WIDTH - 1),
		26675 => to_unsigned(18071, LUT_AMPL_WIDTH - 1),
		26676 => to_unsigned(18068, LUT_AMPL_WIDTH - 1),
		26677 => to_unsigned(18066, LUT_AMPL_WIDTH - 1),
		26678 => to_unsigned(18063, LUT_AMPL_WIDTH - 1),
		26679 => to_unsigned(18060, LUT_AMPL_WIDTH - 1),
		26680 => to_unsigned(18058, LUT_AMPL_WIDTH - 1),
		26681 => to_unsigned(18055, LUT_AMPL_WIDTH - 1),
		26682 => to_unsigned(18053, LUT_AMPL_WIDTH - 1),
		26683 => to_unsigned(18050, LUT_AMPL_WIDTH - 1),
		26684 => to_unsigned(18047, LUT_AMPL_WIDTH - 1),
		26685 => to_unsigned(18045, LUT_AMPL_WIDTH - 1),
		26686 => to_unsigned(18042, LUT_AMPL_WIDTH - 1),
		26687 => to_unsigned(18039, LUT_AMPL_WIDTH - 1),
		26688 => to_unsigned(18037, LUT_AMPL_WIDTH - 1),
		26689 => to_unsigned(18034, LUT_AMPL_WIDTH - 1),
		26690 => to_unsigned(18032, LUT_AMPL_WIDTH - 1),
		26691 => to_unsigned(18029, LUT_AMPL_WIDTH - 1),
		26692 => to_unsigned(18026, LUT_AMPL_WIDTH - 1),
		26693 => to_unsigned(18024, LUT_AMPL_WIDTH - 1),
		26694 => to_unsigned(18021, LUT_AMPL_WIDTH - 1),
		26695 => to_unsigned(18018, LUT_AMPL_WIDTH - 1),
		26696 => to_unsigned(18016, LUT_AMPL_WIDTH - 1),
		26697 => to_unsigned(18013, LUT_AMPL_WIDTH - 1),
		26698 => to_unsigned(18011, LUT_AMPL_WIDTH - 1),
		26699 => to_unsigned(18008, LUT_AMPL_WIDTH - 1),
		26700 => to_unsigned(18005, LUT_AMPL_WIDTH - 1),
		26701 => to_unsigned(18003, LUT_AMPL_WIDTH - 1),
		26702 => to_unsigned(18000, LUT_AMPL_WIDTH - 1),
		26703 => to_unsigned(17997, LUT_AMPL_WIDTH - 1),
		26704 => to_unsigned(17995, LUT_AMPL_WIDTH - 1),
		26705 => to_unsigned(17992, LUT_AMPL_WIDTH - 1),
		26706 => to_unsigned(17990, LUT_AMPL_WIDTH - 1),
		26707 => to_unsigned(17987, LUT_AMPL_WIDTH - 1),
		26708 => to_unsigned(17984, LUT_AMPL_WIDTH - 1),
		26709 => to_unsigned(17982, LUT_AMPL_WIDTH - 1),
		26710 => to_unsigned(17979, LUT_AMPL_WIDTH - 1),
		26711 => to_unsigned(17976, LUT_AMPL_WIDTH - 1),
		26712 => to_unsigned(17974, LUT_AMPL_WIDTH - 1),
		26713 => to_unsigned(17971, LUT_AMPL_WIDTH - 1),
		26714 => to_unsigned(17969, LUT_AMPL_WIDTH - 1),
		26715 => to_unsigned(17966, LUT_AMPL_WIDTH - 1),
		26716 => to_unsigned(17963, LUT_AMPL_WIDTH - 1),
		26717 => to_unsigned(17961, LUT_AMPL_WIDTH - 1),
		26718 => to_unsigned(17958, LUT_AMPL_WIDTH - 1),
		26719 => to_unsigned(17955, LUT_AMPL_WIDTH - 1),
		26720 => to_unsigned(17953, LUT_AMPL_WIDTH - 1),
		26721 => to_unsigned(17950, LUT_AMPL_WIDTH - 1),
		26722 => to_unsigned(17948, LUT_AMPL_WIDTH - 1),
		26723 => to_unsigned(17945, LUT_AMPL_WIDTH - 1),
		26724 => to_unsigned(17942, LUT_AMPL_WIDTH - 1),
		26725 => to_unsigned(17940, LUT_AMPL_WIDTH - 1),
		26726 => to_unsigned(17937, LUT_AMPL_WIDTH - 1),
		26727 => to_unsigned(17934, LUT_AMPL_WIDTH - 1),
		26728 => to_unsigned(17932, LUT_AMPL_WIDTH - 1),
		26729 => to_unsigned(17929, LUT_AMPL_WIDTH - 1),
		26730 => to_unsigned(17927, LUT_AMPL_WIDTH - 1),
		26731 => to_unsigned(17924, LUT_AMPL_WIDTH - 1),
		26732 => to_unsigned(17921, LUT_AMPL_WIDTH - 1),
		26733 => to_unsigned(17919, LUT_AMPL_WIDTH - 1),
		26734 => to_unsigned(17916, LUT_AMPL_WIDTH - 1),
		26735 => to_unsigned(17913, LUT_AMPL_WIDTH - 1),
		26736 => to_unsigned(17911, LUT_AMPL_WIDTH - 1),
		26737 => to_unsigned(17908, LUT_AMPL_WIDTH - 1),
		26738 => to_unsigned(17906, LUT_AMPL_WIDTH - 1),
		26739 => to_unsigned(17903, LUT_AMPL_WIDTH - 1),
		26740 => to_unsigned(17900, LUT_AMPL_WIDTH - 1),
		26741 => to_unsigned(17898, LUT_AMPL_WIDTH - 1),
		26742 => to_unsigned(17895, LUT_AMPL_WIDTH - 1),
		26743 => to_unsigned(17892, LUT_AMPL_WIDTH - 1),
		26744 => to_unsigned(17890, LUT_AMPL_WIDTH - 1),
		26745 => to_unsigned(17887, LUT_AMPL_WIDTH - 1),
		26746 => to_unsigned(17884, LUT_AMPL_WIDTH - 1),
		26747 => to_unsigned(17882, LUT_AMPL_WIDTH - 1),
		26748 => to_unsigned(17879, LUT_AMPL_WIDTH - 1),
		26749 => to_unsigned(17877, LUT_AMPL_WIDTH - 1),
		26750 => to_unsigned(17874, LUT_AMPL_WIDTH - 1),
		26751 => to_unsigned(17871, LUT_AMPL_WIDTH - 1),
		26752 => to_unsigned(17869, LUT_AMPL_WIDTH - 1),
		26753 => to_unsigned(17866, LUT_AMPL_WIDTH - 1),
		26754 => to_unsigned(17863, LUT_AMPL_WIDTH - 1),
		26755 => to_unsigned(17861, LUT_AMPL_WIDTH - 1),
		26756 => to_unsigned(17858, LUT_AMPL_WIDTH - 1),
		26757 => to_unsigned(17855, LUT_AMPL_WIDTH - 1),
		26758 => to_unsigned(17853, LUT_AMPL_WIDTH - 1),
		26759 => to_unsigned(17850, LUT_AMPL_WIDTH - 1),
		26760 => to_unsigned(17848, LUT_AMPL_WIDTH - 1),
		26761 => to_unsigned(17845, LUT_AMPL_WIDTH - 1),
		26762 => to_unsigned(17842, LUT_AMPL_WIDTH - 1),
		26763 => to_unsigned(17840, LUT_AMPL_WIDTH - 1),
		26764 => to_unsigned(17837, LUT_AMPL_WIDTH - 1),
		26765 => to_unsigned(17834, LUT_AMPL_WIDTH - 1),
		26766 => to_unsigned(17832, LUT_AMPL_WIDTH - 1),
		26767 => to_unsigned(17829, LUT_AMPL_WIDTH - 1),
		26768 => to_unsigned(17827, LUT_AMPL_WIDTH - 1),
		26769 => to_unsigned(17824, LUT_AMPL_WIDTH - 1),
		26770 => to_unsigned(17821, LUT_AMPL_WIDTH - 1),
		26771 => to_unsigned(17819, LUT_AMPL_WIDTH - 1),
		26772 => to_unsigned(17816, LUT_AMPL_WIDTH - 1),
		26773 => to_unsigned(17813, LUT_AMPL_WIDTH - 1),
		26774 => to_unsigned(17811, LUT_AMPL_WIDTH - 1),
		26775 => to_unsigned(17808, LUT_AMPL_WIDTH - 1),
		26776 => to_unsigned(17805, LUT_AMPL_WIDTH - 1),
		26777 => to_unsigned(17803, LUT_AMPL_WIDTH - 1),
		26778 => to_unsigned(17800, LUT_AMPL_WIDTH - 1),
		26779 => to_unsigned(17798, LUT_AMPL_WIDTH - 1),
		26780 => to_unsigned(17795, LUT_AMPL_WIDTH - 1),
		26781 => to_unsigned(17792, LUT_AMPL_WIDTH - 1),
		26782 => to_unsigned(17790, LUT_AMPL_WIDTH - 1),
		26783 => to_unsigned(17787, LUT_AMPL_WIDTH - 1),
		26784 => to_unsigned(17784, LUT_AMPL_WIDTH - 1),
		26785 => to_unsigned(17782, LUT_AMPL_WIDTH - 1),
		26786 => to_unsigned(17779, LUT_AMPL_WIDTH - 1),
		26787 => to_unsigned(17776, LUT_AMPL_WIDTH - 1),
		26788 => to_unsigned(17774, LUT_AMPL_WIDTH - 1),
		26789 => to_unsigned(17771, LUT_AMPL_WIDTH - 1),
		26790 => to_unsigned(17768, LUT_AMPL_WIDTH - 1),
		26791 => to_unsigned(17766, LUT_AMPL_WIDTH - 1),
		26792 => to_unsigned(17763, LUT_AMPL_WIDTH - 1),
		26793 => to_unsigned(17761, LUT_AMPL_WIDTH - 1),
		26794 => to_unsigned(17758, LUT_AMPL_WIDTH - 1),
		26795 => to_unsigned(17755, LUT_AMPL_WIDTH - 1),
		26796 => to_unsigned(17753, LUT_AMPL_WIDTH - 1),
		26797 => to_unsigned(17750, LUT_AMPL_WIDTH - 1),
		26798 => to_unsigned(17747, LUT_AMPL_WIDTH - 1),
		26799 => to_unsigned(17745, LUT_AMPL_WIDTH - 1),
		26800 => to_unsigned(17742, LUT_AMPL_WIDTH - 1),
		26801 => to_unsigned(17739, LUT_AMPL_WIDTH - 1),
		26802 => to_unsigned(17737, LUT_AMPL_WIDTH - 1),
		26803 => to_unsigned(17734, LUT_AMPL_WIDTH - 1),
		26804 => to_unsigned(17732, LUT_AMPL_WIDTH - 1),
		26805 => to_unsigned(17729, LUT_AMPL_WIDTH - 1),
		26806 => to_unsigned(17726, LUT_AMPL_WIDTH - 1),
		26807 => to_unsigned(17724, LUT_AMPL_WIDTH - 1),
		26808 => to_unsigned(17721, LUT_AMPL_WIDTH - 1),
		26809 => to_unsigned(17718, LUT_AMPL_WIDTH - 1),
		26810 => to_unsigned(17716, LUT_AMPL_WIDTH - 1),
		26811 => to_unsigned(17713, LUT_AMPL_WIDTH - 1),
		26812 => to_unsigned(17710, LUT_AMPL_WIDTH - 1),
		26813 => to_unsigned(17708, LUT_AMPL_WIDTH - 1),
		26814 => to_unsigned(17705, LUT_AMPL_WIDTH - 1),
		26815 => to_unsigned(17702, LUT_AMPL_WIDTH - 1),
		26816 => to_unsigned(17700, LUT_AMPL_WIDTH - 1),
		26817 => to_unsigned(17697, LUT_AMPL_WIDTH - 1),
		26818 => to_unsigned(17695, LUT_AMPL_WIDTH - 1),
		26819 => to_unsigned(17692, LUT_AMPL_WIDTH - 1),
		26820 => to_unsigned(17689, LUT_AMPL_WIDTH - 1),
		26821 => to_unsigned(17687, LUT_AMPL_WIDTH - 1),
		26822 => to_unsigned(17684, LUT_AMPL_WIDTH - 1),
		26823 => to_unsigned(17681, LUT_AMPL_WIDTH - 1),
		26824 => to_unsigned(17679, LUT_AMPL_WIDTH - 1),
		26825 => to_unsigned(17676, LUT_AMPL_WIDTH - 1),
		26826 => to_unsigned(17673, LUT_AMPL_WIDTH - 1),
		26827 => to_unsigned(17671, LUT_AMPL_WIDTH - 1),
		26828 => to_unsigned(17668, LUT_AMPL_WIDTH - 1),
		26829 => to_unsigned(17665, LUT_AMPL_WIDTH - 1),
		26830 => to_unsigned(17663, LUT_AMPL_WIDTH - 1),
		26831 => to_unsigned(17660, LUT_AMPL_WIDTH - 1),
		26832 => to_unsigned(17657, LUT_AMPL_WIDTH - 1),
		26833 => to_unsigned(17655, LUT_AMPL_WIDTH - 1),
		26834 => to_unsigned(17652, LUT_AMPL_WIDTH - 1),
		26835 => to_unsigned(17650, LUT_AMPL_WIDTH - 1),
		26836 => to_unsigned(17647, LUT_AMPL_WIDTH - 1),
		26837 => to_unsigned(17644, LUT_AMPL_WIDTH - 1),
		26838 => to_unsigned(17642, LUT_AMPL_WIDTH - 1),
		26839 => to_unsigned(17639, LUT_AMPL_WIDTH - 1),
		26840 => to_unsigned(17636, LUT_AMPL_WIDTH - 1),
		26841 => to_unsigned(17634, LUT_AMPL_WIDTH - 1),
		26842 => to_unsigned(17631, LUT_AMPL_WIDTH - 1),
		26843 => to_unsigned(17628, LUT_AMPL_WIDTH - 1),
		26844 => to_unsigned(17626, LUT_AMPL_WIDTH - 1),
		26845 => to_unsigned(17623, LUT_AMPL_WIDTH - 1),
		26846 => to_unsigned(17620, LUT_AMPL_WIDTH - 1),
		26847 => to_unsigned(17618, LUT_AMPL_WIDTH - 1),
		26848 => to_unsigned(17615, LUT_AMPL_WIDTH - 1),
		26849 => to_unsigned(17612, LUT_AMPL_WIDTH - 1),
		26850 => to_unsigned(17610, LUT_AMPL_WIDTH - 1),
		26851 => to_unsigned(17607, LUT_AMPL_WIDTH - 1),
		26852 => to_unsigned(17605, LUT_AMPL_WIDTH - 1),
		26853 => to_unsigned(17602, LUT_AMPL_WIDTH - 1),
		26854 => to_unsigned(17599, LUT_AMPL_WIDTH - 1),
		26855 => to_unsigned(17597, LUT_AMPL_WIDTH - 1),
		26856 => to_unsigned(17594, LUT_AMPL_WIDTH - 1),
		26857 => to_unsigned(17591, LUT_AMPL_WIDTH - 1),
		26858 => to_unsigned(17589, LUT_AMPL_WIDTH - 1),
		26859 => to_unsigned(17586, LUT_AMPL_WIDTH - 1),
		26860 => to_unsigned(17583, LUT_AMPL_WIDTH - 1),
		26861 => to_unsigned(17581, LUT_AMPL_WIDTH - 1),
		26862 => to_unsigned(17578, LUT_AMPL_WIDTH - 1),
		26863 => to_unsigned(17575, LUT_AMPL_WIDTH - 1),
		26864 => to_unsigned(17573, LUT_AMPL_WIDTH - 1),
		26865 => to_unsigned(17570, LUT_AMPL_WIDTH - 1),
		26866 => to_unsigned(17567, LUT_AMPL_WIDTH - 1),
		26867 => to_unsigned(17565, LUT_AMPL_WIDTH - 1),
		26868 => to_unsigned(17562, LUT_AMPL_WIDTH - 1),
		26869 => to_unsigned(17559, LUT_AMPL_WIDTH - 1),
		26870 => to_unsigned(17557, LUT_AMPL_WIDTH - 1),
		26871 => to_unsigned(17554, LUT_AMPL_WIDTH - 1),
		26872 => to_unsigned(17551, LUT_AMPL_WIDTH - 1),
		26873 => to_unsigned(17549, LUT_AMPL_WIDTH - 1),
		26874 => to_unsigned(17546, LUT_AMPL_WIDTH - 1),
		26875 => to_unsigned(17544, LUT_AMPL_WIDTH - 1),
		26876 => to_unsigned(17541, LUT_AMPL_WIDTH - 1),
		26877 => to_unsigned(17538, LUT_AMPL_WIDTH - 1),
		26878 => to_unsigned(17536, LUT_AMPL_WIDTH - 1),
		26879 => to_unsigned(17533, LUT_AMPL_WIDTH - 1),
		26880 => to_unsigned(17530, LUT_AMPL_WIDTH - 1),
		26881 => to_unsigned(17528, LUT_AMPL_WIDTH - 1),
		26882 => to_unsigned(17525, LUT_AMPL_WIDTH - 1),
		26883 => to_unsigned(17522, LUT_AMPL_WIDTH - 1),
		26884 => to_unsigned(17520, LUT_AMPL_WIDTH - 1),
		26885 => to_unsigned(17517, LUT_AMPL_WIDTH - 1),
		26886 => to_unsigned(17514, LUT_AMPL_WIDTH - 1),
		26887 => to_unsigned(17512, LUT_AMPL_WIDTH - 1),
		26888 => to_unsigned(17509, LUT_AMPL_WIDTH - 1),
		26889 => to_unsigned(17506, LUT_AMPL_WIDTH - 1),
		26890 => to_unsigned(17504, LUT_AMPL_WIDTH - 1),
		26891 => to_unsigned(17501, LUT_AMPL_WIDTH - 1),
		26892 => to_unsigned(17498, LUT_AMPL_WIDTH - 1),
		26893 => to_unsigned(17496, LUT_AMPL_WIDTH - 1),
		26894 => to_unsigned(17493, LUT_AMPL_WIDTH - 1),
		26895 => to_unsigned(17490, LUT_AMPL_WIDTH - 1),
		26896 => to_unsigned(17488, LUT_AMPL_WIDTH - 1),
		26897 => to_unsigned(17485, LUT_AMPL_WIDTH - 1),
		26898 => to_unsigned(17482, LUT_AMPL_WIDTH - 1),
		26899 => to_unsigned(17480, LUT_AMPL_WIDTH - 1),
		26900 => to_unsigned(17477, LUT_AMPL_WIDTH - 1),
		26901 => to_unsigned(17474, LUT_AMPL_WIDTH - 1),
		26902 => to_unsigned(17472, LUT_AMPL_WIDTH - 1),
		26903 => to_unsigned(17469, LUT_AMPL_WIDTH - 1),
		26904 => to_unsigned(17467, LUT_AMPL_WIDTH - 1),
		26905 => to_unsigned(17464, LUT_AMPL_WIDTH - 1),
		26906 => to_unsigned(17461, LUT_AMPL_WIDTH - 1),
		26907 => to_unsigned(17459, LUT_AMPL_WIDTH - 1),
		26908 => to_unsigned(17456, LUT_AMPL_WIDTH - 1),
		26909 => to_unsigned(17453, LUT_AMPL_WIDTH - 1),
		26910 => to_unsigned(17451, LUT_AMPL_WIDTH - 1),
		26911 => to_unsigned(17448, LUT_AMPL_WIDTH - 1),
		26912 => to_unsigned(17445, LUT_AMPL_WIDTH - 1),
		26913 => to_unsigned(17443, LUT_AMPL_WIDTH - 1),
		26914 => to_unsigned(17440, LUT_AMPL_WIDTH - 1),
		26915 => to_unsigned(17437, LUT_AMPL_WIDTH - 1),
		26916 => to_unsigned(17435, LUT_AMPL_WIDTH - 1),
		26917 => to_unsigned(17432, LUT_AMPL_WIDTH - 1),
		26918 => to_unsigned(17429, LUT_AMPL_WIDTH - 1),
		26919 => to_unsigned(17427, LUT_AMPL_WIDTH - 1),
		26920 => to_unsigned(17424, LUT_AMPL_WIDTH - 1),
		26921 => to_unsigned(17421, LUT_AMPL_WIDTH - 1),
		26922 => to_unsigned(17419, LUT_AMPL_WIDTH - 1),
		26923 => to_unsigned(17416, LUT_AMPL_WIDTH - 1),
		26924 => to_unsigned(17413, LUT_AMPL_WIDTH - 1),
		26925 => to_unsigned(17411, LUT_AMPL_WIDTH - 1),
		26926 => to_unsigned(17408, LUT_AMPL_WIDTH - 1),
		26927 => to_unsigned(17405, LUT_AMPL_WIDTH - 1),
		26928 => to_unsigned(17403, LUT_AMPL_WIDTH - 1),
		26929 => to_unsigned(17400, LUT_AMPL_WIDTH - 1),
		26930 => to_unsigned(17397, LUT_AMPL_WIDTH - 1),
		26931 => to_unsigned(17395, LUT_AMPL_WIDTH - 1),
		26932 => to_unsigned(17392, LUT_AMPL_WIDTH - 1),
		26933 => to_unsigned(17389, LUT_AMPL_WIDTH - 1),
		26934 => to_unsigned(17387, LUT_AMPL_WIDTH - 1),
		26935 => to_unsigned(17384, LUT_AMPL_WIDTH - 1),
		26936 => to_unsigned(17381, LUT_AMPL_WIDTH - 1),
		26937 => to_unsigned(17379, LUT_AMPL_WIDTH - 1),
		26938 => to_unsigned(17376, LUT_AMPL_WIDTH - 1),
		26939 => to_unsigned(17373, LUT_AMPL_WIDTH - 1),
		26940 => to_unsigned(17371, LUT_AMPL_WIDTH - 1),
		26941 => to_unsigned(17368, LUT_AMPL_WIDTH - 1),
		26942 => to_unsigned(17365, LUT_AMPL_WIDTH - 1),
		26943 => to_unsigned(17363, LUT_AMPL_WIDTH - 1),
		26944 => to_unsigned(17360, LUT_AMPL_WIDTH - 1),
		26945 => to_unsigned(17357, LUT_AMPL_WIDTH - 1),
		26946 => to_unsigned(17355, LUT_AMPL_WIDTH - 1),
		26947 => to_unsigned(17352, LUT_AMPL_WIDTH - 1),
		26948 => to_unsigned(17349, LUT_AMPL_WIDTH - 1),
		26949 => to_unsigned(17347, LUT_AMPL_WIDTH - 1),
		26950 => to_unsigned(17344, LUT_AMPL_WIDTH - 1),
		26951 => to_unsigned(17341, LUT_AMPL_WIDTH - 1),
		26952 => to_unsigned(17339, LUT_AMPL_WIDTH - 1),
		26953 => to_unsigned(17336, LUT_AMPL_WIDTH - 1),
		26954 => to_unsigned(17333, LUT_AMPL_WIDTH - 1),
		26955 => to_unsigned(17331, LUT_AMPL_WIDTH - 1),
		26956 => to_unsigned(17328, LUT_AMPL_WIDTH - 1),
		26957 => to_unsigned(17325, LUT_AMPL_WIDTH - 1),
		26958 => to_unsigned(17323, LUT_AMPL_WIDTH - 1),
		26959 => to_unsigned(17320, LUT_AMPL_WIDTH - 1),
		26960 => to_unsigned(17317, LUT_AMPL_WIDTH - 1),
		26961 => to_unsigned(17315, LUT_AMPL_WIDTH - 1),
		26962 => to_unsigned(17312, LUT_AMPL_WIDTH - 1),
		26963 => to_unsigned(17309, LUT_AMPL_WIDTH - 1),
		26964 => to_unsigned(17307, LUT_AMPL_WIDTH - 1),
		26965 => to_unsigned(17304, LUT_AMPL_WIDTH - 1),
		26966 => to_unsigned(17301, LUT_AMPL_WIDTH - 1),
		26967 => to_unsigned(17299, LUT_AMPL_WIDTH - 1),
		26968 => to_unsigned(17296, LUT_AMPL_WIDTH - 1),
		26969 => to_unsigned(17293, LUT_AMPL_WIDTH - 1),
		26970 => to_unsigned(17291, LUT_AMPL_WIDTH - 1),
		26971 => to_unsigned(17288, LUT_AMPL_WIDTH - 1),
		26972 => to_unsigned(17285, LUT_AMPL_WIDTH - 1),
		26973 => to_unsigned(17283, LUT_AMPL_WIDTH - 1),
		26974 => to_unsigned(17280, LUT_AMPL_WIDTH - 1),
		26975 => to_unsigned(17277, LUT_AMPL_WIDTH - 1),
		26976 => to_unsigned(17275, LUT_AMPL_WIDTH - 1),
		26977 => to_unsigned(17272, LUT_AMPL_WIDTH - 1),
		26978 => to_unsigned(17269, LUT_AMPL_WIDTH - 1),
		26979 => to_unsigned(17267, LUT_AMPL_WIDTH - 1),
		26980 => to_unsigned(17264, LUT_AMPL_WIDTH - 1),
		26981 => to_unsigned(17261, LUT_AMPL_WIDTH - 1),
		26982 => to_unsigned(17259, LUT_AMPL_WIDTH - 1),
		26983 => to_unsigned(17256, LUT_AMPL_WIDTH - 1),
		26984 => to_unsigned(17253, LUT_AMPL_WIDTH - 1),
		26985 => to_unsigned(17251, LUT_AMPL_WIDTH - 1),
		26986 => to_unsigned(17248, LUT_AMPL_WIDTH - 1),
		26987 => to_unsigned(17245, LUT_AMPL_WIDTH - 1),
		26988 => to_unsigned(17243, LUT_AMPL_WIDTH - 1),
		26989 => to_unsigned(17240, LUT_AMPL_WIDTH - 1),
		26990 => to_unsigned(17237, LUT_AMPL_WIDTH - 1),
		26991 => to_unsigned(17235, LUT_AMPL_WIDTH - 1),
		26992 => to_unsigned(17232, LUT_AMPL_WIDTH - 1),
		26993 => to_unsigned(17229, LUT_AMPL_WIDTH - 1),
		26994 => to_unsigned(17227, LUT_AMPL_WIDTH - 1),
		26995 => to_unsigned(17224, LUT_AMPL_WIDTH - 1),
		26996 => to_unsigned(17221, LUT_AMPL_WIDTH - 1),
		26997 => to_unsigned(17219, LUT_AMPL_WIDTH - 1),
		26998 => to_unsigned(17216, LUT_AMPL_WIDTH - 1),
		26999 => to_unsigned(17213, LUT_AMPL_WIDTH - 1),
		27000 => to_unsigned(17211, LUT_AMPL_WIDTH - 1),
		27001 => to_unsigned(17208, LUT_AMPL_WIDTH - 1),
		27002 => to_unsigned(17205, LUT_AMPL_WIDTH - 1),
		27003 => to_unsigned(17203, LUT_AMPL_WIDTH - 1),
		27004 => to_unsigned(17200, LUT_AMPL_WIDTH - 1),
		27005 => to_unsigned(17197, LUT_AMPL_WIDTH - 1),
		27006 => to_unsigned(17195, LUT_AMPL_WIDTH - 1),
		27007 => to_unsigned(17192, LUT_AMPL_WIDTH - 1),
		27008 => to_unsigned(17189, LUT_AMPL_WIDTH - 1),
		27009 => to_unsigned(17187, LUT_AMPL_WIDTH - 1),
		27010 => to_unsigned(17184, LUT_AMPL_WIDTH - 1),
		27011 => to_unsigned(17181, LUT_AMPL_WIDTH - 1),
		27012 => to_unsigned(17179, LUT_AMPL_WIDTH - 1),
		27013 => to_unsigned(17176, LUT_AMPL_WIDTH - 1),
		27014 => to_unsigned(17173, LUT_AMPL_WIDTH - 1),
		27015 => to_unsigned(17171, LUT_AMPL_WIDTH - 1),
		27016 => to_unsigned(17168, LUT_AMPL_WIDTH - 1),
		27017 => to_unsigned(17165, LUT_AMPL_WIDTH - 1),
		27018 => to_unsigned(17162, LUT_AMPL_WIDTH - 1),
		27019 => to_unsigned(17160, LUT_AMPL_WIDTH - 1),
		27020 => to_unsigned(17157, LUT_AMPL_WIDTH - 1),
		27021 => to_unsigned(17154, LUT_AMPL_WIDTH - 1),
		27022 => to_unsigned(17152, LUT_AMPL_WIDTH - 1),
		27023 => to_unsigned(17149, LUT_AMPL_WIDTH - 1),
		27024 => to_unsigned(17146, LUT_AMPL_WIDTH - 1),
		27025 => to_unsigned(17144, LUT_AMPL_WIDTH - 1),
		27026 => to_unsigned(17141, LUT_AMPL_WIDTH - 1),
		27027 => to_unsigned(17138, LUT_AMPL_WIDTH - 1),
		27028 => to_unsigned(17136, LUT_AMPL_WIDTH - 1),
		27029 => to_unsigned(17133, LUT_AMPL_WIDTH - 1),
		27030 => to_unsigned(17130, LUT_AMPL_WIDTH - 1),
		27031 => to_unsigned(17128, LUT_AMPL_WIDTH - 1),
		27032 => to_unsigned(17125, LUT_AMPL_WIDTH - 1),
		27033 => to_unsigned(17122, LUT_AMPL_WIDTH - 1),
		27034 => to_unsigned(17120, LUT_AMPL_WIDTH - 1),
		27035 => to_unsigned(17117, LUT_AMPL_WIDTH - 1),
		27036 => to_unsigned(17114, LUT_AMPL_WIDTH - 1),
		27037 => to_unsigned(17112, LUT_AMPL_WIDTH - 1),
		27038 => to_unsigned(17109, LUT_AMPL_WIDTH - 1),
		27039 => to_unsigned(17106, LUT_AMPL_WIDTH - 1),
		27040 => to_unsigned(17104, LUT_AMPL_WIDTH - 1),
		27041 => to_unsigned(17101, LUT_AMPL_WIDTH - 1),
		27042 => to_unsigned(17098, LUT_AMPL_WIDTH - 1),
		27043 => to_unsigned(17096, LUT_AMPL_WIDTH - 1),
		27044 => to_unsigned(17093, LUT_AMPL_WIDTH - 1),
		27045 => to_unsigned(17090, LUT_AMPL_WIDTH - 1),
		27046 => to_unsigned(17087, LUT_AMPL_WIDTH - 1),
		27047 => to_unsigned(17085, LUT_AMPL_WIDTH - 1),
		27048 => to_unsigned(17082, LUT_AMPL_WIDTH - 1),
		27049 => to_unsigned(17079, LUT_AMPL_WIDTH - 1),
		27050 => to_unsigned(17077, LUT_AMPL_WIDTH - 1),
		27051 => to_unsigned(17074, LUT_AMPL_WIDTH - 1),
		27052 => to_unsigned(17071, LUT_AMPL_WIDTH - 1),
		27053 => to_unsigned(17069, LUT_AMPL_WIDTH - 1),
		27054 => to_unsigned(17066, LUT_AMPL_WIDTH - 1),
		27055 => to_unsigned(17063, LUT_AMPL_WIDTH - 1),
		27056 => to_unsigned(17061, LUT_AMPL_WIDTH - 1),
		27057 => to_unsigned(17058, LUT_AMPL_WIDTH - 1),
		27058 => to_unsigned(17055, LUT_AMPL_WIDTH - 1),
		27059 => to_unsigned(17053, LUT_AMPL_WIDTH - 1),
		27060 => to_unsigned(17050, LUT_AMPL_WIDTH - 1),
		27061 => to_unsigned(17047, LUT_AMPL_WIDTH - 1),
		27062 => to_unsigned(17045, LUT_AMPL_WIDTH - 1),
		27063 => to_unsigned(17042, LUT_AMPL_WIDTH - 1),
		27064 => to_unsigned(17039, LUT_AMPL_WIDTH - 1),
		27065 => to_unsigned(17037, LUT_AMPL_WIDTH - 1),
		27066 => to_unsigned(17034, LUT_AMPL_WIDTH - 1),
		27067 => to_unsigned(17031, LUT_AMPL_WIDTH - 1),
		27068 => to_unsigned(17028, LUT_AMPL_WIDTH - 1),
		27069 => to_unsigned(17026, LUT_AMPL_WIDTH - 1),
		27070 => to_unsigned(17023, LUT_AMPL_WIDTH - 1),
		27071 => to_unsigned(17020, LUT_AMPL_WIDTH - 1),
		27072 => to_unsigned(17018, LUT_AMPL_WIDTH - 1),
		27073 => to_unsigned(17015, LUT_AMPL_WIDTH - 1),
		27074 => to_unsigned(17012, LUT_AMPL_WIDTH - 1),
		27075 => to_unsigned(17010, LUT_AMPL_WIDTH - 1),
		27076 => to_unsigned(17007, LUT_AMPL_WIDTH - 1),
		27077 => to_unsigned(17004, LUT_AMPL_WIDTH - 1),
		27078 => to_unsigned(17002, LUT_AMPL_WIDTH - 1),
		27079 => to_unsigned(16999, LUT_AMPL_WIDTH - 1),
		27080 => to_unsigned(16996, LUT_AMPL_WIDTH - 1),
		27081 => to_unsigned(16994, LUT_AMPL_WIDTH - 1),
		27082 => to_unsigned(16991, LUT_AMPL_WIDTH - 1),
		27083 => to_unsigned(16988, LUT_AMPL_WIDTH - 1),
		27084 => to_unsigned(16986, LUT_AMPL_WIDTH - 1),
		27085 => to_unsigned(16983, LUT_AMPL_WIDTH - 1),
		27086 => to_unsigned(16980, LUT_AMPL_WIDTH - 1),
		27087 => to_unsigned(16977, LUT_AMPL_WIDTH - 1),
		27088 => to_unsigned(16975, LUT_AMPL_WIDTH - 1),
		27089 => to_unsigned(16972, LUT_AMPL_WIDTH - 1),
		27090 => to_unsigned(16969, LUT_AMPL_WIDTH - 1),
		27091 => to_unsigned(16967, LUT_AMPL_WIDTH - 1),
		27092 => to_unsigned(16964, LUT_AMPL_WIDTH - 1),
		27093 => to_unsigned(16961, LUT_AMPL_WIDTH - 1),
		27094 => to_unsigned(16959, LUT_AMPL_WIDTH - 1),
		27095 => to_unsigned(16956, LUT_AMPL_WIDTH - 1),
		27096 => to_unsigned(16953, LUT_AMPL_WIDTH - 1),
		27097 => to_unsigned(16951, LUT_AMPL_WIDTH - 1),
		27098 => to_unsigned(16948, LUT_AMPL_WIDTH - 1),
		27099 => to_unsigned(16945, LUT_AMPL_WIDTH - 1),
		27100 => to_unsigned(16943, LUT_AMPL_WIDTH - 1),
		27101 => to_unsigned(16940, LUT_AMPL_WIDTH - 1),
		27102 => to_unsigned(16937, LUT_AMPL_WIDTH - 1),
		27103 => to_unsigned(16934, LUT_AMPL_WIDTH - 1),
		27104 => to_unsigned(16932, LUT_AMPL_WIDTH - 1),
		27105 => to_unsigned(16929, LUT_AMPL_WIDTH - 1),
		27106 => to_unsigned(16926, LUT_AMPL_WIDTH - 1),
		27107 => to_unsigned(16924, LUT_AMPL_WIDTH - 1),
		27108 => to_unsigned(16921, LUT_AMPL_WIDTH - 1),
		27109 => to_unsigned(16918, LUT_AMPL_WIDTH - 1),
		27110 => to_unsigned(16916, LUT_AMPL_WIDTH - 1),
		27111 => to_unsigned(16913, LUT_AMPL_WIDTH - 1),
		27112 => to_unsigned(16910, LUT_AMPL_WIDTH - 1),
		27113 => to_unsigned(16908, LUT_AMPL_WIDTH - 1),
		27114 => to_unsigned(16905, LUT_AMPL_WIDTH - 1),
		27115 => to_unsigned(16902, LUT_AMPL_WIDTH - 1),
		27116 => to_unsigned(16899, LUT_AMPL_WIDTH - 1),
		27117 => to_unsigned(16897, LUT_AMPL_WIDTH - 1),
		27118 => to_unsigned(16894, LUT_AMPL_WIDTH - 1),
		27119 => to_unsigned(16891, LUT_AMPL_WIDTH - 1),
		27120 => to_unsigned(16889, LUT_AMPL_WIDTH - 1),
		27121 => to_unsigned(16886, LUT_AMPL_WIDTH - 1),
		27122 => to_unsigned(16883, LUT_AMPL_WIDTH - 1),
		27123 => to_unsigned(16881, LUT_AMPL_WIDTH - 1),
		27124 => to_unsigned(16878, LUT_AMPL_WIDTH - 1),
		27125 => to_unsigned(16875, LUT_AMPL_WIDTH - 1),
		27126 => to_unsigned(16873, LUT_AMPL_WIDTH - 1),
		27127 => to_unsigned(16870, LUT_AMPL_WIDTH - 1),
		27128 => to_unsigned(16867, LUT_AMPL_WIDTH - 1),
		27129 => to_unsigned(16864, LUT_AMPL_WIDTH - 1),
		27130 => to_unsigned(16862, LUT_AMPL_WIDTH - 1),
		27131 => to_unsigned(16859, LUT_AMPL_WIDTH - 1),
		27132 => to_unsigned(16856, LUT_AMPL_WIDTH - 1),
		27133 => to_unsigned(16854, LUT_AMPL_WIDTH - 1),
		27134 => to_unsigned(16851, LUT_AMPL_WIDTH - 1),
		27135 => to_unsigned(16848, LUT_AMPL_WIDTH - 1),
		27136 => to_unsigned(16846, LUT_AMPL_WIDTH - 1),
		27137 => to_unsigned(16843, LUT_AMPL_WIDTH - 1),
		27138 => to_unsigned(16840, LUT_AMPL_WIDTH - 1),
		27139 => to_unsigned(16838, LUT_AMPL_WIDTH - 1),
		27140 => to_unsigned(16835, LUT_AMPL_WIDTH - 1),
		27141 => to_unsigned(16832, LUT_AMPL_WIDTH - 1),
		27142 => to_unsigned(16829, LUT_AMPL_WIDTH - 1),
		27143 => to_unsigned(16827, LUT_AMPL_WIDTH - 1),
		27144 => to_unsigned(16824, LUT_AMPL_WIDTH - 1),
		27145 => to_unsigned(16821, LUT_AMPL_WIDTH - 1),
		27146 => to_unsigned(16819, LUT_AMPL_WIDTH - 1),
		27147 => to_unsigned(16816, LUT_AMPL_WIDTH - 1),
		27148 => to_unsigned(16813, LUT_AMPL_WIDTH - 1),
		27149 => to_unsigned(16811, LUT_AMPL_WIDTH - 1),
		27150 => to_unsigned(16808, LUT_AMPL_WIDTH - 1),
		27151 => to_unsigned(16805, LUT_AMPL_WIDTH - 1),
		27152 => to_unsigned(16802, LUT_AMPL_WIDTH - 1),
		27153 => to_unsigned(16800, LUT_AMPL_WIDTH - 1),
		27154 => to_unsigned(16797, LUT_AMPL_WIDTH - 1),
		27155 => to_unsigned(16794, LUT_AMPL_WIDTH - 1),
		27156 => to_unsigned(16792, LUT_AMPL_WIDTH - 1),
		27157 => to_unsigned(16789, LUT_AMPL_WIDTH - 1),
		27158 => to_unsigned(16786, LUT_AMPL_WIDTH - 1),
		27159 => to_unsigned(16784, LUT_AMPL_WIDTH - 1),
		27160 => to_unsigned(16781, LUT_AMPL_WIDTH - 1),
		27161 => to_unsigned(16778, LUT_AMPL_WIDTH - 1),
		27162 => to_unsigned(16775, LUT_AMPL_WIDTH - 1),
		27163 => to_unsigned(16773, LUT_AMPL_WIDTH - 1),
		27164 => to_unsigned(16770, LUT_AMPL_WIDTH - 1),
		27165 => to_unsigned(16767, LUT_AMPL_WIDTH - 1),
		27166 => to_unsigned(16765, LUT_AMPL_WIDTH - 1),
		27167 => to_unsigned(16762, LUT_AMPL_WIDTH - 1),
		27168 => to_unsigned(16759, LUT_AMPL_WIDTH - 1),
		27169 => to_unsigned(16757, LUT_AMPL_WIDTH - 1),
		27170 => to_unsigned(16754, LUT_AMPL_WIDTH - 1),
		27171 => to_unsigned(16751, LUT_AMPL_WIDTH - 1),
		27172 => to_unsigned(16749, LUT_AMPL_WIDTH - 1),
		27173 => to_unsigned(16746, LUT_AMPL_WIDTH - 1),
		27174 => to_unsigned(16743, LUT_AMPL_WIDTH - 1),
		27175 => to_unsigned(16740, LUT_AMPL_WIDTH - 1),
		27176 => to_unsigned(16738, LUT_AMPL_WIDTH - 1),
		27177 => to_unsigned(16735, LUT_AMPL_WIDTH - 1),
		27178 => to_unsigned(16732, LUT_AMPL_WIDTH - 1),
		27179 => to_unsigned(16730, LUT_AMPL_WIDTH - 1),
		27180 => to_unsigned(16727, LUT_AMPL_WIDTH - 1),
		27181 => to_unsigned(16724, LUT_AMPL_WIDTH - 1),
		27182 => to_unsigned(16721, LUT_AMPL_WIDTH - 1),
		27183 => to_unsigned(16719, LUT_AMPL_WIDTH - 1),
		27184 => to_unsigned(16716, LUT_AMPL_WIDTH - 1),
		27185 => to_unsigned(16713, LUT_AMPL_WIDTH - 1),
		27186 => to_unsigned(16711, LUT_AMPL_WIDTH - 1),
		27187 => to_unsigned(16708, LUT_AMPL_WIDTH - 1),
		27188 => to_unsigned(16705, LUT_AMPL_WIDTH - 1),
		27189 => to_unsigned(16703, LUT_AMPL_WIDTH - 1),
		27190 => to_unsigned(16700, LUT_AMPL_WIDTH - 1),
		27191 => to_unsigned(16697, LUT_AMPL_WIDTH - 1),
		27192 => to_unsigned(16694, LUT_AMPL_WIDTH - 1),
		27193 => to_unsigned(16692, LUT_AMPL_WIDTH - 1),
		27194 => to_unsigned(16689, LUT_AMPL_WIDTH - 1),
		27195 => to_unsigned(16686, LUT_AMPL_WIDTH - 1),
		27196 => to_unsigned(16684, LUT_AMPL_WIDTH - 1),
		27197 => to_unsigned(16681, LUT_AMPL_WIDTH - 1),
		27198 => to_unsigned(16678, LUT_AMPL_WIDTH - 1),
		27199 => to_unsigned(16676, LUT_AMPL_WIDTH - 1),
		27200 => to_unsigned(16673, LUT_AMPL_WIDTH - 1),
		27201 => to_unsigned(16670, LUT_AMPL_WIDTH - 1),
		27202 => to_unsigned(16667, LUT_AMPL_WIDTH - 1),
		27203 => to_unsigned(16665, LUT_AMPL_WIDTH - 1),
		27204 => to_unsigned(16662, LUT_AMPL_WIDTH - 1),
		27205 => to_unsigned(16659, LUT_AMPL_WIDTH - 1),
		27206 => to_unsigned(16657, LUT_AMPL_WIDTH - 1),
		27207 => to_unsigned(16654, LUT_AMPL_WIDTH - 1),
		27208 => to_unsigned(16651, LUT_AMPL_WIDTH - 1),
		27209 => to_unsigned(16648, LUT_AMPL_WIDTH - 1),
		27210 => to_unsigned(16646, LUT_AMPL_WIDTH - 1),
		27211 => to_unsigned(16643, LUT_AMPL_WIDTH - 1),
		27212 => to_unsigned(16640, LUT_AMPL_WIDTH - 1),
		27213 => to_unsigned(16638, LUT_AMPL_WIDTH - 1),
		27214 => to_unsigned(16635, LUT_AMPL_WIDTH - 1),
		27215 => to_unsigned(16632, LUT_AMPL_WIDTH - 1),
		27216 => to_unsigned(16630, LUT_AMPL_WIDTH - 1),
		27217 => to_unsigned(16627, LUT_AMPL_WIDTH - 1),
		27218 => to_unsigned(16624, LUT_AMPL_WIDTH - 1),
		27219 => to_unsigned(16621, LUT_AMPL_WIDTH - 1),
		27220 => to_unsigned(16619, LUT_AMPL_WIDTH - 1),
		27221 => to_unsigned(16616, LUT_AMPL_WIDTH - 1),
		27222 => to_unsigned(16613, LUT_AMPL_WIDTH - 1),
		27223 => to_unsigned(16611, LUT_AMPL_WIDTH - 1),
		27224 => to_unsigned(16608, LUT_AMPL_WIDTH - 1),
		27225 => to_unsigned(16605, LUT_AMPL_WIDTH - 1),
		27226 => to_unsigned(16602, LUT_AMPL_WIDTH - 1),
		27227 => to_unsigned(16600, LUT_AMPL_WIDTH - 1),
		27228 => to_unsigned(16597, LUT_AMPL_WIDTH - 1),
		27229 => to_unsigned(16594, LUT_AMPL_WIDTH - 1),
		27230 => to_unsigned(16592, LUT_AMPL_WIDTH - 1),
		27231 => to_unsigned(16589, LUT_AMPL_WIDTH - 1),
		27232 => to_unsigned(16586, LUT_AMPL_WIDTH - 1),
		27233 => to_unsigned(16584, LUT_AMPL_WIDTH - 1),
		27234 => to_unsigned(16581, LUT_AMPL_WIDTH - 1),
		27235 => to_unsigned(16578, LUT_AMPL_WIDTH - 1),
		27236 => to_unsigned(16575, LUT_AMPL_WIDTH - 1),
		27237 => to_unsigned(16573, LUT_AMPL_WIDTH - 1),
		27238 => to_unsigned(16570, LUT_AMPL_WIDTH - 1),
		27239 => to_unsigned(16567, LUT_AMPL_WIDTH - 1),
		27240 => to_unsigned(16565, LUT_AMPL_WIDTH - 1),
		27241 => to_unsigned(16562, LUT_AMPL_WIDTH - 1),
		27242 => to_unsigned(16559, LUT_AMPL_WIDTH - 1),
		27243 => to_unsigned(16556, LUT_AMPL_WIDTH - 1),
		27244 => to_unsigned(16554, LUT_AMPL_WIDTH - 1),
		27245 => to_unsigned(16551, LUT_AMPL_WIDTH - 1),
		27246 => to_unsigned(16548, LUT_AMPL_WIDTH - 1),
		27247 => to_unsigned(16546, LUT_AMPL_WIDTH - 1),
		27248 => to_unsigned(16543, LUT_AMPL_WIDTH - 1),
		27249 => to_unsigned(16540, LUT_AMPL_WIDTH - 1),
		27250 => to_unsigned(16537, LUT_AMPL_WIDTH - 1),
		27251 => to_unsigned(16535, LUT_AMPL_WIDTH - 1),
		27252 => to_unsigned(16532, LUT_AMPL_WIDTH - 1),
		27253 => to_unsigned(16529, LUT_AMPL_WIDTH - 1),
		27254 => to_unsigned(16527, LUT_AMPL_WIDTH - 1),
		27255 => to_unsigned(16524, LUT_AMPL_WIDTH - 1),
		27256 => to_unsigned(16521, LUT_AMPL_WIDTH - 1),
		27257 => to_unsigned(16518, LUT_AMPL_WIDTH - 1),
		27258 => to_unsigned(16516, LUT_AMPL_WIDTH - 1),
		27259 => to_unsigned(16513, LUT_AMPL_WIDTH - 1),
		27260 => to_unsigned(16510, LUT_AMPL_WIDTH - 1),
		27261 => to_unsigned(16508, LUT_AMPL_WIDTH - 1),
		27262 => to_unsigned(16505, LUT_AMPL_WIDTH - 1),
		27263 => to_unsigned(16502, LUT_AMPL_WIDTH - 1),
		27264 => to_unsigned(16499, LUT_AMPL_WIDTH - 1),
		27265 => to_unsigned(16497, LUT_AMPL_WIDTH - 1),
		27266 => to_unsigned(16494, LUT_AMPL_WIDTH - 1),
		27267 => to_unsigned(16491, LUT_AMPL_WIDTH - 1),
		27268 => to_unsigned(16489, LUT_AMPL_WIDTH - 1),
		27269 => to_unsigned(16486, LUT_AMPL_WIDTH - 1),
		27270 => to_unsigned(16483, LUT_AMPL_WIDTH - 1),
		27271 => to_unsigned(16480, LUT_AMPL_WIDTH - 1),
		27272 => to_unsigned(16478, LUT_AMPL_WIDTH - 1),
		27273 => to_unsigned(16475, LUT_AMPL_WIDTH - 1),
		27274 => to_unsigned(16472, LUT_AMPL_WIDTH - 1),
		27275 => to_unsigned(16470, LUT_AMPL_WIDTH - 1),
		27276 => to_unsigned(16467, LUT_AMPL_WIDTH - 1),
		27277 => to_unsigned(16464, LUT_AMPL_WIDTH - 1),
		27278 => to_unsigned(16461, LUT_AMPL_WIDTH - 1),
		27279 => to_unsigned(16459, LUT_AMPL_WIDTH - 1),
		27280 => to_unsigned(16456, LUT_AMPL_WIDTH - 1),
		27281 => to_unsigned(16453, LUT_AMPL_WIDTH - 1),
		27282 => to_unsigned(16451, LUT_AMPL_WIDTH - 1),
		27283 => to_unsigned(16448, LUT_AMPL_WIDTH - 1),
		27284 => to_unsigned(16445, LUT_AMPL_WIDTH - 1),
		27285 => to_unsigned(16442, LUT_AMPL_WIDTH - 1),
		27286 => to_unsigned(16440, LUT_AMPL_WIDTH - 1),
		27287 => to_unsigned(16437, LUT_AMPL_WIDTH - 1),
		27288 => to_unsigned(16434, LUT_AMPL_WIDTH - 1),
		27289 => to_unsigned(16432, LUT_AMPL_WIDTH - 1),
		27290 => to_unsigned(16429, LUT_AMPL_WIDTH - 1),
		27291 => to_unsigned(16426, LUT_AMPL_WIDTH - 1),
		27292 => to_unsigned(16423, LUT_AMPL_WIDTH - 1),
		27293 => to_unsigned(16421, LUT_AMPL_WIDTH - 1),
		27294 => to_unsigned(16418, LUT_AMPL_WIDTH - 1),
		27295 => to_unsigned(16415, LUT_AMPL_WIDTH - 1),
		27296 => to_unsigned(16413, LUT_AMPL_WIDTH - 1),
		27297 => to_unsigned(16410, LUT_AMPL_WIDTH - 1),
		27298 => to_unsigned(16407, LUT_AMPL_WIDTH - 1),
		27299 => to_unsigned(16404, LUT_AMPL_WIDTH - 1),
		27300 => to_unsigned(16402, LUT_AMPL_WIDTH - 1),
		27301 => to_unsigned(16399, LUT_AMPL_WIDTH - 1),
		27302 => to_unsigned(16396, LUT_AMPL_WIDTH - 1),
		27303 => to_unsigned(16393, LUT_AMPL_WIDTH - 1),
		27304 => to_unsigned(16391, LUT_AMPL_WIDTH - 1),
		27305 => to_unsigned(16388, LUT_AMPL_WIDTH - 1),
		27306 => to_unsigned(16385, LUT_AMPL_WIDTH - 1),
		27307 => to_unsigned(16383, LUT_AMPL_WIDTH - 1),
		27308 => to_unsigned(16380, LUT_AMPL_WIDTH - 1),
		27309 => to_unsigned(16377, LUT_AMPL_WIDTH - 1),
		27310 => to_unsigned(16374, LUT_AMPL_WIDTH - 1),
		27311 => to_unsigned(16372, LUT_AMPL_WIDTH - 1),
		27312 => to_unsigned(16369, LUT_AMPL_WIDTH - 1),
		27313 => to_unsigned(16366, LUT_AMPL_WIDTH - 1),
		27314 => to_unsigned(16364, LUT_AMPL_WIDTH - 1),
		27315 => to_unsigned(16361, LUT_AMPL_WIDTH - 1),
		27316 => to_unsigned(16358, LUT_AMPL_WIDTH - 1),
		27317 => to_unsigned(16355, LUT_AMPL_WIDTH - 1),
		27318 => to_unsigned(16353, LUT_AMPL_WIDTH - 1),
		27319 => to_unsigned(16350, LUT_AMPL_WIDTH - 1),
		27320 => to_unsigned(16347, LUT_AMPL_WIDTH - 1),
		27321 => to_unsigned(16344, LUT_AMPL_WIDTH - 1),
		27322 => to_unsigned(16342, LUT_AMPL_WIDTH - 1),
		27323 => to_unsigned(16339, LUT_AMPL_WIDTH - 1),
		27324 => to_unsigned(16336, LUT_AMPL_WIDTH - 1),
		27325 => to_unsigned(16334, LUT_AMPL_WIDTH - 1),
		27326 => to_unsigned(16331, LUT_AMPL_WIDTH - 1),
		27327 => to_unsigned(16328, LUT_AMPL_WIDTH - 1),
		27328 => to_unsigned(16325, LUT_AMPL_WIDTH - 1),
		27329 => to_unsigned(16323, LUT_AMPL_WIDTH - 1),
		27330 => to_unsigned(16320, LUT_AMPL_WIDTH - 1),
		27331 => to_unsigned(16317, LUT_AMPL_WIDTH - 1),
		27332 => to_unsigned(16315, LUT_AMPL_WIDTH - 1),
		27333 => to_unsigned(16312, LUT_AMPL_WIDTH - 1),
		27334 => to_unsigned(16309, LUT_AMPL_WIDTH - 1),
		27335 => to_unsigned(16306, LUT_AMPL_WIDTH - 1),
		27336 => to_unsigned(16304, LUT_AMPL_WIDTH - 1),
		27337 => to_unsigned(16301, LUT_AMPL_WIDTH - 1),
		27338 => to_unsigned(16298, LUT_AMPL_WIDTH - 1),
		27339 => to_unsigned(16295, LUT_AMPL_WIDTH - 1),
		27340 => to_unsigned(16293, LUT_AMPL_WIDTH - 1),
		27341 => to_unsigned(16290, LUT_AMPL_WIDTH - 1),
		27342 => to_unsigned(16287, LUT_AMPL_WIDTH - 1),
		27343 => to_unsigned(16285, LUT_AMPL_WIDTH - 1),
		27344 => to_unsigned(16282, LUT_AMPL_WIDTH - 1),
		27345 => to_unsigned(16279, LUT_AMPL_WIDTH - 1),
		27346 => to_unsigned(16276, LUT_AMPL_WIDTH - 1),
		27347 => to_unsigned(16274, LUT_AMPL_WIDTH - 1),
		27348 => to_unsigned(16271, LUT_AMPL_WIDTH - 1),
		27349 => to_unsigned(16268, LUT_AMPL_WIDTH - 1),
		27350 => to_unsigned(16265, LUT_AMPL_WIDTH - 1),
		27351 => to_unsigned(16263, LUT_AMPL_WIDTH - 1),
		27352 => to_unsigned(16260, LUT_AMPL_WIDTH - 1),
		27353 => to_unsigned(16257, LUT_AMPL_WIDTH - 1),
		27354 => to_unsigned(16255, LUT_AMPL_WIDTH - 1),
		27355 => to_unsigned(16252, LUT_AMPL_WIDTH - 1),
		27356 => to_unsigned(16249, LUT_AMPL_WIDTH - 1),
		27357 => to_unsigned(16246, LUT_AMPL_WIDTH - 1),
		27358 => to_unsigned(16244, LUT_AMPL_WIDTH - 1),
		27359 => to_unsigned(16241, LUT_AMPL_WIDTH - 1),
		27360 => to_unsigned(16238, LUT_AMPL_WIDTH - 1),
		27361 => to_unsigned(16235, LUT_AMPL_WIDTH - 1),
		27362 => to_unsigned(16233, LUT_AMPL_WIDTH - 1),
		27363 => to_unsigned(16230, LUT_AMPL_WIDTH - 1),
		27364 => to_unsigned(16227, LUT_AMPL_WIDTH - 1),
		27365 => to_unsigned(16225, LUT_AMPL_WIDTH - 1),
		27366 => to_unsigned(16222, LUT_AMPL_WIDTH - 1),
		27367 => to_unsigned(16219, LUT_AMPL_WIDTH - 1),
		27368 => to_unsigned(16216, LUT_AMPL_WIDTH - 1),
		27369 => to_unsigned(16214, LUT_AMPL_WIDTH - 1),
		27370 => to_unsigned(16211, LUT_AMPL_WIDTH - 1),
		27371 => to_unsigned(16208, LUT_AMPL_WIDTH - 1),
		27372 => to_unsigned(16205, LUT_AMPL_WIDTH - 1),
		27373 => to_unsigned(16203, LUT_AMPL_WIDTH - 1),
		27374 => to_unsigned(16200, LUT_AMPL_WIDTH - 1),
		27375 => to_unsigned(16197, LUT_AMPL_WIDTH - 1),
		27376 => to_unsigned(16195, LUT_AMPL_WIDTH - 1),
		27377 => to_unsigned(16192, LUT_AMPL_WIDTH - 1),
		27378 => to_unsigned(16189, LUT_AMPL_WIDTH - 1),
		27379 => to_unsigned(16186, LUT_AMPL_WIDTH - 1),
		27380 => to_unsigned(16184, LUT_AMPL_WIDTH - 1),
		27381 => to_unsigned(16181, LUT_AMPL_WIDTH - 1),
		27382 => to_unsigned(16178, LUT_AMPL_WIDTH - 1),
		27383 => to_unsigned(16175, LUT_AMPL_WIDTH - 1),
		27384 => to_unsigned(16173, LUT_AMPL_WIDTH - 1),
		27385 => to_unsigned(16170, LUT_AMPL_WIDTH - 1),
		27386 => to_unsigned(16167, LUT_AMPL_WIDTH - 1),
		27387 => to_unsigned(16164, LUT_AMPL_WIDTH - 1),
		27388 => to_unsigned(16162, LUT_AMPL_WIDTH - 1),
		27389 => to_unsigned(16159, LUT_AMPL_WIDTH - 1),
		27390 => to_unsigned(16156, LUT_AMPL_WIDTH - 1),
		27391 => to_unsigned(16154, LUT_AMPL_WIDTH - 1),
		27392 => to_unsigned(16151, LUT_AMPL_WIDTH - 1),
		27393 => to_unsigned(16148, LUT_AMPL_WIDTH - 1),
		27394 => to_unsigned(16145, LUT_AMPL_WIDTH - 1),
		27395 => to_unsigned(16143, LUT_AMPL_WIDTH - 1),
		27396 => to_unsigned(16140, LUT_AMPL_WIDTH - 1),
		27397 => to_unsigned(16137, LUT_AMPL_WIDTH - 1),
		27398 => to_unsigned(16134, LUT_AMPL_WIDTH - 1),
		27399 => to_unsigned(16132, LUT_AMPL_WIDTH - 1),
		27400 => to_unsigned(16129, LUT_AMPL_WIDTH - 1),
		27401 => to_unsigned(16126, LUT_AMPL_WIDTH - 1),
		27402 => to_unsigned(16123, LUT_AMPL_WIDTH - 1),
		27403 => to_unsigned(16121, LUT_AMPL_WIDTH - 1),
		27404 => to_unsigned(16118, LUT_AMPL_WIDTH - 1),
		27405 => to_unsigned(16115, LUT_AMPL_WIDTH - 1),
		27406 => to_unsigned(16113, LUT_AMPL_WIDTH - 1),
		27407 => to_unsigned(16110, LUT_AMPL_WIDTH - 1),
		27408 => to_unsigned(16107, LUT_AMPL_WIDTH - 1),
		27409 => to_unsigned(16104, LUT_AMPL_WIDTH - 1),
		27410 => to_unsigned(16102, LUT_AMPL_WIDTH - 1),
		27411 => to_unsigned(16099, LUT_AMPL_WIDTH - 1),
		27412 => to_unsigned(16096, LUT_AMPL_WIDTH - 1),
		27413 => to_unsigned(16093, LUT_AMPL_WIDTH - 1),
		27414 => to_unsigned(16091, LUT_AMPL_WIDTH - 1),
		27415 => to_unsigned(16088, LUT_AMPL_WIDTH - 1),
		27416 => to_unsigned(16085, LUT_AMPL_WIDTH - 1),
		27417 => to_unsigned(16082, LUT_AMPL_WIDTH - 1),
		27418 => to_unsigned(16080, LUT_AMPL_WIDTH - 1),
		27419 => to_unsigned(16077, LUT_AMPL_WIDTH - 1),
		27420 => to_unsigned(16074, LUT_AMPL_WIDTH - 1),
		27421 => to_unsigned(16071, LUT_AMPL_WIDTH - 1),
		27422 => to_unsigned(16069, LUT_AMPL_WIDTH - 1),
		27423 => to_unsigned(16066, LUT_AMPL_WIDTH - 1),
		27424 => to_unsigned(16063, LUT_AMPL_WIDTH - 1),
		27425 => to_unsigned(16061, LUT_AMPL_WIDTH - 1),
		27426 => to_unsigned(16058, LUT_AMPL_WIDTH - 1),
		27427 => to_unsigned(16055, LUT_AMPL_WIDTH - 1),
		27428 => to_unsigned(16052, LUT_AMPL_WIDTH - 1),
		27429 => to_unsigned(16050, LUT_AMPL_WIDTH - 1),
		27430 => to_unsigned(16047, LUT_AMPL_WIDTH - 1),
		27431 => to_unsigned(16044, LUT_AMPL_WIDTH - 1),
		27432 => to_unsigned(16041, LUT_AMPL_WIDTH - 1),
		27433 => to_unsigned(16039, LUT_AMPL_WIDTH - 1),
		27434 => to_unsigned(16036, LUT_AMPL_WIDTH - 1),
		27435 => to_unsigned(16033, LUT_AMPL_WIDTH - 1),
		27436 => to_unsigned(16030, LUT_AMPL_WIDTH - 1),
		27437 => to_unsigned(16028, LUT_AMPL_WIDTH - 1),
		27438 => to_unsigned(16025, LUT_AMPL_WIDTH - 1),
		27439 => to_unsigned(16022, LUT_AMPL_WIDTH - 1),
		27440 => to_unsigned(16019, LUT_AMPL_WIDTH - 1),
		27441 => to_unsigned(16017, LUT_AMPL_WIDTH - 1),
		27442 => to_unsigned(16014, LUT_AMPL_WIDTH - 1),
		27443 => to_unsigned(16011, LUT_AMPL_WIDTH - 1),
		27444 => to_unsigned(16008, LUT_AMPL_WIDTH - 1),
		27445 => to_unsigned(16006, LUT_AMPL_WIDTH - 1),
		27446 => to_unsigned(16003, LUT_AMPL_WIDTH - 1),
		27447 => to_unsigned(16000, LUT_AMPL_WIDTH - 1),
		27448 => to_unsigned(15997, LUT_AMPL_WIDTH - 1),
		27449 => to_unsigned(15995, LUT_AMPL_WIDTH - 1),
		27450 => to_unsigned(15992, LUT_AMPL_WIDTH - 1),
		27451 => to_unsigned(15989, LUT_AMPL_WIDTH - 1),
		27452 => to_unsigned(15987, LUT_AMPL_WIDTH - 1),
		27453 => to_unsigned(15984, LUT_AMPL_WIDTH - 1),
		27454 => to_unsigned(15981, LUT_AMPL_WIDTH - 1),
		27455 => to_unsigned(15978, LUT_AMPL_WIDTH - 1),
		27456 => to_unsigned(15976, LUT_AMPL_WIDTH - 1),
		27457 => to_unsigned(15973, LUT_AMPL_WIDTH - 1),
		27458 => to_unsigned(15970, LUT_AMPL_WIDTH - 1),
		27459 => to_unsigned(15967, LUT_AMPL_WIDTH - 1),
		27460 => to_unsigned(15965, LUT_AMPL_WIDTH - 1),
		27461 => to_unsigned(15962, LUT_AMPL_WIDTH - 1),
		27462 => to_unsigned(15959, LUT_AMPL_WIDTH - 1),
		27463 => to_unsigned(15956, LUT_AMPL_WIDTH - 1),
		27464 => to_unsigned(15954, LUT_AMPL_WIDTH - 1),
		27465 => to_unsigned(15951, LUT_AMPL_WIDTH - 1),
		27466 => to_unsigned(15948, LUT_AMPL_WIDTH - 1),
		27467 => to_unsigned(15945, LUT_AMPL_WIDTH - 1),
		27468 => to_unsigned(15943, LUT_AMPL_WIDTH - 1),
		27469 => to_unsigned(15940, LUT_AMPL_WIDTH - 1),
		27470 => to_unsigned(15937, LUT_AMPL_WIDTH - 1),
		27471 => to_unsigned(15934, LUT_AMPL_WIDTH - 1),
		27472 => to_unsigned(15932, LUT_AMPL_WIDTH - 1),
		27473 => to_unsigned(15929, LUT_AMPL_WIDTH - 1),
		27474 => to_unsigned(15926, LUT_AMPL_WIDTH - 1),
		27475 => to_unsigned(15923, LUT_AMPL_WIDTH - 1),
		27476 => to_unsigned(15921, LUT_AMPL_WIDTH - 1),
		27477 => to_unsigned(15918, LUT_AMPL_WIDTH - 1),
		27478 => to_unsigned(15915, LUT_AMPL_WIDTH - 1),
		27479 => to_unsigned(15912, LUT_AMPL_WIDTH - 1),
		27480 => to_unsigned(15910, LUT_AMPL_WIDTH - 1),
		27481 => to_unsigned(15907, LUT_AMPL_WIDTH - 1),
		27482 => to_unsigned(15904, LUT_AMPL_WIDTH - 1),
		27483 => to_unsigned(15901, LUT_AMPL_WIDTH - 1),
		27484 => to_unsigned(15899, LUT_AMPL_WIDTH - 1),
		27485 => to_unsigned(15896, LUT_AMPL_WIDTH - 1),
		27486 => to_unsigned(15893, LUT_AMPL_WIDTH - 1),
		27487 => to_unsigned(15890, LUT_AMPL_WIDTH - 1),
		27488 => to_unsigned(15888, LUT_AMPL_WIDTH - 1),
		27489 => to_unsigned(15885, LUT_AMPL_WIDTH - 1),
		27490 => to_unsigned(15882, LUT_AMPL_WIDTH - 1),
		27491 => to_unsigned(15879, LUT_AMPL_WIDTH - 1),
		27492 => to_unsigned(15877, LUT_AMPL_WIDTH - 1),
		27493 => to_unsigned(15874, LUT_AMPL_WIDTH - 1),
		27494 => to_unsigned(15871, LUT_AMPL_WIDTH - 1),
		27495 => to_unsigned(15868, LUT_AMPL_WIDTH - 1),
		27496 => to_unsigned(15866, LUT_AMPL_WIDTH - 1),
		27497 => to_unsigned(15863, LUT_AMPL_WIDTH - 1),
		27498 => to_unsigned(15860, LUT_AMPL_WIDTH - 1),
		27499 => to_unsigned(15857, LUT_AMPL_WIDTH - 1),
		27500 => to_unsigned(15855, LUT_AMPL_WIDTH - 1),
		27501 => to_unsigned(15852, LUT_AMPL_WIDTH - 1),
		27502 => to_unsigned(15849, LUT_AMPL_WIDTH - 1),
		27503 => to_unsigned(15846, LUT_AMPL_WIDTH - 1),
		27504 => to_unsigned(15844, LUT_AMPL_WIDTH - 1),
		27505 => to_unsigned(15841, LUT_AMPL_WIDTH - 1),
		27506 => to_unsigned(15838, LUT_AMPL_WIDTH - 1),
		27507 => to_unsigned(15835, LUT_AMPL_WIDTH - 1),
		27508 => to_unsigned(15833, LUT_AMPL_WIDTH - 1),
		27509 => to_unsigned(15830, LUT_AMPL_WIDTH - 1),
		27510 => to_unsigned(15827, LUT_AMPL_WIDTH - 1),
		27511 => to_unsigned(15824, LUT_AMPL_WIDTH - 1),
		27512 => to_unsigned(15822, LUT_AMPL_WIDTH - 1),
		27513 => to_unsigned(15819, LUT_AMPL_WIDTH - 1),
		27514 => to_unsigned(15816, LUT_AMPL_WIDTH - 1),
		27515 => to_unsigned(15813, LUT_AMPL_WIDTH - 1),
		27516 => to_unsigned(15811, LUT_AMPL_WIDTH - 1),
		27517 => to_unsigned(15808, LUT_AMPL_WIDTH - 1),
		27518 => to_unsigned(15805, LUT_AMPL_WIDTH - 1),
		27519 => to_unsigned(15802, LUT_AMPL_WIDTH - 1),
		27520 => to_unsigned(15800, LUT_AMPL_WIDTH - 1),
		27521 => to_unsigned(15797, LUT_AMPL_WIDTH - 1),
		27522 => to_unsigned(15794, LUT_AMPL_WIDTH - 1),
		27523 => to_unsigned(15791, LUT_AMPL_WIDTH - 1),
		27524 => to_unsigned(15789, LUT_AMPL_WIDTH - 1),
		27525 => to_unsigned(15786, LUT_AMPL_WIDTH - 1),
		27526 => to_unsigned(15783, LUT_AMPL_WIDTH - 1),
		27527 => to_unsigned(15780, LUT_AMPL_WIDTH - 1),
		27528 => to_unsigned(15778, LUT_AMPL_WIDTH - 1),
		27529 => to_unsigned(15775, LUT_AMPL_WIDTH - 1),
		27530 => to_unsigned(15772, LUT_AMPL_WIDTH - 1),
		27531 => to_unsigned(15769, LUT_AMPL_WIDTH - 1),
		27532 => to_unsigned(15767, LUT_AMPL_WIDTH - 1),
		27533 => to_unsigned(15764, LUT_AMPL_WIDTH - 1),
		27534 => to_unsigned(15761, LUT_AMPL_WIDTH - 1),
		27535 => to_unsigned(15758, LUT_AMPL_WIDTH - 1),
		27536 => to_unsigned(15756, LUT_AMPL_WIDTH - 1),
		27537 => to_unsigned(15753, LUT_AMPL_WIDTH - 1),
		27538 => to_unsigned(15750, LUT_AMPL_WIDTH - 1),
		27539 => to_unsigned(15747, LUT_AMPL_WIDTH - 1),
		27540 => to_unsigned(15745, LUT_AMPL_WIDTH - 1),
		27541 => to_unsigned(15742, LUT_AMPL_WIDTH - 1),
		27542 => to_unsigned(15739, LUT_AMPL_WIDTH - 1),
		27543 => to_unsigned(15736, LUT_AMPL_WIDTH - 1),
		27544 => to_unsigned(15734, LUT_AMPL_WIDTH - 1),
		27545 => to_unsigned(15731, LUT_AMPL_WIDTH - 1),
		27546 => to_unsigned(15728, LUT_AMPL_WIDTH - 1),
		27547 => to_unsigned(15725, LUT_AMPL_WIDTH - 1),
		27548 => to_unsigned(15723, LUT_AMPL_WIDTH - 1),
		27549 => to_unsigned(15720, LUT_AMPL_WIDTH - 1),
		27550 => to_unsigned(15717, LUT_AMPL_WIDTH - 1),
		27551 => to_unsigned(15714, LUT_AMPL_WIDTH - 1),
		27552 => to_unsigned(15712, LUT_AMPL_WIDTH - 1),
		27553 => to_unsigned(15709, LUT_AMPL_WIDTH - 1),
		27554 => to_unsigned(15706, LUT_AMPL_WIDTH - 1),
		27555 => to_unsigned(15703, LUT_AMPL_WIDTH - 1),
		27556 => to_unsigned(15701, LUT_AMPL_WIDTH - 1),
		27557 => to_unsigned(15698, LUT_AMPL_WIDTH - 1),
		27558 => to_unsigned(15695, LUT_AMPL_WIDTH - 1),
		27559 => to_unsigned(15692, LUT_AMPL_WIDTH - 1),
		27560 => to_unsigned(15690, LUT_AMPL_WIDTH - 1),
		27561 => to_unsigned(15687, LUT_AMPL_WIDTH - 1),
		27562 => to_unsigned(15684, LUT_AMPL_WIDTH - 1),
		27563 => to_unsigned(15681, LUT_AMPL_WIDTH - 1),
		27564 => to_unsigned(15678, LUT_AMPL_WIDTH - 1),
		27565 => to_unsigned(15676, LUT_AMPL_WIDTH - 1),
		27566 => to_unsigned(15673, LUT_AMPL_WIDTH - 1),
		27567 => to_unsigned(15670, LUT_AMPL_WIDTH - 1),
		27568 => to_unsigned(15667, LUT_AMPL_WIDTH - 1),
		27569 => to_unsigned(15665, LUT_AMPL_WIDTH - 1),
		27570 => to_unsigned(15662, LUT_AMPL_WIDTH - 1),
		27571 => to_unsigned(15659, LUT_AMPL_WIDTH - 1),
		27572 => to_unsigned(15656, LUT_AMPL_WIDTH - 1),
		27573 => to_unsigned(15654, LUT_AMPL_WIDTH - 1),
		27574 => to_unsigned(15651, LUT_AMPL_WIDTH - 1),
		27575 => to_unsigned(15648, LUT_AMPL_WIDTH - 1),
		27576 => to_unsigned(15645, LUT_AMPL_WIDTH - 1),
		27577 => to_unsigned(15643, LUT_AMPL_WIDTH - 1),
		27578 => to_unsigned(15640, LUT_AMPL_WIDTH - 1),
		27579 => to_unsigned(15637, LUT_AMPL_WIDTH - 1),
		27580 => to_unsigned(15634, LUT_AMPL_WIDTH - 1),
		27581 => to_unsigned(15632, LUT_AMPL_WIDTH - 1),
		27582 => to_unsigned(15629, LUT_AMPL_WIDTH - 1),
		27583 => to_unsigned(15626, LUT_AMPL_WIDTH - 1),
		27584 => to_unsigned(15623, LUT_AMPL_WIDTH - 1),
		27585 => to_unsigned(15621, LUT_AMPL_WIDTH - 1),
		27586 => to_unsigned(15618, LUT_AMPL_WIDTH - 1),
		27587 => to_unsigned(15615, LUT_AMPL_WIDTH - 1),
		27588 => to_unsigned(15612, LUT_AMPL_WIDTH - 1),
		27589 => to_unsigned(15609, LUT_AMPL_WIDTH - 1),
		27590 => to_unsigned(15607, LUT_AMPL_WIDTH - 1),
		27591 => to_unsigned(15604, LUT_AMPL_WIDTH - 1),
		27592 => to_unsigned(15601, LUT_AMPL_WIDTH - 1),
		27593 => to_unsigned(15598, LUT_AMPL_WIDTH - 1),
		27594 => to_unsigned(15596, LUT_AMPL_WIDTH - 1),
		27595 => to_unsigned(15593, LUT_AMPL_WIDTH - 1),
		27596 => to_unsigned(15590, LUT_AMPL_WIDTH - 1),
		27597 => to_unsigned(15587, LUT_AMPL_WIDTH - 1),
		27598 => to_unsigned(15585, LUT_AMPL_WIDTH - 1),
		27599 => to_unsigned(15582, LUT_AMPL_WIDTH - 1),
		27600 => to_unsigned(15579, LUT_AMPL_WIDTH - 1),
		27601 => to_unsigned(15576, LUT_AMPL_WIDTH - 1),
		27602 => to_unsigned(15574, LUT_AMPL_WIDTH - 1),
		27603 => to_unsigned(15571, LUT_AMPL_WIDTH - 1),
		27604 => to_unsigned(15568, LUT_AMPL_WIDTH - 1),
		27605 => to_unsigned(15565, LUT_AMPL_WIDTH - 1),
		27606 => to_unsigned(15562, LUT_AMPL_WIDTH - 1),
		27607 => to_unsigned(15560, LUT_AMPL_WIDTH - 1),
		27608 => to_unsigned(15557, LUT_AMPL_WIDTH - 1),
		27609 => to_unsigned(15554, LUT_AMPL_WIDTH - 1),
		27610 => to_unsigned(15551, LUT_AMPL_WIDTH - 1),
		27611 => to_unsigned(15549, LUT_AMPL_WIDTH - 1),
		27612 => to_unsigned(15546, LUT_AMPL_WIDTH - 1),
		27613 => to_unsigned(15543, LUT_AMPL_WIDTH - 1),
		27614 => to_unsigned(15540, LUT_AMPL_WIDTH - 1),
		27615 => to_unsigned(15538, LUT_AMPL_WIDTH - 1),
		27616 => to_unsigned(15535, LUT_AMPL_WIDTH - 1),
		27617 => to_unsigned(15532, LUT_AMPL_WIDTH - 1),
		27618 => to_unsigned(15529, LUT_AMPL_WIDTH - 1),
		27619 => to_unsigned(15527, LUT_AMPL_WIDTH - 1),
		27620 => to_unsigned(15524, LUT_AMPL_WIDTH - 1),
		27621 => to_unsigned(15521, LUT_AMPL_WIDTH - 1),
		27622 => to_unsigned(15518, LUT_AMPL_WIDTH - 1),
		27623 => to_unsigned(15515, LUT_AMPL_WIDTH - 1),
		27624 => to_unsigned(15513, LUT_AMPL_WIDTH - 1),
		27625 => to_unsigned(15510, LUT_AMPL_WIDTH - 1),
		27626 => to_unsigned(15507, LUT_AMPL_WIDTH - 1),
		27627 => to_unsigned(15504, LUT_AMPL_WIDTH - 1),
		27628 => to_unsigned(15502, LUT_AMPL_WIDTH - 1),
		27629 => to_unsigned(15499, LUT_AMPL_WIDTH - 1),
		27630 => to_unsigned(15496, LUT_AMPL_WIDTH - 1),
		27631 => to_unsigned(15493, LUT_AMPL_WIDTH - 1),
		27632 => to_unsigned(15491, LUT_AMPL_WIDTH - 1),
		27633 => to_unsigned(15488, LUT_AMPL_WIDTH - 1),
		27634 => to_unsigned(15485, LUT_AMPL_WIDTH - 1),
		27635 => to_unsigned(15482, LUT_AMPL_WIDTH - 1),
		27636 => to_unsigned(15479, LUT_AMPL_WIDTH - 1),
		27637 => to_unsigned(15477, LUT_AMPL_WIDTH - 1),
		27638 => to_unsigned(15474, LUT_AMPL_WIDTH - 1),
		27639 => to_unsigned(15471, LUT_AMPL_WIDTH - 1),
		27640 => to_unsigned(15468, LUT_AMPL_WIDTH - 1),
		27641 => to_unsigned(15466, LUT_AMPL_WIDTH - 1),
		27642 => to_unsigned(15463, LUT_AMPL_WIDTH - 1),
		27643 => to_unsigned(15460, LUT_AMPL_WIDTH - 1),
		27644 => to_unsigned(15457, LUT_AMPL_WIDTH - 1),
		27645 => to_unsigned(15455, LUT_AMPL_WIDTH - 1),
		27646 => to_unsigned(15452, LUT_AMPL_WIDTH - 1),
		27647 => to_unsigned(15449, LUT_AMPL_WIDTH - 1),
		27648 => to_unsigned(15446, LUT_AMPL_WIDTH - 1),
		27649 => to_unsigned(15443, LUT_AMPL_WIDTH - 1),
		27650 => to_unsigned(15441, LUT_AMPL_WIDTH - 1),
		27651 => to_unsigned(15438, LUT_AMPL_WIDTH - 1),
		27652 => to_unsigned(15435, LUT_AMPL_WIDTH - 1),
		27653 => to_unsigned(15432, LUT_AMPL_WIDTH - 1),
		27654 => to_unsigned(15430, LUT_AMPL_WIDTH - 1),
		27655 => to_unsigned(15427, LUT_AMPL_WIDTH - 1),
		27656 => to_unsigned(15424, LUT_AMPL_WIDTH - 1),
		27657 => to_unsigned(15421, LUT_AMPL_WIDTH - 1),
		27658 => to_unsigned(15419, LUT_AMPL_WIDTH - 1),
		27659 => to_unsigned(15416, LUT_AMPL_WIDTH - 1),
		27660 => to_unsigned(15413, LUT_AMPL_WIDTH - 1),
		27661 => to_unsigned(15410, LUT_AMPL_WIDTH - 1),
		27662 => to_unsigned(15407, LUT_AMPL_WIDTH - 1),
		27663 => to_unsigned(15405, LUT_AMPL_WIDTH - 1),
		27664 => to_unsigned(15402, LUT_AMPL_WIDTH - 1),
		27665 => to_unsigned(15399, LUT_AMPL_WIDTH - 1),
		27666 => to_unsigned(15396, LUT_AMPL_WIDTH - 1),
		27667 => to_unsigned(15394, LUT_AMPL_WIDTH - 1),
		27668 => to_unsigned(15391, LUT_AMPL_WIDTH - 1),
		27669 => to_unsigned(15388, LUT_AMPL_WIDTH - 1),
		27670 => to_unsigned(15385, LUT_AMPL_WIDTH - 1),
		27671 => to_unsigned(15382, LUT_AMPL_WIDTH - 1),
		27672 => to_unsigned(15380, LUT_AMPL_WIDTH - 1),
		27673 => to_unsigned(15377, LUT_AMPL_WIDTH - 1),
		27674 => to_unsigned(15374, LUT_AMPL_WIDTH - 1),
		27675 => to_unsigned(15371, LUT_AMPL_WIDTH - 1),
		27676 => to_unsigned(15369, LUT_AMPL_WIDTH - 1),
		27677 => to_unsigned(15366, LUT_AMPL_WIDTH - 1),
		27678 => to_unsigned(15363, LUT_AMPL_WIDTH - 1),
		27679 => to_unsigned(15360, LUT_AMPL_WIDTH - 1),
		27680 => to_unsigned(15358, LUT_AMPL_WIDTH - 1),
		27681 => to_unsigned(15355, LUT_AMPL_WIDTH - 1),
		27682 => to_unsigned(15352, LUT_AMPL_WIDTH - 1),
		27683 => to_unsigned(15349, LUT_AMPL_WIDTH - 1),
		27684 => to_unsigned(15346, LUT_AMPL_WIDTH - 1),
		27685 => to_unsigned(15344, LUT_AMPL_WIDTH - 1),
		27686 => to_unsigned(15341, LUT_AMPL_WIDTH - 1),
		27687 => to_unsigned(15338, LUT_AMPL_WIDTH - 1),
		27688 => to_unsigned(15335, LUT_AMPL_WIDTH - 1),
		27689 => to_unsigned(15333, LUT_AMPL_WIDTH - 1),
		27690 => to_unsigned(15330, LUT_AMPL_WIDTH - 1),
		27691 => to_unsigned(15327, LUT_AMPL_WIDTH - 1),
		27692 => to_unsigned(15324, LUT_AMPL_WIDTH - 1),
		27693 => to_unsigned(15321, LUT_AMPL_WIDTH - 1),
		27694 => to_unsigned(15319, LUT_AMPL_WIDTH - 1),
		27695 => to_unsigned(15316, LUT_AMPL_WIDTH - 1),
		27696 => to_unsigned(15313, LUT_AMPL_WIDTH - 1),
		27697 => to_unsigned(15310, LUT_AMPL_WIDTH - 1),
		27698 => to_unsigned(15308, LUT_AMPL_WIDTH - 1),
		27699 => to_unsigned(15305, LUT_AMPL_WIDTH - 1),
		27700 => to_unsigned(15302, LUT_AMPL_WIDTH - 1),
		27701 => to_unsigned(15299, LUT_AMPL_WIDTH - 1),
		27702 => to_unsigned(15296, LUT_AMPL_WIDTH - 1),
		27703 => to_unsigned(15294, LUT_AMPL_WIDTH - 1),
		27704 => to_unsigned(15291, LUT_AMPL_WIDTH - 1),
		27705 => to_unsigned(15288, LUT_AMPL_WIDTH - 1),
		27706 => to_unsigned(15285, LUT_AMPL_WIDTH - 1),
		27707 => to_unsigned(15283, LUT_AMPL_WIDTH - 1),
		27708 => to_unsigned(15280, LUT_AMPL_WIDTH - 1),
		27709 => to_unsigned(15277, LUT_AMPL_WIDTH - 1),
		27710 => to_unsigned(15274, LUT_AMPL_WIDTH - 1),
		27711 => to_unsigned(15271, LUT_AMPL_WIDTH - 1),
		27712 => to_unsigned(15269, LUT_AMPL_WIDTH - 1),
		27713 => to_unsigned(15266, LUT_AMPL_WIDTH - 1),
		27714 => to_unsigned(15263, LUT_AMPL_WIDTH - 1),
		27715 => to_unsigned(15260, LUT_AMPL_WIDTH - 1),
		27716 => to_unsigned(15258, LUT_AMPL_WIDTH - 1),
		27717 => to_unsigned(15255, LUT_AMPL_WIDTH - 1),
		27718 => to_unsigned(15252, LUT_AMPL_WIDTH - 1),
		27719 => to_unsigned(15249, LUT_AMPL_WIDTH - 1),
		27720 => to_unsigned(15246, LUT_AMPL_WIDTH - 1),
		27721 => to_unsigned(15244, LUT_AMPL_WIDTH - 1),
		27722 => to_unsigned(15241, LUT_AMPL_WIDTH - 1),
		27723 => to_unsigned(15238, LUT_AMPL_WIDTH - 1),
		27724 => to_unsigned(15235, LUT_AMPL_WIDTH - 1),
		27725 => to_unsigned(15233, LUT_AMPL_WIDTH - 1),
		27726 => to_unsigned(15230, LUT_AMPL_WIDTH - 1),
		27727 => to_unsigned(15227, LUT_AMPL_WIDTH - 1),
		27728 => to_unsigned(15224, LUT_AMPL_WIDTH - 1),
		27729 => to_unsigned(15221, LUT_AMPL_WIDTH - 1),
		27730 => to_unsigned(15219, LUT_AMPL_WIDTH - 1),
		27731 => to_unsigned(15216, LUT_AMPL_WIDTH - 1),
		27732 => to_unsigned(15213, LUT_AMPL_WIDTH - 1),
		27733 => to_unsigned(15210, LUT_AMPL_WIDTH - 1),
		27734 => to_unsigned(15207, LUT_AMPL_WIDTH - 1),
		27735 => to_unsigned(15205, LUT_AMPL_WIDTH - 1),
		27736 => to_unsigned(15202, LUT_AMPL_WIDTH - 1),
		27737 => to_unsigned(15199, LUT_AMPL_WIDTH - 1),
		27738 => to_unsigned(15196, LUT_AMPL_WIDTH - 1),
		27739 => to_unsigned(15194, LUT_AMPL_WIDTH - 1),
		27740 => to_unsigned(15191, LUT_AMPL_WIDTH - 1),
		27741 => to_unsigned(15188, LUT_AMPL_WIDTH - 1),
		27742 => to_unsigned(15185, LUT_AMPL_WIDTH - 1),
		27743 => to_unsigned(15182, LUT_AMPL_WIDTH - 1),
		27744 => to_unsigned(15180, LUT_AMPL_WIDTH - 1),
		27745 => to_unsigned(15177, LUT_AMPL_WIDTH - 1),
		27746 => to_unsigned(15174, LUT_AMPL_WIDTH - 1),
		27747 => to_unsigned(15171, LUT_AMPL_WIDTH - 1),
		27748 => to_unsigned(15168, LUT_AMPL_WIDTH - 1),
		27749 => to_unsigned(15166, LUT_AMPL_WIDTH - 1),
		27750 => to_unsigned(15163, LUT_AMPL_WIDTH - 1),
		27751 => to_unsigned(15160, LUT_AMPL_WIDTH - 1),
		27752 => to_unsigned(15157, LUT_AMPL_WIDTH - 1),
		27753 => to_unsigned(15155, LUT_AMPL_WIDTH - 1),
		27754 => to_unsigned(15152, LUT_AMPL_WIDTH - 1),
		27755 => to_unsigned(15149, LUT_AMPL_WIDTH - 1),
		27756 => to_unsigned(15146, LUT_AMPL_WIDTH - 1),
		27757 => to_unsigned(15143, LUT_AMPL_WIDTH - 1),
		27758 => to_unsigned(15141, LUT_AMPL_WIDTH - 1),
		27759 => to_unsigned(15138, LUT_AMPL_WIDTH - 1),
		27760 => to_unsigned(15135, LUT_AMPL_WIDTH - 1),
		27761 => to_unsigned(15132, LUT_AMPL_WIDTH - 1),
		27762 => to_unsigned(15129, LUT_AMPL_WIDTH - 1),
		27763 => to_unsigned(15127, LUT_AMPL_WIDTH - 1),
		27764 => to_unsigned(15124, LUT_AMPL_WIDTH - 1),
		27765 => to_unsigned(15121, LUT_AMPL_WIDTH - 1),
		27766 => to_unsigned(15118, LUT_AMPL_WIDTH - 1),
		27767 => to_unsigned(15116, LUT_AMPL_WIDTH - 1),
		27768 => to_unsigned(15113, LUT_AMPL_WIDTH - 1),
		27769 => to_unsigned(15110, LUT_AMPL_WIDTH - 1),
		27770 => to_unsigned(15107, LUT_AMPL_WIDTH - 1),
		27771 => to_unsigned(15104, LUT_AMPL_WIDTH - 1),
		27772 => to_unsigned(15102, LUT_AMPL_WIDTH - 1),
		27773 => to_unsigned(15099, LUT_AMPL_WIDTH - 1),
		27774 => to_unsigned(15096, LUT_AMPL_WIDTH - 1),
		27775 => to_unsigned(15093, LUT_AMPL_WIDTH - 1),
		27776 => to_unsigned(15090, LUT_AMPL_WIDTH - 1),
		27777 => to_unsigned(15088, LUT_AMPL_WIDTH - 1),
		27778 => to_unsigned(15085, LUT_AMPL_WIDTH - 1),
		27779 => to_unsigned(15082, LUT_AMPL_WIDTH - 1),
		27780 => to_unsigned(15079, LUT_AMPL_WIDTH - 1),
		27781 => to_unsigned(15077, LUT_AMPL_WIDTH - 1),
		27782 => to_unsigned(15074, LUT_AMPL_WIDTH - 1),
		27783 => to_unsigned(15071, LUT_AMPL_WIDTH - 1),
		27784 => to_unsigned(15068, LUT_AMPL_WIDTH - 1),
		27785 => to_unsigned(15065, LUT_AMPL_WIDTH - 1),
		27786 => to_unsigned(15063, LUT_AMPL_WIDTH - 1),
		27787 => to_unsigned(15060, LUT_AMPL_WIDTH - 1),
		27788 => to_unsigned(15057, LUT_AMPL_WIDTH - 1),
		27789 => to_unsigned(15054, LUT_AMPL_WIDTH - 1),
		27790 => to_unsigned(15051, LUT_AMPL_WIDTH - 1),
		27791 => to_unsigned(15049, LUT_AMPL_WIDTH - 1),
		27792 => to_unsigned(15046, LUT_AMPL_WIDTH - 1),
		27793 => to_unsigned(15043, LUT_AMPL_WIDTH - 1),
		27794 => to_unsigned(15040, LUT_AMPL_WIDTH - 1),
		27795 => to_unsigned(15037, LUT_AMPL_WIDTH - 1),
		27796 => to_unsigned(15035, LUT_AMPL_WIDTH - 1),
		27797 => to_unsigned(15032, LUT_AMPL_WIDTH - 1),
		27798 => to_unsigned(15029, LUT_AMPL_WIDTH - 1),
		27799 => to_unsigned(15026, LUT_AMPL_WIDTH - 1),
		27800 => to_unsigned(15024, LUT_AMPL_WIDTH - 1),
		27801 => to_unsigned(15021, LUT_AMPL_WIDTH - 1),
		27802 => to_unsigned(15018, LUT_AMPL_WIDTH - 1),
		27803 => to_unsigned(15015, LUT_AMPL_WIDTH - 1),
		27804 => to_unsigned(15012, LUT_AMPL_WIDTH - 1),
		27805 => to_unsigned(15010, LUT_AMPL_WIDTH - 1),
		27806 => to_unsigned(15007, LUT_AMPL_WIDTH - 1),
		27807 => to_unsigned(15004, LUT_AMPL_WIDTH - 1),
		27808 => to_unsigned(15001, LUT_AMPL_WIDTH - 1),
		27809 => to_unsigned(14998, LUT_AMPL_WIDTH - 1),
		27810 => to_unsigned(14996, LUT_AMPL_WIDTH - 1),
		27811 => to_unsigned(14993, LUT_AMPL_WIDTH - 1),
		27812 => to_unsigned(14990, LUT_AMPL_WIDTH - 1),
		27813 => to_unsigned(14987, LUT_AMPL_WIDTH - 1),
		27814 => to_unsigned(14984, LUT_AMPL_WIDTH - 1),
		27815 => to_unsigned(14982, LUT_AMPL_WIDTH - 1),
		27816 => to_unsigned(14979, LUT_AMPL_WIDTH - 1),
		27817 => to_unsigned(14976, LUT_AMPL_WIDTH - 1),
		27818 => to_unsigned(14973, LUT_AMPL_WIDTH - 1),
		27819 => to_unsigned(14970, LUT_AMPL_WIDTH - 1),
		27820 => to_unsigned(14968, LUT_AMPL_WIDTH - 1),
		27821 => to_unsigned(14965, LUT_AMPL_WIDTH - 1),
		27822 => to_unsigned(14962, LUT_AMPL_WIDTH - 1),
		27823 => to_unsigned(14959, LUT_AMPL_WIDTH - 1),
		27824 => to_unsigned(14956, LUT_AMPL_WIDTH - 1),
		27825 => to_unsigned(14954, LUT_AMPL_WIDTH - 1),
		27826 => to_unsigned(14951, LUT_AMPL_WIDTH - 1),
		27827 => to_unsigned(14948, LUT_AMPL_WIDTH - 1),
		27828 => to_unsigned(14945, LUT_AMPL_WIDTH - 1),
		27829 => to_unsigned(14942, LUT_AMPL_WIDTH - 1),
		27830 => to_unsigned(14940, LUT_AMPL_WIDTH - 1),
		27831 => to_unsigned(14937, LUT_AMPL_WIDTH - 1),
		27832 => to_unsigned(14934, LUT_AMPL_WIDTH - 1),
		27833 => to_unsigned(14931, LUT_AMPL_WIDTH - 1),
		27834 => to_unsigned(14929, LUT_AMPL_WIDTH - 1),
		27835 => to_unsigned(14926, LUT_AMPL_WIDTH - 1),
		27836 => to_unsigned(14923, LUT_AMPL_WIDTH - 1),
		27837 => to_unsigned(14920, LUT_AMPL_WIDTH - 1),
		27838 => to_unsigned(14917, LUT_AMPL_WIDTH - 1),
		27839 => to_unsigned(14915, LUT_AMPL_WIDTH - 1),
		27840 => to_unsigned(14912, LUT_AMPL_WIDTH - 1),
		27841 => to_unsigned(14909, LUT_AMPL_WIDTH - 1),
		27842 => to_unsigned(14906, LUT_AMPL_WIDTH - 1),
		27843 => to_unsigned(14903, LUT_AMPL_WIDTH - 1),
		27844 => to_unsigned(14901, LUT_AMPL_WIDTH - 1),
		27845 => to_unsigned(14898, LUT_AMPL_WIDTH - 1),
		27846 => to_unsigned(14895, LUT_AMPL_WIDTH - 1),
		27847 => to_unsigned(14892, LUT_AMPL_WIDTH - 1),
		27848 => to_unsigned(14889, LUT_AMPL_WIDTH - 1),
		27849 => to_unsigned(14887, LUT_AMPL_WIDTH - 1),
		27850 => to_unsigned(14884, LUT_AMPL_WIDTH - 1),
		27851 => to_unsigned(14881, LUT_AMPL_WIDTH - 1),
		27852 => to_unsigned(14878, LUT_AMPL_WIDTH - 1),
		27853 => to_unsigned(14875, LUT_AMPL_WIDTH - 1),
		27854 => to_unsigned(14873, LUT_AMPL_WIDTH - 1),
		27855 => to_unsigned(14870, LUT_AMPL_WIDTH - 1),
		27856 => to_unsigned(14867, LUT_AMPL_WIDTH - 1),
		27857 => to_unsigned(14864, LUT_AMPL_WIDTH - 1),
		27858 => to_unsigned(14861, LUT_AMPL_WIDTH - 1),
		27859 => to_unsigned(14859, LUT_AMPL_WIDTH - 1),
		27860 => to_unsigned(14856, LUT_AMPL_WIDTH - 1),
		27861 => to_unsigned(14853, LUT_AMPL_WIDTH - 1),
		27862 => to_unsigned(14850, LUT_AMPL_WIDTH - 1),
		27863 => to_unsigned(14847, LUT_AMPL_WIDTH - 1),
		27864 => to_unsigned(14845, LUT_AMPL_WIDTH - 1),
		27865 => to_unsigned(14842, LUT_AMPL_WIDTH - 1),
		27866 => to_unsigned(14839, LUT_AMPL_WIDTH - 1),
		27867 => to_unsigned(14836, LUT_AMPL_WIDTH - 1),
		27868 => to_unsigned(14833, LUT_AMPL_WIDTH - 1),
		27869 => to_unsigned(14831, LUT_AMPL_WIDTH - 1),
		27870 => to_unsigned(14828, LUT_AMPL_WIDTH - 1),
		27871 => to_unsigned(14825, LUT_AMPL_WIDTH - 1),
		27872 => to_unsigned(14822, LUT_AMPL_WIDTH - 1),
		27873 => to_unsigned(14819, LUT_AMPL_WIDTH - 1),
		27874 => to_unsigned(14817, LUT_AMPL_WIDTH - 1),
		27875 => to_unsigned(14814, LUT_AMPL_WIDTH - 1),
		27876 => to_unsigned(14811, LUT_AMPL_WIDTH - 1),
		27877 => to_unsigned(14808, LUT_AMPL_WIDTH - 1),
		27878 => to_unsigned(14805, LUT_AMPL_WIDTH - 1),
		27879 => to_unsigned(14803, LUT_AMPL_WIDTH - 1),
		27880 => to_unsigned(14800, LUT_AMPL_WIDTH - 1),
		27881 => to_unsigned(14797, LUT_AMPL_WIDTH - 1),
		27882 => to_unsigned(14794, LUT_AMPL_WIDTH - 1),
		27883 => to_unsigned(14791, LUT_AMPL_WIDTH - 1),
		27884 => to_unsigned(14789, LUT_AMPL_WIDTH - 1),
		27885 => to_unsigned(14786, LUT_AMPL_WIDTH - 1),
		27886 => to_unsigned(14783, LUT_AMPL_WIDTH - 1),
		27887 => to_unsigned(14780, LUT_AMPL_WIDTH - 1),
		27888 => to_unsigned(14777, LUT_AMPL_WIDTH - 1),
		27889 => to_unsigned(14774, LUT_AMPL_WIDTH - 1),
		27890 => to_unsigned(14772, LUT_AMPL_WIDTH - 1),
		27891 => to_unsigned(14769, LUT_AMPL_WIDTH - 1),
		27892 => to_unsigned(14766, LUT_AMPL_WIDTH - 1),
		27893 => to_unsigned(14763, LUT_AMPL_WIDTH - 1),
		27894 => to_unsigned(14760, LUT_AMPL_WIDTH - 1),
		27895 => to_unsigned(14758, LUT_AMPL_WIDTH - 1),
		27896 => to_unsigned(14755, LUT_AMPL_WIDTH - 1),
		27897 => to_unsigned(14752, LUT_AMPL_WIDTH - 1),
		27898 => to_unsigned(14749, LUT_AMPL_WIDTH - 1),
		27899 => to_unsigned(14746, LUT_AMPL_WIDTH - 1),
		27900 => to_unsigned(14744, LUT_AMPL_WIDTH - 1),
		27901 => to_unsigned(14741, LUT_AMPL_WIDTH - 1),
		27902 => to_unsigned(14738, LUT_AMPL_WIDTH - 1),
		27903 => to_unsigned(14735, LUT_AMPL_WIDTH - 1),
		27904 => to_unsigned(14732, LUT_AMPL_WIDTH - 1),
		27905 => to_unsigned(14730, LUT_AMPL_WIDTH - 1),
		27906 => to_unsigned(14727, LUT_AMPL_WIDTH - 1),
		27907 => to_unsigned(14724, LUT_AMPL_WIDTH - 1),
		27908 => to_unsigned(14721, LUT_AMPL_WIDTH - 1),
		27909 => to_unsigned(14718, LUT_AMPL_WIDTH - 1),
		27910 => to_unsigned(14716, LUT_AMPL_WIDTH - 1),
		27911 => to_unsigned(14713, LUT_AMPL_WIDTH - 1),
		27912 => to_unsigned(14710, LUT_AMPL_WIDTH - 1),
		27913 => to_unsigned(14707, LUT_AMPL_WIDTH - 1),
		27914 => to_unsigned(14704, LUT_AMPL_WIDTH - 1),
		27915 => to_unsigned(14702, LUT_AMPL_WIDTH - 1),
		27916 => to_unsigned(14699, LUT_AMPL_WIDTH - 1),
		27917 => to_unsigned(14696, LUT_AMPL_WIDTH - 1),
		27918 => to_unsigned(14693, LUT_AMPL_WIDTH - 1),
		27919 => to_unsigned(14690, LUT_AMPL_WIDTH - 1),
		27920 => to_unsigned(14688, LUT_AMPL_WIDTH - 1),
		27921 => to_unsigned(14685, LUT_AMPL_WIDTH - 1),
		27922 => to_unsigned(14682, LUT_AMPL_WIDTH - 1),
		27923 => to_unsigned(14679, LUT_AMPL_WIDTH - 1),
		27924 => to_unsigned(14676, LUT_AMPL_WIDTH - 1),
		27925 => to_unsigned(14673, LUT_AMPL_WIDTH - 1),
		27926 => to_unsigned(14671, LUT_AMPL_WIDTH - 1),
		27927 => to_unsigned(14668, LUT_AMPL_WIDTH - 1),
		27928 => to_unsigned(14665, LUT_AMPL_WIDTH - 1),
		27929 => to_unsigned(14662, LUT_AMPL_WIDTH - 1),
		27930 => to_unsigned(14659, LUT_AMPL_WIDTH - 1),
		27931 => to_unsigned(14657, LUT_AMPL_WIDTH - 1),
		27932 => to_unsigned(14654, LUT_AMPL_WIDTH - 1),
		27933 => to_unsigned(14651, LUT_AMPL_WIDTH - 1),
		27934 => to_unsigned(14648, LUT_AMPL_WIDTH - 1),
		27935 => to_unsigned(14645, LUT_AMPL_WIDTH - 1),
		27936 => to_unsigned(14643, LUT_AMPL_WIDTH - 1),
		27937 => to_unsigned(14640, LUT_AMPL_WIDTH - 1),
		27938 => to_unsigned(14637, LUT_AMPL_WIDTH - 1),
		27939 => to_unsigned(14634, LUT_AMPL_WIDTH - 1),
		27940 => to_unsigned(14631, LUT_AMPL_WIDTH - 1),
		27941 => to_unsigned(14628, LUT_AMPL_WIDTH - 1),
		27942 => to_unsigned(14626, LUT_AMPL_WIDTH - 1),
		27943 => to_unsigned(14623, LUT_AMPL_WIDTH - 1),
		27944 => to_unsigned(14620, LUT_AMPL_WIDTH - 1),
		27945 => to_unsigned(14617, LUT_AMPL_WIDTH - 1),
		27946 => to_unsigned(14614, LUT_AMPL_WIDTH - 1),
		27947 => to_unsigned(14612, LUT_AMPL_WIDTH - 1),
		27948 => to_unsigned(14609, LUT_AMPL_WIDTH - 1),
		27949 => to_unsigned(14606, LUT_AMPL_WIDTH - 1),
		27950 => to_unsigned(14603, LUT_AMPL_WIDTH - 1),
		27951 => to_unsigned(14600, LUT_AMPL_WIDTH - 1),
		27952 => to_unsigned(14598, LUT_AMPL_WIDTH - 1),
		27953 => to_unsigned(14595, LUT_AMPL_WIDTH - 1),
		27954 => to_unsigned(14592, LUT_AMPL_WIDTH - 1),
		27955 => to_unsigned(14589, LUT_AMPL_WIDTH - 1),
		27956 => to_unsigned(14586, LUT_AMPL_WIDTH - 1),
		27957 => to_unsigned(14584, LUT_AMPL_WIDTH - 1),
		27958 => to_unsigned(14581, LUT_AMPL_WIDTH - 1),
		27959 => to_unsigned(14578, LUT_AMPL_WIDTH - 1),
		27960 => to_unsigned(14575, LUT_AMPL_WIDTH - 1),
		27961 => to_unsigned(14572, LUT_AMPL_WIDTH - 1),
		27962 => to_unsigned(14569, LUT_AMPL_WIDTH - 1),
		27963 => to_unsigned(14567, LUT_AMPL_WIDTH - 1),
		27964 => to_unsigned(14564, LUT_AMPL_WIDTH - 1),
		27965 => to_unsigned(14561, LUT_AMPL_WIDTH - 1),
		27966 => to_unsigned(14558, LUT_AMPL_WIDTH - 1),
		27967 => to_unsigned(14555, LUT_AMPL_WIDTH - 1),
		27968 => to_unsigned(14553, LUT_AMPL_WIDTH - 1),
		27969 => to_unsigned(14550, LUT_AMPL_WIDTH - 1),
		27970 => to_unsigned(14547, LUT_AMPL_WIDTH - 1),
		27971 => to_unsigned(14544, LUT_AMPL_WIDTH - 1),
		27972 => to_unsigned(14541, LUT_AMPL_WIDTH - 1),
		27973 => to_unsigned(14538, LUT_AMPL_WIDTH - 1),
		27974 => to_unsigned(14536, LUT_AMPL_WIDTH - 1),
		27975 => to_unsigned(14533, LUT_AMPL_WIDTH - 1),
		27976 => to_unsigned(14530, LUT_AMPL_WIDTH - 1),
		27977 => to_unsigned(14527, LUT_AMPL_WIDTH - 1),
		27978 => to_unsigned(14524, LUT_AMPL_WIDTH - 1),
		27979 => to_unsigned(14522, LUT_AMPL_WIDTH - 1),
		27980 => to_unsigned(14519, LUT_AMPL_WIDTH - 1),
		27981 => to_unsigned(14516, LUT_AMPL_WIDTH - 1),
		27982 => to_unsigned(14513, LUT_AMPL_WIDTH - 1),
		27983 => to_unsigned(14510, LUT_AMPL_WIDTH - 1),
		27984 => to_unsigned(14507, LUT_AMPL_WIDTH - 1),
		27985 => to_unsigned(14505, LUT_AMPL_WIDTH - 1),
		27986 => to_unsigned(14502, LUT_AMPL_WIDTH - 1),
		27987 => to_unsigned(14499, LUT_AMPL_WIDTH - 1),
		27988 => to_unsigned(14496, LUT_AMPL_WIDTH - 1),
		27989 => to_unsigned(14493, LUT_AMPL_WIDTH - 1),
		27990 => to_unsigned(14491, LUT_AMPL_WIDTH - 1),
		27991 => to_unsigned(14488, LUT_AMPL_WIDTH - 1),
		27992 => to_unsigned(14485, LUT_AMPL_WIDTH - 1),
		27993 => to_unsigned(14482, LUT_AMPL_WIDTH - 1),
		27994 => to_unsigned(14479, LUT_AMPL_WIDTH - 1),
		27995 => to_unsigned(14477, LUT_AMPL_WIDTH - 1),
		27996 => to_unsigned(14474, LUT_AMPL_WIDTH - 1),
		27997 => to_unsigned(14471, LUT_AMPL_WIDTH - 1),
		27998 => to_unsigned(14468, LUT_AMPL_WIDTH - 1),
		27999 => to_unsigned(14465, LUT_AMPL_WIDTH - 1),
		28000 => to_unsigned(14462, LUT_AMPL_WIDTH - 1),
		28001 => to_unsigned(14460, LUT_AMPL_WIDTH - 1),
		28002 => to_unsigned(14457, LUT_AMPL_WIDTH - 1),
		28003 => to_unsigned(14454, LUT_AMPL_WIDTH - 1),
		28004 => to_unsigned(14451, LUT_AMPL_WIDTH - 1),
		28005 => to_unsigned(14448, LUT_AMPL_WIDTH - 1),
		28006 => to_unsigned(14445, LUT_AMPL_WIDTH - 1),
		28007 => to_unsigned(14443, LUT_AMPL_WIDTH - 1),
		28008 => to_unsigned(14440, LUT_AMPL_WIDTH - 1),
		28009 => to_unsigned(14437, LUT_AMPL_WIDTH - 1),
		28010 => to_unsigned(14434, LUT_AMPL_WIDTH - 1),
		28011 => to_unsigned(14431, LUT_AMPL_WIDTH - 1),
		28012 => to_unsigned(14429, LUT_AMPL_WIDTH - 1),
		28013 => to_unsigned(14426, LUT_AMPL_WIDTH - 1),
		28014 => to_unsigned(14423, LUT_AMPL_WIDTH - 1),
		28015 => to_unsigned(14420, LUT_AMPL_WIDTH - 1),
		28016 => to_unsigned(14417, LUT_AMPL_WIDTH - 1),
		28017 => to_unsigned(14414, LUT_AMPL_WIDTH - 1),
		28018 => to_unsigned(14412, LUT_AMPL_WIDTH - 1),
		28019 => to_unsigned(14409, LUT_AMPL_WIDTH - 1),
		28020 => to_unsigned(14406, LUT_AMPL_WIDTH - 1),
		28021 => to_unsigned(14403, LUT_AMPL_WIDTH - 1),
		28022 => to_unsigned(14400, LUT_AMPL_WIDTH - 1),
		28023 => to_unsigned(14398, LUT_AMPL_WIDTH - 1),
		28024 => to_unsigned(14395, LUT_AMPL_WIDTH - 1),
		28025 => to_unsigned(14392, LUT_AMPL_WIDTH - 1),
		28026 => to_unsigned(14389, LUT_AMPL_WIDTH - 1),
		28027 => to_unsigned(14386, LUT_AMPL_WIDTH - 1),
		28028 => to_unsigned(14383, LUT_AMPL_WIDTH - 1),
		28029 => to_unsigned(14381, LUT_AMPL_WIDTH - 1),
		28030 => to_unsigned(14378, LUT_AMPL_WIDTH - 1),
		28031 => to_unsigned(14375, LUT_AMPL_WIDTH - 1),
		28032 => to_unsigned(14372, LUT_AMPL_WIDTH - 1),
		28033 => to_unsigned(14369, LUT_AMPL_WIDTH - 1),
		28034 => to_unsigned(14366, LUT_AMPL_WIDTH - 1),
		28035 => to_unsigned(14364, LUT_AMPL_WIDTH - 1),
		28036 => to_unsigned(14361, LUT_AMPL_WIDTH - 1),
		28037 => to_unsigned(14358, LUT_AMPL_WIDTH - 1),
		28038 => to_unsigned(14355, LUT_AMPL_WIDTH - 1),
		28039 => to_unsigned(14352, LUT_AMPL_WIDTH - 1),
		28040 => to_unsigned(14350, LUT_AMPL_WIDTH - 1),
		28041 => to_unsigned(14347, LUT_AMPL_WIDTH - 1),
		28042 => to_unsigned(14344, LUT_AMPL_WIDTH - 1),
		28043 => to_unsigned(14341, LUT_AMPL_WIDTH - 1),
		28044 => to_unsigned(14338, LUT_AMPL_WIDTH - 1),
		28045 => to_unsigned(14335, LUT_AMPL_WIDTH - 1),
		28046 => to_unsigned(14333, LUT_AMPL_WIDTH - 1),
		28047 => to_unsigned(14330, LUT_AMPL_WIDTH - 1),
		28048 => to_unsigned(14327, LUT_AMPL_WIDTH - 1),
		28049 => to_unsigned(14324, LUT_AMPL_WIDTH - 1),
		28050 => to_unsigned(14321, LUT_AMPL_WIDTH - 1),
		28051 => to_unsigned(14318, LUT_AMPL_WIDTH - 1),
		28052 => to_unsigned(14316, LUT_AMPL_WIDTH - 1),
		28053 => to_unsigned(14313, LUT_AMPL_WIDTH - 1),
		28054 => to_unsigned(14310, LUT_AMPL_WIDTH - 1),
		28055 => to_unsigned(14307, LUT_AMPL_WIDTH - 1),
		28056 => to_unsigned(14304, LUT_AMPL_WIDTH - 1),
		28057 => to_unsigned(14302, LUT_AMPL_WIDTH - 1),
		28058 => to_unsigned(14299, LUT_AMPL_WIDTH - 1),
		28059 => to_unsigned(14296, LUT_AMPL_WIDTH - 1),
		28060 => to_unsigned(14293, LUT_AMPL_WIDTH - 1),
		28061 => to_unsigned(14290, LUT_AMPL_WIDTH - 1),
		28062 => to_unsigned(14287, LUT_AMPL_WIDTH - 1),
		28063 => to_unsigned(14285, LUT_AMPL_WIDTH - 1),
		28064 => to_unsigned(14282, LUT_AMPL_WIDTH - 1),
		28065 => to_unsigned(14279, LUT_AMPL_WIDTH - 1),
		28066 => to_unsigned(14276, LUT_AMPL_WIDTH - 1),
		28067 => to_unsigned(14273, LUT_AMPL_WIDTH - 1),
		28068 => to_unsigned(14270, LUT_AMPL_WIDTH - 1),
		28069 => to_unsigned(14268, LUT_AMPL_WIDTH - 1),
		28070 => to_unsigned(14265, LUT_AMPL_WIDTH - 1),
		28071 => to_unsigned(14262, LUT_AMPL_WIDTH - 1),
		28072 => to_unsigned(14259, LUT_AMPL_WIDTH - 1),
		28073 => to_unsigned(14256, LUT_AMPL_WIDTH - 1),
		28074 => to_unsigned(14253, LUT_AMPL_WIDTH - 1),
		28075 => to_unsigned(14251, LUT_AMPL_WIDTH - 1),
		28076 => to_unsigned(14248, LUT_AMPL_WIDTH - 1),
		28077 => to_unsigned(14245, LUT_AMPL_WIDTH - 1),
		28078 => to_unsigned(14242, LUT_AMPL_WIDTH - 1),
		28079 => to_unsigned(14239, LUT_AMPL_WIDTH - 1),
		28080 => to_unsigned(14236, LUT_AMPL_WIDTH - 1),
		28081 => to_unsigned(14234, LUT_AMPL_WIDTH - 1),
		28082 => to_unsigned(14231, LUT_AMPL_WIDTH - 1),
		28083 => to_unsigned(14228, LUT_AMPL_WIDTH - 1),
		28084 => to_unsigned(14225, LUT_AMPL_WIDTH - 1),
		28085 => to_unsigned(14222, LUT_AMPL_WIDTH - 1),
		28086 => to_unsigned(14219, LUT_AMPL_WIDTH - 1),
		28087 => to_unsigned(14217, LUT_AMPL_WIDTH - 1),
		28088 => to_unsigned(14214, LUT_AMPL_WIDTH - 1),
		28089 => to_unsigned(14211, LUT_AMPL_WIDTH - 1),
		28090 => to_unsigned(14208, LUT_AMPL_WIDTH - 1),
		28091 => to_unsigned(14205, LUT_AMPL_WIDTH - 1),
		28092 => to_unsigned(14203, LUT_AMPL_WIDTH - 1),
		28093 => to_unsigned(14200, LUT_AMPL_WIDTH - 1),
		28094 => to_unsigned(14197, LUT_AMPL_WIDTH - 1),
		28095 => to_unsigned(14194, LUT_AMPL_WIDTH - 1),
		28096 => to_unsigned(14191, LUT_AMPL_WIDTH - 1),
		28097 => to_unsigned(14188, LUT_AMPL_WIDTH - 1),
		28098 => to_unsigned(14186, LUT_AMPL_WIDTH - 1),
		28099 => to_unsigned(14183, LUT_AMPL_WIDTH - 1),
		28100 => to_unsigned(14180, LUT_AMPL_WIDTH - 1),
		28101 => to_unsigned(14177, LUT_AMPL_WIDTH - 1),
		28102 => to_unsigned(14174, LUT_AMPL_WIDTH - 1),
		28103 => to_unsigned(14171, LUT_AMPL_WIDTH - 1),
		28104 => to_unsigned(14169, LUT_AMPL_WIDTH - 1),
		28105 => to_unsigned(14166, LUT_AMPL_WIDTH - 1),
		28106 => to_unsigned(14163, LUT_AMPL_WIDTH - 1),
		28107 => to_unsigned(14160, LUT_AMPL_WIDTH - 1),
		28108 => to_unsigned(14157, LUT_AMPL_WIDTH - 1),
		28109 => to_unsigned(14154, LUT_AMPL_WIDTH - 1),
		28110 => to_unsigned(14152, LUT_AMPL_WIDTH - 1),
		28111 => to_unsigned(14149, LUT_AMPL_WIDTH - 1),
		28112 => to_unsigned(14146, LUT_AMPL_WIDTH - 1),
		28113 => to_unsigned(14143, LUT_AMPL_WIDTH - 1),
		28114 => to_unsigned(14140, LUT_AMPL_WIDTH - 1),
		28115 => to_unsigned(14137, LUT_AMPL_WIDTH - 1),
		28116 => to_unsigned(14135, LUT_AMPL_WIDTH - 1),
		28117 => to_unsigned(14132, LUT_AMPL_WIDTH - 1),
		28118 => to_unsigned(14129, LUT_AMPL_WIDTH - 1),
		28119 => to_unsigned(14126, LUT_AMPL_WIDTH - 1),
		28120 => to_unsigned(14123, LUT_AMPL_WIDTH - 1),
		28121 => to_unsigned(14120, LUT_AMPL_WIDTH - 1),
		28122 => to_unsigned(14118, LUT_AMPL_WIDTH - 1),
		28123 => to_unsigned(14115, LUT_AMPL_WIDTH - 1),
		28124 => to_unsigned(14112, LUT_AMPL_WIDTH - 1),
		28125 => to_unsigned(14109, LUT_AMPL_WIDTH - 1),
		28126 => to_unsigned(14106, LUT_AMPL_WIDTH - 1),
		28127 => to_unsigned(14103, LUT_AMPL_WIDTH - 1),
		28128 => to_unsigned(14101, LUT_AMPL_WIDTH - 1),
		28129 => to_unsigned(14098, LUT_AMPL_WIDTH - 1),
		28130 => to_unsigned(14095, LUT_AMPL_WIDTH - 1),
		28131 => to_unsigned(14092, LUT_AMPL_WIDTH - 1),
		28132 => to_unsigned(14089, LUT_AMPL_WIDTH - 1),
		28133 => to_unsigned(14086, LUT_AMPL_WIDTH - 1),
		28134 => to_unsigned(14083, LUT_AMPL_WIDTH - 1),
		28135 => to_unsigned(14081, LUT_AMPL_WIDTH - 1),
		28136 => to_unsigned(14078, LUT_AMPL_WIDTH - 1),
		28137 => to_unsigned(14075, LUT_AMPL_WIDTH - 1),
		28138 => to_unsigned(14072, LUT_AMPL_WIDTH - 1),
		28139 => to_unsigned(14069, LUT_AMPL_WIDTH - 1),
		28140 => to_unsigned(14066, LUT_AMPL_WIDTH - 1),
		28141 => to_unsigned(14064, LUT_AMPL_WIDTH - 1),
		28142 => to_unsigned(14061, LUT_AMPL_WIDTH - 1),
		28143 => to_unsigned(14058, LUT_AMPL_WIDTH - 1),
		28144 => to_unsigned(14055, LUT_AMPL_WIDTH - 1),
		28145 => to_unsigned(14052, LUT_AMPL_WIDTH - 1),
		28146 => to_unsigned(14049, LUT_AMPL_WIDTH - 1),
		28147 => to_unsigned(14047, LUT_AMPL_WIDTH - 1),
		28148 => to_unsigned(14044, LUT_AMPL_WIDTH - 1),
		28149 => to_unsigned(14041, LUT_AMPL_WIDTH - 1),
		28150 => to_unsigned(14038, LUT_AMPL_WIDTH - 1),
		28151 => to_unsigned(14035, LUT_AMPL_WIDTH - 1),
		28152 => to_unsigned(14032, LUT_AMPL_WIDTH - 1),
		28153 => to_unsigned(14030, LUT_AMPL_WIDTH - 1),
		28154 => to_unsigned(14027, LUT_AMPL_WIDTH - 1),
		28155 => to_unsigned(14024, LUT_AMPL_WIDTH - 1),
		28156 => to_unsigned(14021, LUT_AMPL_WIDTH - 1),
		28157 => to_unsigned(14018, LUT_AMPL_WIDTH - 1),
		28158 => to_unsigned(14015, LUT_AMPL_WIDTH - 1),
		28159 => to_unsigned(14013, LUT_AMPL_WIDTH - 1),
		28160 => to_unsigned(14010, LUT_AMPL_WIDTH - 1),
		28161 => to_unsigned(14007, LUT_AMPL_WIDTH - 1),
		28162 => to_unsigned(14004, LUT_AMPL_WIDTH - 1),
		28163 => to_unsigned(14001, LUT_AMPL_WIDTH - 1),
		28164 => to_unsigned(13998, LUT_AMPL_WIDTH - 1),
		28165 => to_unsigned(13995, LUT_AMPL_WIDTH - 1),
		28166 => to_unsigned(13993, LUT_AMPL_WIDTH - 1),
		28167 => to_unsigned(13990, LUT_AMPL_WIDTH - 1),
		28168 => to_unsigned(13987, LUT_AMPL_WIDTH - 1),
		28169 => to_unsigned(13984, LUT_AMPL_WIDTH - 1),
		28170 => to_unsigned(13981, LUT_AMPL_WIDTH - 1),
		28171 => to_unsigned(13978, LUT_AMPL_WIDTH - 1),
		28172 => to_unsigned(13976, LUT_AMPL_WIDTH - 1),
		28173 => to_unsigned(13973, LUT_AMPL_WIDTH - 1),
		28174 => to_unsigned(13970, LUT_AMPL_WIDTH - 1),
		28175 => to_unsigned(13967, LUT_AMPL_WIDTH - 1),
		28176 => to_unsigned(13964, LUT_AMPL_WIDTH - 1),
		28177 => to_unsigned(13961, LUT_AMPL_WIDTH - 1),
		28178 => to_unsigned(13959, LUT_AMPL_WIDTH - 1),
		28179 => to_unsigned(13956, LUT_AMPL_WIDTH - 1),
		28180 => to_unsigned(13953, LUT_AMPL_WIDTH - 1),
		28181 => to_unsigned(13950, LUT_AMPL_WIDTH - 1),
		28182 => to_unsigned(13947, LUT_AMPL_WIDTH - 1),
		28183 => to_unsigned(13944, LUT_AMPL_WIDTH - 1),
		28184 => to_unsigned(13942, LUT_AMPL_WIDTH - 1),
		28185 => to_unsigned(13939, LUT_AMPL_WIDTH - 1),
		28186 => to_unsigned(13936, LUT_AMPL_WIDTH - 1),
		28187 => to_unsigned(13933, LUT_AMPL_WIDTH - 1),
		28188 => to_unsigned(13930, LUT_AMPL_WIDTH - 1),
		28189 => to_unsigned(13927, LUT_AMPL_WIDTH - 1),
		28190 => to_unsigned(13924, LUT_AMPL_WIDTH - 1),
		28191 => to_unsigned(13922, LUT_AMPL_WIDTH - 1),
		28192 => to_unsigned(13919, LUT_AMPL_WIDTH - 1),
		28193 => to_unsigned(13916, LUT_AMPL_WIDTH - 1),
		28194 => to_unsigned(13913, LUT_AMPL_WIDTH - 1),
		28195 => to_unsigned(13910, LUT_AMPL_WIDTH - 1),
		28196 => to_unsigned(13907, LUT_AMPL_WIDTH - 1),
		28197 => to_unsigned(13905, LUT_AMPL_WIDTH - 1),
		28198 => to_unsigned(13902, LUT_AMPL_WIDTH - 1),
		28199 => to_unsigned(13899, LUT_AMPL_WIDTH - 1),
		28200 => to_unsigned(13896, LUT_AMPL_WIDTH - 1),
		28201 => to_unsigned(13893, LUT_AMPL_WIDTH - 1),
		28202 => to_unsigned(13890, LUT_AMPL_WIDTH - 1),
		28203 => to_unsigned(13887, LUT_AMPL_WIDTH - 1),
		28204 => to_unsigned(13885, LUT_AMPL_WIDTH - 1),
		28205 => to_unsigned(13882, LUT_AMPL_WIDTH - 1),
		28206 => to_unsigned(13879, LUT_AMPL_WIDTH - 1),
		28207 => to_unsigned(13876, LUT_AMPL_WIDTH - 1),
		28208 => to_unsigned(13873, LUT_AMPL_WIDTH - 1),
		28209 => to_unsigned(13870, LUT_AMPL_WIDTH - 1),
		28210 => to_unsigned(13868, LUT_AMPL_WIDTH - 1),
		28211 => to_unsigned(13865, LUT_AMPL_WIDTH - 1),
		28212 => to_unsigned(13862, LUT_AMPL_WIDTH - 1),
		28213 => to_unsigned(13859, LUT_AMPL_WIDTH - 1),
		28214 => to_unsigned(13856, LUT_AMPL_WIDTH - 1),
		28215 => to_unsigned(13853, LUT_AMPL_WIDTH - 1),
		28216 => to_unsigned(13850, LUT_AMPL_WIDTH - 1),
		28217 => to_unsigned(13848, LUT_AMPL_WIDTH - 1),
		28218 => to_unsigned(13845, LUT_AMPL_WIDTH - 1),
		28219 => to_unsigned(13842, LUT_AMPL_WIDTH - 1),
		28220 => to_unsigned(13839, LUT_AMPL_WIDTH - 1),
		28221 => to_unsigned(13836, LUT_AMPL_WIDTH - 1),
		28222 => to_unsigned(13833, LUT_AMPL_WIDTH - 1),
		28223 => to_unsigned(13831, LUT_AMPL_WIDTH - 1),
		28224 => to_unsigned(13828, LUT_AMPL_WIDTH - 1),
		28225 => to_unsigned(13825, LUT_AMPL_WIDTH - 1),
		28226 => to_unsigned(13822, LUT_AMPL_WIDTH - 1),
		28227 => to_unsigned(13819, LUT_AMPL_WIDTH - 1),
		28228 => to_unsigned(13816, LUT_AMPL_WIDTH - 1),
		28229 => to_unsigned(13813, LUT_AMPL_WIDTH - 1),
		28230 => to_unsigned(13811, LUT_AMPL_WIDTH - 1),
		28231 => to_unsigned(13808, LUT_AMPL_WIDTH - 1),
		28232 => to_unsigned(13805, LUT_AMPL_WIDTH - 1),
		28233 => to_unsigned(13802, LUT_AMPL_WIDTH - 1),
		28234 => to_unsigned(13799, LUT_AMPL_WIDTH - 1),
		28235 => to_unsigned(13796, LUT_AMPL_WIDTH - 1),
		28236 => to_unsigned(13793, LUT_AMPL_WIDTH - 1),
		28237 => to_unsigned(13791, LUT_AMPL_WIDTH - 1),
		28238 => to_unsigned(13788, LUT_AMPL_WIDTH - 1),
		28239 => to_unsigned(13785, LUT_AMPL_WIDTH - 1),
		28240 => to_unsigned(13782, LUT_AMPL_WIDTH - 1),
		28241 => to_unsigned(13779, LUT_AMPL_WIDTH - 1),
		28242 => to_unsigned(13776, LUT_AMPL_WIDTH - 1),
		28243 => to_unsigned(13774, LUT_AMPL_WIDTH - 1),
		28244 => to_unsigned(13771, LUT_AMPL_WIDTH - 1),
		28245 => to_unsigned(13768, LUT_AMPL_WIDTH - 1),
		28246 => to_unsigned(13765, LUT_AMPL_WIDTH - 1),
		28247 => to_unsigned(13762, LUT_AMPL_WIDTH - 1),
		28248 => to_unsigned(13759, LUT_AMPL_WIDTH - 1),
		28249 => to_unsigned(13756, LUT_AMPL_WIDTH - 1),
		28250 => to_unsigned(13754, LUT_AMPL_WIDTH - 1),
		28251 => to_unsigned(13751, LUT_AMPL_WIDTH - 1),
		28252 => to_unsigned(13748, LUT_AMPL_WIDTH - 1),
		28253 => to_unsigned(13745, LUT_AMPL_WIDTH - 1),
		28254 => to_unsigned(13742, LUT_AMPL_WIDTH - 1),
		28255 => to_unsigned(13739, LUT_AMPL_WIDTH - 1),
		28256 => to_unsigned(13736, LUT_AMPL_WIDTH - 1),
		28257 => to_unsigned(13734, LUT_AMPL_WIDTH - 1),
		28258 => to_unsigned(13731, LUT_AMPL_WIDTH - 1),
		28259 => to_unsigned(13728, LUT_AMPL_WIDTH - 1),
		28260 => to_unsigned(13725, LUT_AMPL_WIDTH - 1),
		28261 => to_unsigned(13722, LUT_AMPL_WIDTH - 1),
		28262 => to_unsigned(13719, LUT_AMPL_WIDTH - 1),
		28263 => to_unsigned(13717, LUT_AMPL_WIDTH - 1),
		28264 => to_unsigned(13714, LUT_AMPL_WIDTH - 1),
		28265 => to_unsigned(13711, LUT_AMPL_WIDTH - 1),
		28266 => to_unsigned(13708, LUT_AMPL_WIDTH - 1),
		28267 => to_unsigned(13705, LUT_AMPL_WIDTH - 1),
		28268 => to_unsigned(13702, LUT_AMPL_WIDTH - 1),
		28269 => to_unsigned(13699, LUT_AMPL_WIDTH - 1),
		28270 => to_unsigned(13697, LUT_AMPL_WIDTH - 1),
		28271 => to_unsigned(13694, LUT_AMPL_WIDTH - 1),
		28272 => to_unsigned(13691, LUT_AMPL_WIDTH - 1),
		28273 => to_unsigned(13688, LUT_AMPL_WIDTH - 1),
		28274 => to_unsigned(13685, LUT_AMPL_WIDTH - 1),
		28275 => to_unsigned(13682, LUT_AMPL_WIDTH - 1),
		28276 => to_unsigned(13679, LUT_AMPL_WIDTH - 1),
		28277 => to_unsigned(13677, LUT_AMPL_WIDTH - 1),
		28278 => to_unsigned(13674, LUT_AMPL_WIDTH - 1),
		28279 => to_unsigned(13671, LUT_AMPL_WIDTH - 1),
		28280 => to_unsigned(13668, LUT_AMPL_WIDTH - 1),
		28281 => to_unsigned(13665, LUT_AMPL_WIDTH - 1),
		28282 => to_unsigned(13662, LUT_AMPL_WIDTH - 1),
		28283 => to_unsigned(13659, LUT_AMPL_WIDTH - 1),
		28284 => to_unsigned(13657, LUT_AMPL_WIDTH - 1),
		28285 => to_unsigned(13654, LUT_AMPL_WIDTH - 1),
		28286 => to_unsigned(13651, LUT_AMPL_WIDTH - 1),
		28287 => to_unsigned(13648, LUT_AMPL_WIDTH - 1),
		28288 => to_unsigned(13645, LUT_AMPL_WIDTH - 1),
		28289 => to_unsigned(13642, LUT_AMPL_WIDTH - 1),
		28290 => to_unsigned(13639, LUT_AMPL_WIDTH - 1),
		28291 => to_unsigned(13637, LUT_AMPL_WIDTH - 1),
		28292 => to_unsigned(13634, LUT_AMPL_WIDTH - 1),
		28293 => to_unsigned(13631, LUT_AMPL_WIDTH - 1),
		28294 => to_unsigned(13628, LUT_AMPL_WIDTH - 1),
		28295 => to_unsigned(13625, LUT_AMPL_WIDTH - 1),
		28296 => to_unsigned(13622, LUT_AMPL_WIDTH - 1),
		28297 => to_unsigned(13619, LUT_AMPL_WIDTH - 1),
		28298 => to_unsigned(13617, LUT_AMPL_WIDTH - 1),
		28299 => to_unsigned(13614, LUT_AMPL_WIDTH - 1),
		28300 => to_unsigned(13611, LUT_AMPL_WIDTH - 1),
		28301 => to_unsigned(13608, LUT_AMPL_WIDTH - 1),
		28302 => to_unsigned(13605, LUT_AMPL_WIDTH - 1),
		28303 => to_unsigned(13602, LUT_AMPL_WIDTH - 1),
		28304 => to_unsigned(13599, LUT_AMPL_WIDTH - 1),
		28305 => to_unsigned(13597, LUT_AMPL_WIDTH - 1),
		28306 => to_unsigned(13594, LUT_AMPL_WIDTH - 1),
		28307 => to_unsigned(13591, LUT_AMPL_WIDTH - 1),
		28308 => to_unsigned(13588, LUT_AMPL_WIDTH - 1),
		28309 => to_unsigned(13585, LUT_AMPL_WIDTH - 1),
		28310 => to_unsigned(13582, LUT_AMPL_WIDTH - 1),
		28311 => to_unsigned(13579, LUT_AMPL_WIDTH - 1),
		28312 => to_unsigned(13577, LUT_AMPL_WIDTH - 1),
		28313 => to_unsigned(13574, LUT_AMPL_WIDTH - 1),
		28314 => to_unsigned(13571, LUT_AMPL_WIDTH - 1),
		28315 => to_unsigned(13568, LUT_AMPL_WIDTH - 1),
		28316 => to_unsigned(13565, LUT_AMPL_WIDTH - 1),
		28317 => to_unsigned(13562, LUT_AMPL_WIDTH - 1),
		28318 => to_unsigned(13559, LUT_AMPL_WIDTH - 1),
		28319 => to_unsigned(13557, LUT_AMPL_WIDTH - 1),
		28320 => to_unsigned(13554, LUT_AMPL_WIDTH - 1),
		28321 => to_unsigned(13551, LUT_AMPL_WIDTH - 1),
		28322 => to_unsigned(13548, LUT_AMPL_WIDTH - 1),
		28323 => to_unsigned(13545, LUT_AMPL_WIDTH - 1),
		28324 => to_unsigned(13542, LUT_AMPL_WIDTH - 1),
		28325 => to_unsigned(13539, LUT_AMPL_WIDTH - 1),
		28326 => to_unsigned(13537, LUT_AMPL_WIDTH - 1),
		28327 => to_unsigned(13534, LUT_AMPL_WIDTH - 1),
		28328 => to_unsigned(13531, LUT_AMPL_WIDTH - 1),
		28329 => to_unsigned(13528, LUT_AMPL_WIDTH - 1),
		28330 => to_unsigned(13525, LUT_AMPL_WIDTH - 1),
		28331 => to_unsigned(13522, LUT_AMPL_WIDTH - 1),
		28332 => to_unsigned(13519, LUT_AMPL_WIDTH - 1),
		28333 => to_unsigned(13516, LUT_AMPL_WIDTH - 1),
		28334 => to_unsigned(13514, LUT_AMPL_WIDTH - 1),
		28335 => to_unsigned(13511, LUT_AMPL_WIDTH - 1),
		28336 => to_unsigned(13508, LUT_AMPL_WIDTH - 1),
		28337 => to_unsigned(13505, LUT_AMPL_WIDTH - 1),
		28338 => to_unsigned(13502, LUT_AMPL_WIDTH - 1),
		28339 => to_unsigned(13499, LUT_AMPL_WIDTH - 1),
		28340 => to_unsigned(13496, LUT_AMPL_WIDTH - 1),
		28341 => to_unsigned(13494, LUT_AMPL_WIDTH - 1),
		28342 => to_unsigned(13491, LUT_AMPL_WIDTH - 1),
		28343 => to_unsigned(13488, LUT_AMPL_WIDTH - 1),
		28344 => to_unsigned(13485, LUT_AMPL_WIDTH - 1),
		28345 => to_unsigned(13482, LUT_AMPL_WIDTH - 1),
		28346 => to_unsigned(13479, LUT_AMPL_WIDTH - 1),
		28347 => to_unsigned(13476, LUT_AMPL_WIDTH - 1),
		28348 => to_unsigned(13474, LUT_AMPL_WIDTH - 1),
		28349 => to_unsigned(13471, LUT_AMPL_WIDTH - 1),
		28350 => to_unsigned(13468, LUT_AMPL_WIDTH - 1),
		28351 => to_unsigned(13465, LUT_AMPL_WIDTH - 1),
		28352 => to_unsigned(13462, LUT_AMPL_WIDTH - 1),
		28353 => to_unsigned(13459, LUT_AMPL_WIDTH - 1),
		28354 => to_unsigned(13456, LUT_AMPL_WIDTH - 1),
		28355 => to_unsigned(13454, LUT_AMPL_WIDTH - 1),
		28356 => to_unsigned(13451, LUT_AMPL_WIDTH - 1),
		28357 => to_unsigned(13448, LUT_AMPL_WIDTH - 1),
		28358 => to_unsigned(13445, LUT_AMPL_WIDTH - 1),
		28359 => to_unsigned(13442, LUT_AMPL_WIDTH - 1),
		28360 => to_unsigned(13439, LUT_AMPL_WIDTH - 1),
		28361 => to_unsigned(13436, LUT_AMPL_WIDTH - 1),
		28362 => to_unsigned(13433, LUT_AMPL_WIDTH - 1),
		28363 => to_unsigned(13431, LUT_AMPL_WIDTH - 1),
		28364 => to_unsigned(13428, LUT_AMPL_WIDTH - 1),
		28365 => to_unsigned(13425, LUT_AMPL_WIDTH - 1),
		28366 => to_unsigned(13422, LUT_AMPL_WIDTH - 1),
		28367 => to_unsigned(13419, LUT_AMPL_WIDTH - 1),
		28368 => to_unsigned(13416, LUT_AMPL_WIDTH - 1),
		28369 => to_unsigned(13413, LUT_AMPL_WIDTH - 1),
		28370 => to_unsigned(13411, LUT_AMPL_WIDTH - 1),
		28371 => to_unsigned(13408, LUT_AMPL_WIDTH - 1),
		28372 => to_unsigned(13405, LUT_AMPL_WIDTH - 1),
		28373 => to_unsigned(13402, LUT_AMPL_WIDTH - 1),
		28374 => to_unsigned(13399, LUT_AMPL_WIDTH - 1),
		28375 => to_unsigned(13396, LUT_AMPL_WIDTH - 1),
		28376 => to_unsigned(13393, LUT_AMPL_WIDTH - 1),
		28377 => to_unsigned(13390, LUT_AMPL_WIDTH - 1),
		28378 => to_unsigned(13388, LUT_AMPL_WIDTH - 1),
		28379 => to_unsigned(13385, LUT_AMPL_WIDTH - 1),
		28380 => to_unsigned(13382, LUT_AMPL_WIDTH - 1),
		28381 => to_unsigned(13379, LUT_AMPL_WIDTH - 1),
		28382 => to_unsigned(13376, LUT_AMPL_WIDTH - 1),
		28383 => to_unsigned(13373, LUT_AMPL_WIDTH - 1),
		28384 => to_unsigned(13370, LUT_AMPL_WIDTH - 1),
		28385 => to_unsigned(13368, LUT_AMPL_WIDTH - 1),
		28386 => to_unsigned(13365, LUT_AMPL_WIDTH - 1),
		28387 => to_unsigned(13362, LUT_AMPL_WIDTH - 1),
		28388 => to_unsigned(13359, LUT_AMPL_WIDTH - 1),
		28389 => to_unsigned(13356, LUT_AMPL_WIDTH - 1),
		28390 => to_unsigned(13353, LUT_AMPL_WIDTH - 1),
		28391 => to_unsigned(13350, LUT_AMPL_WIDTH - 1),
		28392 => to_unsigned(13347, LUT_AMPL_WIDTH - 1),
		28393 => to_unsigned(13345, LUT_AMPL_WIDTH - 1),
		28394 => to_unsigned(13342, LUT_AMPL_WIDTH - 1),
		28395 => to_unsigned(13339, LUT_AMPL_WIDTH - 1),
		28396 => to_unsigned(13336, LUT_AMPL_WIDTH - 1),
		28397 => to_unsigned(13333, LUT_AMPL_WIDTH - 1),
		28398 => to_unsigned(13330, LUT_AMPL_WIDTH - 1),
		28399 => to_unsigned(13327, LUT_AMPL_WIDTH - 1),
		28400 => to_unsigned(13324, LUT_AMPL_WIDTH - 1),
		28401 => to_unsigned(13322, LUT_AMPL_WIDTH - 1),
		28402 => to_unsigned(13319, LUT_AMPL_WIDTH - 1),
		28403 => to_unsigned(13316, LUT_AMPL_WIDTH - 1),
		28404 => to_unsigned(13313, LUT_AMPL_WIDTH - 1),
		28405 => to_unsigned(13310, LUT_AMPL_WIDTH - 1),
		28406 => to_unsigned(13307, LUT_AMPL_WIDTH - 1),
		28407 => to_unsigned(13304, LUT_AMPL_WIDTH - 1),
		28408 => to_unsigned(13302, LUT_AMPL_WIDTH - 1),
		28409 => to_unsigned(13299, LUT_AMPL_WIDTH - 1),
		28410 => to_unsigned(13296, LUT_AMPL_WIDTH - 1),
		28411 => to_unsigned(13293, LUT_AMPL_WIDTH - 1),
		28412 => to_unsigned(13290, LUT_AMPL_WIDTH - 1),
		28413 => to_unsigned(13287, LUT_AMPL_WIDTH - 1),
		28414 => to_unsigned(13284, LUT_AMPL_WIDTH - 1),
		28415 => to_unsigned(13281, LUT_AMPL_WIDTH - 1),
		28416 => to_unsigned(13279, LUT_AMPL_WIDTH - 1),
		28417 => to_unsigned(13276, LUT_AMPL_WIDTH - 1),
		28418 => to_unsigned(13273, LUT_AMPL_WIDTH - 1),
		28419 => to_unsigned(13270, LUT_AMPL_WIDTH - 1),
		28420 => to_unsigned(13267, LUT_AMPL_WIDTH - 1),
		28421 => to_unsigned(13264, LUT_AMPL_WIDTH - 1),
		28422 => to_unsigned(13261, LUT_AMPL_WIDTH - 1),
		28423 => to_unsigned(13258, LUT_AMPL_WIDTH - 1),
		28424 => to_unsigned(13256, LUT_AMPL_WIDTH - 1),
		28425 => to_unsigned(13253, LUT_AMPL_WIDTH - 1),
		28426 => to_unsigned(13250, LUT_AMPL_WIDTH - 1),
		28427 => to_unsigned(13247, LUT_AMPL_WIDTH - 1),
		28428 => to_unsigned(13244, LUT_AMPL_WIDTH - 1),
		28429 => to_unsigned(13241, LUT_AMPL_WIDTH - 1),
		28430 => to_unsigned(13238, LUT_AMPL_WIDTH - 1),
		28431 => to_unsigned(13235, LUT_AMPL_WIDTH - 1),
		28432 => to_unsigned(13233, LUT_AMPL_WIDTH - 1),
		28433 => to_unsigned(13230, LUT_AMPL_WIDTH - 1),
		28434 => to_unsigned(13227, LUT_AMPL_WIDTH - 1),
		28435 => to_unsigned(13224, LUT_AMPL_WIDTH - 1),
		28436 => to_unsigned(13221, LUT_AMPL_WIDTH - 1),
		28437 => to_unsigned(13218, LUT_AMPL_WIDTH - 1),
		28438 => to_unsigned(13215, LUT_AMPL_WIDTH - 1),
		28439 => to_unsigned(13212, LUT_AMPL_WIDTH - 1),
		28440 => to_unsigned(13210, LUT_AMPL_WIDTH - 1),
		28441 => to_unsigned(13207, LUT_AMPL_WIDTH - 1),
		28442 => to_unsigned(13204, LUT_AMPL_WIDTH - 1),
		28443 => to_unsigned(13201, LUT_AMPL_WIDTH - 1),
		28444 => to_unsigned(13198, LUT_AMPL_WIDTH - 1),
		28445 => to_unsigned(13195, LUT_AMPL_WIDTH - 1),
		28446 => to_unsigned(13192, LUT_AMPL_WIDTH - 1),
		28447 => to_unsigned(13189, LUT_AMPL_WIDTH - 1),
		28448 => to_unsigned(13187, LUT_AMPL_WIDTH - 1),
		28449 => to_unsigned(13184, LUT_AMPL_WIDTH - 1),
		28450 => to_unsigned(13181, LUT_AMPL_WIDTH - 1),
		28451 => to_unsigned(13178, LUT_AMPL_WIDTH - 1),
		28452 => to_unsigned(13175, LUT_AMPL_WIDTH - 1),
		28453 => to_unsigned(13172, LUT_AMPL_WIDTH - 1),
		28454 => to_unsigned(13169, LUT_AMPL_WIDTH - 1),
		28455 => to_unsigned(13166, LUT_AMPL_WIDTH - 1),
		28456 => to_unsigned(13164, LUT_AMPL_WIDTH - 1),
		28457 => to_unsigned(13161, LUT_AMPL_WIDTH - 1),
		28458 => to_unsigned(13158, LUT_AMPL_WIDTH - 1),
		28459 => to_unsigned(13155, LUT_AMPL_WIDTH - 1),
		28460 => to_unsigned(13152, LUT_AMPL_WIDTH - 1),
		28461 => to_unsigned(13149, LUT_AMPL_WIDTH - 1),
		28462 => to_unsigned(13146, LUT_AMPL_WIDTH - 1),
		28463 => to_unsigned(13143, LUT_AMPL_WIDTH - 1),
		28464 => to_unsigned(13141, LUT_AMPL_WIDTH - 1),
		28465 => to_unsigned(13138, LUT_AMPL_WIDTH - 1),
		28466 => to_unsigned(13135, LUT_AMPL_WIDTH - 1),
		28467 => to_unsigned(13132, LUT_AMPL_WIDTH - 1),
		28468 => to_unsigned(13129, LUT_AMPL_WIDTH - 1),
		28469 => to_unsigned(13126, LUT_AMPL_WIDTH - 1),
		28470 => to_unsigned(13123, LUT_AMPL_WIDTH - 1),
		28471 => to_unsigned(13120, LUT_AMPL_WIDTH - 1),
		28472 => to_unsigned(13118, LUT_AMPL_WIDTH - 1),
		28473 => to_unsigned(13115, LUT_AMPL_WIDTH - 1),
		28474 => to_unsigned(13112, LUT_AMPL_WIDTH - 1),
		28475 => to_unsigned(13109, LUT_AMPL_WIDTH - 1),
		28476 => to_unsigned(13106, LUT_AMPL_WIDTH - 1),
		28477 => to_unsigned(13103, LUT_AMPL_WIDTH - 1),
		28478 => to_unsigned(13100, LUT_AMPL_WIDTH - 1),
		28479 => to_unsigned(13097, LUT_AMPL_WIDTH - 1),
		28480 => to_unsigned(13094, LUT_AMPL_WIDTH - 1),
		28481 => to_unsigned(13092, LUT_AMPL_WIDTH - 1),
		28482 => to_unsigned(13089, LUT_AMPL_WIDTH - 1),
		28483 => to_unsigned(13086, LUT_AMPL_WIDTH - 1),
		28484 => to_unsigned(13083, LUT_AMPL_WIDTH - 1),
		28485 => to_unsigned(13080, LUT_AMPL_WIDTH - 1),
		28486 => to_unsigned(13077, LUT_AMPL_WIDTH - 1),
		28487 => to_unsigned(13074, LUT_AMPL_WIDTH - 1),
		28488 => to_unsigned(13071, LUT_AMPL_WIDTH - 1),
		28489 => to_unsigned(13069, LUT_AMPL_WIDTH - 1),
		28490 => to_unsigned(13066, LUT_AMPL_WIDTH - 1),
		28491 => to_unsigned(13063, LUT_AMPL_WIDTH - 1),
		28492 => to_unsigned(13060, LUT_AMPL_WIDTH - 1),
		28493 => to_unsigned(13057, LUT_AMPL_WIDTH - 1),
		28494 => to_unsigned(13054, LUT_AMPL_WIDTH - 1),
		28495 => to_unsigned(13051, LUT_AMPL_WIDTH - 1),
		28496 => to_unsigned(13048, LUT_AMPL_WIDTH - 1),
		28497 => to_unsigned(13046, LUT_AMPL_WIDTH - 1),
		28498 => to_unsigned(13043, LUT_AMPL_WIDTH - 1),
		28499 => to_unsigned(13040, LUT_AMPL_WIDTH - 1),
		28500 => to_unsigned(13037, LUT_AMPL_WIDTH - 1),
		28501 => to_unsigned(13034, LUT_AMPL_WIDTH - 1),
		28502 => to_unsigned(13031, LUT_AMPL_WIDTH - 1),
		28503 => to_unsigned(13028, LUT_AMPL_WIDTH - 1),
		28504 => to_unsigned(13025, LUT_AMPL_WIDTH - 1),
		28505 => to_unsigned(13022, LUT_AMPL_WIDTH - 1),
		28506 => to_unsigned(13020, LUT_AMPL_WIDTH - 1),
		28507 => to_unsigned(13017, LUT_AMPL_WIDTH - 1),
		28508 => to_unsigned(13014, LUT_AMPL_WIDTH - 1),
		28509 => to_unsigned(13011, LUT_AMPL_WIDTH - 1),
		28510 => to_unsigned(13008, LUT_AMPL_WIDTH - 1),
		28511 => to_unsigned(13005, LUT_AMPL_WIDTH - 1),
		28512 => to_unsigned(13002, LUT_AMPL_WIDTH - 1),
		28513 => to_unsigned(12999, LUT_AMPL_WIDTH - 1),
		28514 => to_unsigned(12997, LUT_AMPL_WIDTH - 1),
		28515 => to_unsigned(12994, LUT_AMPL_WIDTH - 1),
		28516 => to_unsigned(12991, LUT_AMPL_WIDTH - 1),
		28517 => to_unsigned(12988, LUT_AMPL_WIDTH - 1),
		28518 => to_unsigned(12985, LUT_AMPL_WIDTH - 1),
		28519 => to_unsigned(12982, LUT_AMPL_WIDTH - 1),
		28520 => to_unsigned(12979, LUT_AMPL_WIDTH - 1),
		28521 => to_unsigned(12976, LUT_AMPL_WIDTH - 1),
		28522 => to_unsigned(12973, LUT_AMPL_WIDTH - 1),
		28523 => to_unsigned(12971, LUT_AMPL_WIDTH - 1),
		28524 => to_unsigned(12968, LUT_AMPL_WIDTH - 1),
		28525 => to_unsigned(12965, LUT_AMPL_WIDTH - 1),
		28526 => to_unsigned(12962, LUT_AMPL_WIDTH - 1),
		28527 => to_unsigned(12959, LUT_AMPL_WIDTH - 1),
		28528 => to_unsigned(12956, LUT_AMPL_WIDTH - 1),
		28529 => to_unsigned(12953, LUT_AMPL_WIDTH - 1),
		28530 => to_unsigned(12950, LUT_AMPL_WIDTH - 1),
		28531 => to_unsigned(12947, LUT_AMPL_WIDTH - 1),
		28532 => to_unsigned(12945, LUT_AMPL_WIDTH - 1),
		28533 => to_unsigned(12942, LUT_AMPL_WIDTH - 1),
		28534 => to_unsigned(12939, LUT_AMPL_WIDTH - 1),
		28535 => to_unsigned(12936, LUT_AMPL_WIDTH - 1),
		28536 => to_unsigned(12933, LUT_AMPL_WIDTH - 1),
		28537 => to_unsigned(12930, LUT_AMPL_WIDTH - 1),
		28538 => to_unsigned(12927, LUT_AMPL_WIDTH - 1),
		28539 => to_unsigned(12924, LUT_AMPL_WIDTH - 1),
		28540 => to_unsigned(12921, LUT_AMPL_WIDTH - 1),
		28541 => to_unsigned(12919, LUT_AMPL_WIDTH - 1),
		28542 => to_unsigned(12916, LUT_AMPL_WIDTH - 1),
		28543 => to_unsigned(12913, LUT_AMPL_WIDTH - 1),
		28544 => to_unsigned(12910, LUT_AMPL_WIDTH - 1),
		28545 => to_unsigned(12907, LUT_AMPL_WIDTH - 1),
		28546 => to_unsigned(12904, LUT_AMPL_WIDTH - 1),
		28547 => to_unsigned(12901, LUT_AMPL_WIDTH - 1),
		28548 => to_unsigned(12898, LUT_AMPL_WIDTH - 1),
		28549 => to_unsigned(12895, LUT_AMPL_WIDTH - 1),
		28550 => to_unsigned(12893, LUT_AMPL_WIDTH - 1),
		28551 => to_unsigned(12890, LUT_AMPL_WIDTH - 1),
		28552 => to_unsigned(12887, LUT_AMPL_WIDTH - 1),
		28553 => to_unsigned(12884, LUT_AMPL_WIDTH - 1),
		28554 => to_unsigned(12881, LUT_AMPL_WIDTH - 1),
		28555 => to_unsigned(12878, LUT_AMPL_WIDTH - 1),
		28556 => to_unsigned(12875, LUT_AMPL_WIDTH - 1),
		28557 => to_unsigned(12872, LUT_AMPL_WIDTH - 1),
		28558 => to_unsigned(12870, LUT_AMPL_WIDTH - 1),
		28559 => to_unsigned(12867, LUT_AMPL_WIDTH - 1),
		28560 => to_unsigned(12864, LUT_AMPL_WIDTH - 1),
		28561 => to_unsigned(12861, LUT_AMPL_WIDTH - 1),
		28562 => to_unsigned(12858, LUT_AMPL_WIDTH - 1),
		28563 => to_unsigned(12855, LUT_AMPL_WIDTH - 1),
		28564 => to_unsigned(12852, LUT_AMPL_WIDTH - 1),
		28565 => to_unsigned(12849, LUT_AMPL_WIDTH - 1),
		28566 => to_unsigned(12846, LUT_AMPL_WIDTH - 1),
		28567 => to_unsigned(12843, LUT_AMPL_WIDTH - 1),
		28568 => to_unsigned(12841, LUT_AMPL_WIDTH - 1),
		28569 => to_unsigned(12838, LUT_AMPL_WIDTH - 1),
		28570 => to_unsigned(12835, LUT_AMPL_WIDTH - 1),
		28571 => to_unsigned(12832, LUT_AMPL_WIDTH - 1),
		28572 => to_unsigned(12829, LUT_AMPL_WIDTH - 1),
		28573 => to_unsigned(12826, LUT_AMPL_WIDTH - 1),
		28574 => to_unsigned(12823, LUT_AMPL_WIDTH - 1),
		28575 => to_unsigned(12820, LUT_AMPL_WIDTH - 1),
		28576 => to_unsigned(12817, LUT_AMPL_WIDTH - 1),
		28577 => to_unsigned(12815, LUT_AMPL_WIDTH - 1),
		28578 => to_unsigned(12812, LUT_AMPL_WIDTH - 1),
		28579 => to_unsigned(12809, LUT_AMPL_WIDTH - 1),
		28580 => to_unsigned(12806, LUT_AMPL_WIDTH - 1),
		28581 => to_unsigned(12803, LUT_AMPL_WIDTH - 1),
		28582 => to_unsigned(12800, LUT_AMPL_WIDTH - 1),
		28583 => to_unsigned(12797, LUT_AMPL_WIDTH - 1),
		28584 => to_unsigned(12794, LUT_AMPL_WIDTH - 1),
		28585 => to_unsigned(12791, LUT_AMPL_WIDTH - 1),
		28586 => to_unsigned(12789, LUT_AMPL_WIDTH - 1),
		28587 => to_unsigned(12786, LUT_AMPL_WIDTH - 1),
		28588 => to_unsigned(12783, LUT_AMPL_WIDTH - 1),
		28589 => to_unsigned(12780, LUT_AMPL_WIDTH - 1),
		28590 => to_unsigned(12777, LUT_AMPL_WIDTH - 1),
		28591 => to_unsigned(12774, LUT_AMPL_WIDTH - 1),
		28592 => to_unsigned(12771, LUT_AMPL_WIDTH - 1),
		28593 => to_unsigned(12768, LUT_AMPL_WIDTH - 1),
		28594 => to_unsigned(12765, LUT_AMPL_WIDTH - 1),
		28595 => to_unsigned(12763, LUT_AMPL_WIDTH - 1),
		28596 => to_unsigned(12760, LUT_AMPL_WIDTH - 1),
		28597 => to_unsigned(12757, LUT_AMPL_WIDTH - 1),
		28598 => to_unsigned(12754, LUT_AMPL_WIDTH - 1),
		28599 => to_unsigned(12751, LUT_AMPL_WIDTH - 1),
		28600 => to_unsigned(12748, LUT_AMPL_WIDTH - 1),
		28601 => to_unsigned(12745, LUT_AMPL_WIDTH - 1),
		28602 => to_unsigned(12742, LUT_AMPL_WIDTH - 1),
		28603 => to_unsigned(12739, LUT_AMPL_WIDTH - 1),
		28604 => to_unsigned(12736, LUT_AMPL_WIDTH - 1),
		28605 => to_unsigned(12734, LUT_AMPL_WIDTH - 1),
		28606 => to_unsigned(12731, LUT_AMPL_WIDTH - 1),
		28607 => to_unsigned(12728, LUT_AMPL_WIDTH - 1),
		28608 => to_unsigned(12725, LUT_AMPL_WIDTH - 1),
		28609 => to_unsigned(12722, LUT_AMPL_WIDTH - 1),
		28610 => to_unsigned(12719, LUT_AMPL_WIDTH - 1),
		28611 => to_unsigned(12716, LUT_AMPL_WIDTH - 1),
		28612 => to_unsigned(12713, LUT_AMPL_WIDTH - 1),
		28613 => to_unsigned(12710, LUT_AMPL_WIDTH - 1),
		28614 => to_unsigned(12708, LUT_AMPL_WIDTH - 1),
		28615 => to_unsigned(12705, LUT_AMPL_WIDTH - 1),
		28616 => to_unsigned(12702, LUT_AMPL_WIDTH - 1),
		28617 => to_unsigned(12699, LUT_AMPL_WIDTH - 1),
		28618 => to_unsigned(12696, LUT_AMPL_WIDTH - 1),
		28619 => to_unsigned(12693, LUT_AMPL_WIDTH - 1),
		28620 => to_unsigned(12690, LUT_AMPL_WIDTH - 1),
		28621 => to_unsigned(12687, LUT_AMPL_WIDTH - 1),
		28622 => to_unsigned(12684, LUT_AMPL_WIDTH - 1),
		28623 => to_unsigned(12681, LUT_AMPL_WIDTH - 1),
		28624 => to_unsigned(12679, LUT_AMPL_WIDTH - 1),
		28625 => to_unsigned(12676, LUT_AMPL_WIDTH - 1),
		28626 => to_unsigned(12673, LUT_AMPL_WIDTH - 1),
		28627 => to_unsigned(12670, LUT_AMPL_WIDTH - 1),
		28628 => to_unsigned(12667, LUT_AMPL_WIDTH - 1),
		28629 => to_unsigned(12664, LUT_AMPL_WIDTH - 1),
		28630 => to_unsigned(12661, LUT_AMPL_WIDTH - 1),
		28631 => to_unsigned(12658, LUT_AMPL_WIDTH - 1),
		28632 => to_unsigned(12655, LUT_AMPL_WIDTH - 1),
		28633 => to_unsigned(12652, LUT_AMPL_WIDTH - 1),
		28634 => to_unsigned(12650, LUT_AMPL_WIDTH - 1),
		28635 => to_unsigned(12647, LUT_AMPL_WIDTH - 1),
		28636 => to_unsigned(12644, LUT_AMPL_WIDTH - 1),
		28637 => to_unsigned(12641, LUT_AMPL_WIDTH - 1),
		28638 => to_unsigned(12638, LUT_AMPL_WIDTH - 1),
		28639 => to_unsigned(12635, LUT_AMPL_WIDTH - 1),
		28640 => to_unsigned(12632, LUT_AMPL_WIDTH - 1),
		28641 => to_unsigned(12629, LUT_AMPL_WIDTH - 1),
		28642 => to_unsigned(12626, LUT_AMPL_WIDTH - 1),
		28643 => to_unsigned(12624, LUT_AMPL_WIDTH - 1),
		28644 => to_unsigned(12621, LUT_AMPL_WIDTH - 1),
		28645 => to_unsigned(12618, LUT_AMPL_WIDTH - 1),
		28646 => to_unsigned(12615, LUT_AMPL_WIDTH - 1),
		28647 => to_unsigned(12612, LUT_AMPL_WIDTH - 1),
		28648 => to_unsigned(12609, LUT_AMPL_WIDTH - 1),
		28649 => to_unsigned(12606, LUT_AMPL_WIDTH - 1),
		28650 => to_unsigned(12603, LUT_AMPL_WIDTH - 1),
		28651 => to_unsigned(12600, LUT_AMPL_WIDTH - 1),
		28652 => to_unsigned(12597, LUT_AMPL_WIDTH - 1),
		28653 => to_unsigned(12595, LUT_AMPL_WIDTH - 1),
		28654 => to_unsigned(12592, LUT_AMPL_WIDTH - 1),
		28655 => to_unsigned(12589, LUT_AMPL_WIDTH - 1),
		28656 => to_unsigned(12586, LUT_AMPL_WIDTH - 1),
		28657 => to_unsigned(12583, LUT_AMPL_WIDTH - 1),
		28658 => to_unsigned(12580, LUT_AMPL_WIDTH - 1),
		28659 => to_unsigned(12577, LUT_AMPL_WIDTH - 1),
		28660 => to_unsigned(12574, LUT_AMPL_WIDTH - 1),
		28661 => to_unsigned(12571, LUT_AMPL_WIDTH - 1),
		28662 => to_unsigned(12568, LUT_AMPL_WIDTH - 1),
		28663 => to_unsigned(12566, LUT_AMPL_WIDTH - 1),
		28664 => to_unsigned(12563, LUT_AMPL_WIDTH - 1),
		28665 => to_unsigned(12560, LUT_AMPL_WIDTH - 1),
		28666 => to_unsigned(12557, LUT_AMPL_WIDTH - 1),
		28667 => to_unsigned(12554, LUT_AMPL_WIDTH - 1),
		28668 => to_unsigned(12551, LUT_AMPL_WIDTH - 1),
		28669 => to_unsigned(12548, LUT_AMPL_WIDTH - 1),
		28670 => to_unsigned(12545, LUT_AMPL_WIDTH - 1),
		28671 => to_unsigned(12542, LUT_AMPL_WIDTH - 1),
		28672 => to_unsigned(12539, LUT_AMPL_WIDTH - 1),
		28673 => to_unsigned(12536, LUT_AMPL_WIDTH - 1),
		28674 => to_unsigned(12534, LUT_AMPL_WIDTH - 1),
		28675 => to_unsigned(12531, LUT_AMPL_WIDTH - 1),
		28676 => to_unsigned(12528, LUT_AMPL_WIDTH - 1),
		28677 => to_unsigned(12525, LUT_AMPL_WIDTH - 1),
		28678 => to_unsigned(12522, LUT_AMPL_WIDTH - 1),
		28679 => to_unsigned(12519, LUT_AMPL_WIDTH - 1),
		28680 => to_unsigned(12516, LUT_AMPL_WIDTH - 1),
		28681 => to_unsigned(12513, LUT_AMPL_WIDTH - 1),
		28682 => to_unsigned(12510, LUT_AMPL_WIDTH - 1),
		28683 => to_unsigned(12507, LUT_AMPL_WIDTH - 1),
		28684 => to_unsigned(12505, LUT_AMPL_WIDTH - 1),
		28685 => to_unsigned(12502, LUT_AMPL_WIDTH - 1),
		28686 => to_unsigned(12499, LUT_AMPL_WIDTH - 1),
		28687 => to_unsigned(12496, LUT_AMPL_WIDTH - 1),
		28688 => to_unsigned(12493, LUT_AMPL_WIDTH - 1),
		28689 => to_unsigned(12490, LUT_AMPL_WIDTH - 1),
		28690 => to_unsigned(12487, LUT_AMPL_WIDTH - 1),
		28691 => to_unsigned(12484, LUT_AMPL_WIDTH - 1),
		28692 => to_unsigned(12481, LUT_AMPL_WIDTH - 1),
		28693 => to_unsigned(12478, LUT_AMPL_WIDTH - 1),
		28694 => to_unsigned(12476, LUT_AMPL_WIDTH - 1),
		28695 => to_unsigned(12473, LUT_AMPL_WIDTH - 1),
		28696 => to_unsigned(12470, LUT_AMPL_WIDTH - 1),
		28697 => to_unsigned(12467, LUT_AMPL_WIDTH - 1),
		28698 => to_unsigned(12464, LUT_AMPL_WIDTH - 1),
		28699 => to_unsigned(12461, LUT_AMPL_WIDTH - 1),
		28700 => to_unsigned(12458, LUT_AMPL_WIDTH - 1),
		28701 => to_unsigned(12455, LUT_AMPL_WIDTH - 1),
		28702 => to_unsigned(12452, LUT_AMPL_WIDTH - 1),
		28703 => to_unsigned(12449, LUT_AMPL_WIDTH - 1),
		28704 => to_unsigned(12446, LUT_AMPL_WIDTH - 1),
		28705 => to_unsigned(12444, LUT_AMPL_WIDTH - 1),
		28706 => to_unsigned(12441, LUT_AMPL_WIDTH - 1),
		28707 => to_unsigned(12438, LUT_AMPL_WIDTH - 1),
		28708 => to_unsigned(12435, LUT_AMPL_WIDTH - 1),
		28709 => to_unsigned(12432, LUT_AMPL_WIDTH - 1),
		28710 => to_unsigned(12429, LUT_AMPL_WIDTH - 1),
		28711 => to_unsigned(12426, LUT_AMPL_WIDTH - 1),
		28712 => to_unsigned(12423, LUT_AMPL_WIDTH - 1),
		28713 => to_unsigned(12420, LUT_AMPL_WIDTH - 1),
		28714 => to_unsigned(12417, LUT_AMPL_WIDTH - 1),
		28715 => to_unsigned(12414, LUT_AMPL_WIDTH - 1),
		28716 => to_unsigned(12412, LUT_AMPL_WIDTH - 1),
		28717 => to_unsigned(12409, LUT_AMPL_WIDTH - 1),
		28718 => to_unsigned(12406, LUT_AMPL_WIDTH - 1),
		28719 => to_unsigned(12403, LUT_AMPL_WIDTH - 1),
		28720 => to_unsigned(12400, LUT_AMPL_WIDTH - 1),
		28721 => to_unsigned(12397, LUT_AMPL_WIDTH - 1),
		28722 => to_unsigned(12394, LUT_AMPL_WIDTH - 1),
		28723 => to_unsigned(12391, LUT_AMPL_WIDTH - 1),
		28724 => to_unsigned(12388, LUT_AMPL_WIDTH - 1),
		28725 => to_unsigned(12385, LUT_AMPL_WIDTH - 1),
		28726 => to_unsigned(12382, LUT_AMPL_WIDTH - 1),
		28727 => to_unsigned(12380, LUT_AMPL_WIDTH - 1),
		28728 => to_unsigned(12377, LUT_AMPL_WIDTH - 1),
		28729 => to_unsigned(12374, LUT_AMPL_WIDTH - 1),
		28730 => to_unsigned(12371, LUT_AMPL_WIDTH - 1),
		28731 => to_unsigned(12368, LUT_AMPL_WIDTH - 1),
		28732 => to_unsigned(12365, LUT_AMPL_WIDTH - 1),
		28733 => to_unsigned(12362, LUT_AMPL_WIDTH - 1),
		28734 => to_unsigned(12359, LUT_AMPL_WIDTH - 1),
		28735 => to_unsigned(12356, LUT_AMPL_WIDTH - 1),
		28736 => to_unsigned(12353, LUT_AMPL_WIDTH - 1),
		28737 => to_unsigned(12350, LUT_AMPL_WIDTH - 1),
		28738 => to_unsigned(12348, LUT_AMPL_WIDTH - 1),
		28739 => to_unsigned(12345, LUT_AMPL_WIDTH - 1),
		28740 => to_unsigned(12342, LUT_AMPL_WIDTH - 1),
		28741 => to_unsigned(12339, LUT_AMPL_WIDTH - 1),
		28742 => to_unsigned(12336, LUT_AMPL_WIDTH - 1),
		28743 => to_unsigned(12333, LUT_AMPL_WIDTH - 1),
		28744 => to_unsigned(12330, LUT_AMPL_WIDTH - 1),
		28745 => to_unsigned(12327, LUT_AMPL_WIDTH - 1),
		28746 => to_unsigned(12324, LUT_AMPL_WIDTH - 1),
		28747 => to_unsigned(12321, LUT_AMPL_WIDTH - 1),
		28748 => to_unsigned(12318, LUT_AMPL_WIDTH - 1),
		28749 => to_unsigned(12316, LUT_AMPL_WIDTH - 1),
		28750 => to_unsigned(12313, LUT_AMPL_WIDTH - 1),
		28751 => to_unsigned(12310, LUT_AMPL_WIDTH - 1),
		28752 => to_unsigned(12307, LUT_AMPL_WIDTH - 1),
		28753 => to_unsigned(12304, LUT_AMPL_WIDTH - 1),
		28754 => to_unsigned(12301, LUT_AMPL_WIDTH - 1),
		28755 => to_unsigned(12298, LUT_AMPL_WIDTH - 1),
		28756 => to_unsigned(12295, LUT_AMPL_WIDTH - 1),
		28757 => to_unsigned(12292, LUT_AMPL_WIDTH - 1),
		28758 => to_unsigned(12289, LUT_AMPL_WIDTH - 1),
		28759 => to_unsigned(12286, LUT_AMPL_WIDTH - 1),
		28760 => to_unsigned(12284, LUT_AMPL_WIDTH - 1),
		28761 => to_unsigned(12281, LUT_AMPL_WIDTH - 1),
		28762 => to_unsigned(12278, LUT_AMPL_WIDTH - 1),
		28763 => to_unsigned(12275, LUT_AMPL_WIDTH - 1),
		28764 => to_unsigned(12272, LUT_AMPL_WIDTH - 1),
		28765 => to_unsigned(12269, LUT_AMPL_WIDTH - 1),
		28766 => to_unsigned(12266, LUT_AMPL_WIDTH - 1),
		28767 => to_unsigned(12263, LUT_AMPL_WIDTH - 1),
		28768 => to_unsigned(12260, LUT_AMPL_WIDTH - 1),
		28769 => to_unsigned(12257, LUT_AMPL_WIDTH - 1),
		28770 => to_unsigned(12254, LUT_AMPL_WIDTH - 1),
		28771 => to_unsigned(12251, LUT_AMPL_WIDTH - 1),
		28772 => to_unsigned(12249, LUT_AMPL_WIDTH - 1),
		28773 => to_unsigned(12246, LUT_AMPL_WIDTH - 1),
		28774 => to_unsigned(12243, LUT_AMPL_WIDTH - 1),
		28775 => to_unsigned(12240, LUT_AMPL_WIDTH - 1),
		28776 => to_unsigned(12237, LUT_AMPL_WIDTH - 1),
		28777 => to_unsigned(12234, LUT_AMPL_WIDTH - 1),
		28778 => to_unsigned(12231, LUT_AMPL_WIDTH - 1),
		28779 => to_unsigned(12228, LUT_AMPL_WIDTH - 1),
		28780 => to_unsigned(12225, LUT_AMPL_WIDTH - 1),
		28781 => to_unsigned(12222, LUT_AMPL_WIDTH - 1),
		28782 => to_unsigned(12219, LUT_AMPL_WIDTH - 1),
		28783 => to_unsigned(12217, LUT_AMPL_WIDTH - 1),
		28784 => to_unsigned(12214, LUT_AMPL_WIDTH - 1),
		28785 => to_unsigned(12211, LUT_AMPL_WIDTH - 1),
		28786 => to_unsigned(12208, LUT_AMPL_WIDTH - 1),
		28787 => to_unsigned(12205, LUT_AMPL_WIDTH - 1),
		28788 => to_unsigned(12202, LUT_AMPL_WIDTH - 1),
		28789 => to_unsigned(12199, LUT_AMPL_WIDTH - 1),
		28790 => to_unsigned(12196, LUT_AMPL_WIDTH - 1),
		28791 => to_unsigned(12193, LUT_AMPL_WIDTH - 1),
		28792 => to_unsigned(12190, LUT_AMPL_WIDTH - 1),
		28793 => to_unsigned(12187, LUT_AMPL_WIDTH - 1),
		28794 => to_unsigned(12184, LUT_AMPL_WIDTH - 1),
		28795 => to_unsigned(12182, LUT_AMPL_WIDTH - 1),
		28796 => to_unsigned(12179, LUT_AMPL_WIDTH - 1),
		28797 => to_unsigned(12176, LUT_AMPL_WIDTH - 1),
		28798 => to_unsigned(12173, LUT_AMPL_WIDTH - 1),
		28799 => to_unsigned(12170, LUT_AMPL_WIDTH - 1),
		28800 => to_unsigned(12167, LUT_AMPL_WIDTH - 1),
		28801 => to_unsigned(12164, LUT_AMPL_WIDTH - 1),
		28802 => to_unsigned(12161, LUT_AMPL_WIDTH - 1),
		28803 => to_unsigned(12158, LUT_AMPL_WIDTH - 1),
		28804 => to_unsigned(12155, LUT_AMPL_WIDTH - 1),
		28805 => to_unsigned(12152, LUT_AMPL_WIDTH - 1),
		28806 => to_unsigned(12149, LUT_AMPL_WIDTH - 1),
		28807 => to_unsigned(12147, LUT_AMPL_WIDTH - 1),
		28808 => to_unsigned(12144, LUT_AMPL_WIDTH - 1),
		28809 => to_unsigned(12141, LUT_AMPL_WIDTH - 1),
		28810 => to_unsigned(12138, LUT_AMPL_WIDTH - 1),
		28811 => to_unsigned(12135, LUT_AMPL_WIDTH - 1),
		28812 => to_unsigned(12132, LUT_AMPL_WIDTH - 1),
		28813 => to_unsigned(12129, LUT_AMPL_WIDTH - 1),
		28814 => to_unsigned(12126, LUT_AMPL_WIDTH - 1),
		28815 => to_unsigned(12123, LUT_AMPL_WIDTH - 1),
		28816 => to_unsigned(12120, LUT_AMPL_WIDTH - 1),
		28817 => to_unsigned(12117, LUT_AMPL_WIDTH - 1),
		28818 => to_unsigned(12114, LUT_AMPL_WIDTH - 1),
		28819 => to_unsigned(12112, LUT_AMPL_WIDTH - 1),
		28820 => to_unsigned(12109, LUT_AMPL_WIDTH - 1),
		28821 => to_unsigned(12106, LUT_AMPL_WIDTH - 1),
		28822 => to_unsigned(12103, LUT_AMPL_WIDTH - 1),
		28823 => to_unsigned(12100, LUT_AMPL_WIDTH - 1),
		28824 => to_unsigned(12097, LUT_AMPL_WIDTH - 1),
		28825 => to_unsigned(12094, LUT_AMPL_WIDTH - 1),
		28826 => to_unsigned(12091, LUT_AMPL_WIDTH - 1),
		28827 => to_unsigned(12088, LUT_AMPL_WIDTH - 1),
		28828 => to_unsigned(12085, LUT_AMPL_WIDTH - 1),
		28829 => to_unsigned(12082, LUT_AMPL_WIDTH - 1),
		28830 => to_unsigned(12079, LUT_AMPL_WIDTH - 1),
		28831 => to_unsigned(12076, LUT_AMPL_WIDTH - 1),
		28832 => to_unsigned(12074, LUT_AMPL_WIDTH - 1),
		28833 => to_unsigned(12071, LUT_AMPL_WIDTH - 1),
		28834 => to_unsigned(12068, LUT_AMPL_WIDTH - 1),
		28835 => to_unsigned(12065, LUT_AMPL_WIDTH - 1),
		28836 => to_unsigned(12062, LUT_AMPL_WIDTH - 1),
		28837 => to_unsigned(12059, LUT_AMPL_WIDTH - 1),
		28838 => to_unsigned(12056, LUT_AMPL_WIDTH - 1),
		28839 => to_unsigned(12053, LUT_AMPL_WIDTH - 1),
		28840 => to_unsigned(12050, LUT_AMPL_WIDTH - 1),
		28841 => to_unsigned(12047, LUT_AMPL_WIDTH - 1),
		28842 => to_unsigned(12044, LUT_AMPL_WIDTH - 1),
		28843 => to_unsigned(12041, LUT_AMPL_WIDTH - 1),
		28844 => to_unsigned(12038, LUT_AMPL_WIDTH - 1),
		28845 => to_unsigned(12036, LUT_AMPL_WIDTH - 1),
		28846 => to_unsigned(12033, LUT_AMPL_WIDTH - 1),
		28847 => to_unsigned(12030, LUT_AMPL_WIDTH - 1),
		28848 => to_unsigned(12027, LUT_AMPL_WIDTH - 1),
		28849 => to_unsigned(12024, LUT_AMPL_WIDTH - 1),
		28850 => to_unsigned(12021, LUT_AMPL_WIDTH - 1),
		28851 => to_unsigned(12018, LUT_AMPL_WIDTH - 1),
		28852 => to_unsigned(12015, LUT_AMPL_WIDTH - 1),
		28853 => to_unsigned(12012, LUT_AMPL_WIDTH - 1),
		28854 => to_unsigned(12009, LUT_AMPL_WIDTH - 1),
		28855 => to_unsigned(12006, LUT_AMPL_WIDTH - 1),
		28856 => to_unsigned(12003, LUT_AMPL_WIDTH - 1),
		28857 => to_unsigned(12001, LUT_AMPL_WIDTH - 1),
		28858 => to_unsigned(11998, LUT_AMPL_WIDTH - 1),
		28859 => to_unsigned(11995, LUT_AMPL_WIDTH - 1),
		28860 => to_unsigned(11992, LUT_AMPL_WIDTH - 1),
		28861 => to_unsigned(11989, LUT_AMPL_WIDTH - 1),
		28862 => to_unsigned(11986, LUT_AMPL_WIDTH - 1),
		28863 => to_unsigned(11983, LUT_AMPL_WIDTH - 1),
		28864 => to_unsigned(11980, LUT_AMPL_WIDTH - 1),
		28865 => to_unsigned(11977, LUT_AMPL_WIDTH - 1),
		28866 => to_unsigned(11974, LUT_AMPL_WIDTH - 1),
		28867 => to_unsigned(11971, LUT_AMPL_WIDTH - 1),
		28868 => to_unsigned(11968, LUT_AMPL_WIDTH - 1),
		28869 => to_unsigned(11965, LUT_AMPL_WIDTH - 1),
		28870 => to_unsigned(11962, LUT_AMPL_WIDTH - 1),
		28871 => to_unsigned(11960, LUT_AMPL_WIDTH - 1),
		28872 => to_unsigned(11957, LUT_AMPL_WIDTH - 1),
		28873 => to_unsigned(11954, LUT_AMPL_WIDTH - 1),
		28874 => to_unsigned(11951, LUT_AMPL_WIDTH - 1),
		28875 => to_unsigned(11948, LUT_AMPL_WIDTH - 1),
		28876 => to_unsigned(11945, LUT_AMPL_WIDTH - 1),
		28877 => to_unsigned(11942, LUT_AMPL_WIDTH - 1),
		28878 => to_unsigned(11939, LUT_AMPL_WIDTH - 1),
		28879 => to_unsigned(11936, LUT_AMPL_WIDTH - 1),
		28880 => to_unsigned(11933, LUT_AMPL_WIDTH - 1),
		28881 => to_unsigned(11930, LUT_AMPL_WIDTH - 1),
		28882 => to_unsigned(11927, LUT_AMPL_WIDTH - 1),
		28883 => to_unsigned(11924, LUT_AMPL_WIDTH - 1),
		28884 => to_unsigned(11922, LUT_AMPL_WIDTH - 1),
		28885 => to_unsigned(11919, LUT_AMPL_WIDTH - 1),
		28886 => to_unsigned(11916, LUT_AMPL_WIDTH - 1),
		28887 => to_unsigned(11913, LUT_AMPL_WIDTH - 1),
		28888 => to_unsigned(11910, LUT_AMPL_WIDTH - 1),
		28889 => to_unsigned(11907, LUT_AMPL_WIDTH - 1),
		28890 => to_unsigned(11904, LUT_AMPL_WIDTH - 1),
		28891 => to_unsigned(11901, LUT_AMPL_WIDTH - 1),
		28892 => to_unsigned(11898, LUT_AMPL_WIDTH - 1),
		28893 => to_unsigned(11895, LUT_AMPL_WIDTH - 1),
		28894 => to_unsigned(11892, LUT_AMPL_WIDTH - 1),
		28895 => to_unsigned(11889, LUT_AMPL_WIDTH - 1),
		28896 => to_unsigned(11886, LUT_AMPL_WIDTH - 1),
		28897 => to_unsigned(11883, LUT_AMPL_WIDTH - 1),
		28898 => to_unsigned(11881, LUT_AMPL_WIDTH - 1),
		28899 => to_unsigned(11878, LUT_AMPL_WIDTH - 1),
		28900 => to_unsigned(11875, LUT_AMPL_WIDTH - 1),
		28901 => to_unsigned(11872, LUT_AMPL_WIDTH - 1),
		28902 => to_unsigned(11869, LUT_AMPL_WIDTH - 1),
		28903 => to_unsigned(11866, LUT_AMPL_WIDTH - 1),
		28904 => to_unsigned(11863, LUT_AMPL_WIDTH - 1),
		28905 => to_unsigned(11860, LUT_AMPL_WIDTH - 1),
		28906 => to_unsigned(11857, LUT_AMPL_WIDTH - 1),
		28907 => to_unsigned(11854, LUT_AMPL_WIDTH - 1),
		28908 => to_unsigned(11851, LUT_AMPL_WIDTH - 1),
		28909 => to_unsigned(11848, LUT_AMPL_WIDTH - 1),
		28910 => to_unsigned(11845, LUT_AMPL_WIDTH - 1),
		28911 => to_unsigned(11842, LUT_AMPL_WIDTH - 1),
		28912 => to_unsigned(11840, LUT_AMPL_WIDTH - 1),
		28913 => to_unsigned(11837, LUT_AMPL_WIDTH - 1),
		28914 => to_unsigned(11834, LUT_AMPL_WIDTH - 1),
		28915 => to_unsigned(11831, LUT_AMPL_WIDTH - 1),
		28916 => to_unsigned(11828, LUT_AMPL_WIDTH - 1),
		28917 => to_unsigned(11825, LUT_AMPL_WIDTH - 1),
		28918 => to_unsigned(11822, LUT_AMPL_WIDTH - 1),
		28919 => to_unsigned(11819, LUT_AMPL_WIDTH - 1),
		28920 => to_unsigned(11816, LUT_AMPL_WIDTH - 1),
		28921 => to_unsigned(11813, LUT_AMPL_WIDTH - 1),
		28922 => to_unsigned(11810, LUT_AMPL_WIDTH - 1),
		28923 => to_unsigned(11807, LUT_AMPL_WIDTH - 1),
		28924 => to_unsigned(11804, LUT_AMPL_WIDTH - 1),
		28925 => to_unsigned(11801, LUT_AMPL_WIDTH - 1),
		28926 => to_unsigned(11799, LUT_AMPL_WIDTH - 1),
		28927 => to_unsigned(11796, LUT_AMPL_WIDTH - 1),
		28928 => to_unsigned(11793, LUT_AMPL_WIDTH - 1),
		28929 => to_unsigned(11790, LUT_AMPL_WIDTH - 1),
		28930 => to_unsigned(11787, LUT_AMPL_WIDTH - 1),
		28931 => to_unsigned(11784, LUT_AMPL_WIDTH - 1),
		28932 => to_unsigned(11781, LUT_AMPL_WIDTH - 1),
		28933 => to_unsigned(11778, LUT_AMPL_WIDTH - 1),
		28934 => to_unsigned(11775, LUT_AMPL_WIDTH - 1),
		28935 => to_unsigned(11772, LUT_AMPL_WIDTH - 1),
		28936 => to_unsigned(11769, LUT_AMPL_WIDTH - 1),
		28937 => to_unsigned(11766, LUT_AMPL_WIDTH - 1),
		28938 => to_unsigned(11763, LUT_AMPL_WIDTH - 1),
		28939 => to_unsigned(11760, LUT_AMPL_WIDTH - 1),
		28940 => to_unsigned(11758, LUT_AMPL_WIDTH - 1),
		28941 => to_unsigned(11755, LUT_AMPL_WIDTH - 1),
		28942 => to_unsigned(11752, LUT_AMPL_WIDTH - 1),
		28943 => to_unsigned(11749, LUT_AMPL_WIDTH - 1),
		28944 => to_unsigned(11746, LUT_AMPL_WIDTH - 1),
		28945 => to_unsigned(11743, LUT_AMPL_WIDTH - 1),
		28946 => to_unsigned(11740, LUT_AMPL_WIDTH - 1),
		28947 => to_unsigned(11737, LUT_AMPL_WIDTH - 1),
		28948 => to_unsigned(11734, LUT_AMPL_WIDTH - 1),
		28949 => to_unsigned(11731, LUT_AMPL_WIDTH - 1),
		28950 => to_unsigned(11728, LUT_AMPL_WIDTH - 1),
		28951 => to_unsigned(11725, LUT_AMPL_WIDTH - 1),
		28952 => to_unsigned(11722, LUT_AMPL_WIDTH - 1),
		28953 => to_unsigned(11719, LUT_AMPL_WIDTH - 1),
		28954 => to_unsigned(11716, LUT_AMPL_WIDTH - 1),
		28955 => to_unsigned(11714, LUT_AMPL_WIDTH - 1),
		28956 => to_unsigned(11711, LUT_AMPL_WIDTH - 1),
		28957 => to_unsigned(11708, LUT_AMPL_WIDTH - 1),
		28958 => to_unsigned(11705, LUT_AMPL_WIDTH - 1),
		28959 => to_unsigned(11702, LUT_AMPL_WIDTH - 1),
		28960 => to_unsigned(11699, LUT_AMPL_WIDTH - 1),
		28961 => to_unsigned(11696, LUT_AMPL_WIDTH - 1),
		28962 => to_unsigned(11693, LUT_AMPL_WIDTH - 1),
		28963 => to_unsigned(11690, LUT_AMPL_WIDTH - 1),
		28964 => to_unsigned(11687, LUT_AMPL_WIDTH - 1),
		28965 => to_unsigned(11684, LUT_AMPL_WIDTH - 1),
		28966 => to_unsigned(11681, LUT_AMPL_WIDTH - 1),
		28967 => to_unsigned(11678, LUT_AMPL_WIDTH - 1),
		28968 => to_unsigned(11675, LUT_AMPL_WIDTH - 1),
		28969 => to_unsigned(11672, LUT_AMPL_WIDTH - 1),
		28970 => to_unsigned(11669, LUT_AMPL_WIDTH - 1),
		28971 => to_unsigned(11667, LUT_AMPL_WIDTH - 1),
		28972 => to_unsigned(11664, LUT_AMPL_WIDTH - 1),
		28973 => to_unsigned(11661, LUT_AMPL_WIDTH - 1),
		28974 => to_unsigned(11658, LUT_AMPL_WIDTH - 1),
		28975 => to_unsigned(11655, LUT_AMPL_WIDTH - 1),
		28976 => to_unsigned(11652, LUT_AMPL_WIDTH - 1),
		28977 => to_unsigned(11649, LUT_AMPL_WIDTH - 1),
		28978 => to_unsigned(11646, LUT_AMPL_WIDTH - 1),
		28979 => to_unsigned(11643, LUT_AMPL_WIDTH - 1),
		28980 => to_unsigned(11640, LUT_AMPL_WIDTH - 1),
		28981 => to_unsigned(11637, LUT_AMPL_WIDTH - 1),
		28982 => to_unsigned(11634, LUT_AMPL_WIDTH - 1),
		28983 => to_unsigned(11631, LUT_AMPL_WIDTH - 1),
		28984 => to_unsigned(11628, LUT_AMPL_WIDTH - 1),
		28985 => to_unsigned(11625, LUT_AMPL_WIDTH - 1),
		28986 => to_unsigned(11623, LUT_AMPL_WIDTH - 1),
		28987 => to_unsigned(11620, LUT_AMPL_WIDTH - 1),
		28988 => to_unsigned(11617, LUT_AMPL_WIDTH - 1),
		28989 => to_unsigned(11614, LUT_AMPL_WIDTH - 1),
		28990 => to_unsigned(11611, LUT_AMPL_WIDTH - 1),
		28991 => to_unsigned(11608, LUT_AMPL_WIDTH - 1),
		28992 => to_unsigned(11605, LUT_AMPL_WIDTH - 1),
		28993 => to_unsigned(11602, LUT_AMPL_WIDTH - 1),
		28994 => to_unsigned(11599, LUT_AMPL_WIDTH - 1),
		28995 => to_unsigned(11596, LUT_AMPL_WIDTH - 1),
		28996 => to_unsigned(11593, LUT_AMPL_WIDTH - 1),
		28997 => to_unsigned(11590, LUT_AMPL_WIDTH - 1),
		28998 => to_unsigned(11587, LUT_AMPL_WIDTH - 1),
		28999 => to_unsigned(11584, LUT_AMPL_WIDTH - 1),
		29000 => to_unsigned(11581, LUT_AMPL_WIDTH - 1),
		29001 => to_unsigned(11578, LUT_AMPL_WIDTH - 1),
		29002 => to_unsigned(11575, LUT_AMPL_WIDTH - 1),
		29003 => to_unsigned(11573, LUT_AMPL_WIDTH - 1),
		29004 => to_unsigned(11570, LUT_AMPL_WIDTH - 1),
		29005 => to_unsigned(11567, LUT_AMPL_WIDTH - 1),
		29006 => to_unsigned(11564, LUT_AMPL_WIDTH - 1),
		29007 => to_unsigned(11561, LUT_AMPL_WIDTH - 1),
		29008 => to_unsigned(11558, LUT_AMPL_WIDTH - 1),
		29009 => to_unsigned(11555, LUT_AMPL_WIDTH - 1),
		29010 => to_unsigned(11552, LUT_AMPL_WIDTH - 1),
		29011 => to_unsigned(11549, LUT_AMPL_WIDTH - 1),
		29012 => to_unsigned(11546, LUT_AMPL_WIDTH - 1),
		29013 => to_unsigned(11543, LUT_AMPL_WIDTH - 1),
		29014 => to_unsigned(11540, LUT_AMPL_WIDTH - 1),
		29015 => to_unsigned(11537, LUT_AMPL_WIDTH - 1),
		29016 => to_unsigned(11534, LUT_AMPL_WIDTH - 1),
		29017 => to_unsigned(11531, LUT_AMPL_WIDTH - 1),
		29018 => to_unsigned(11528, LUT_AMPL_WIDTH - 1),
		29019 => to_unsigned(11526, LUT_AMPL_WIDTH - 1),
		29020 => to_unsigned(11523, LUT_AMPL_WIDTH - 1),
		29021 => to_unsigned(11520, LUT_AMPL_WIDTH - 1),
		29022 => to_unsigned(11517, LUT_AMPL_WIDTH - 1),
		29023 => to_unsigned(11514, LUT_AMPL_WIDTH - 1),
		29024 => to_unsigned(11511, LUT_AMPL_WIDTH - 1),
		29025 => to_unsigned(11508, LUT_AMPL_WIDTH - 1),
		29026 => to_unsigned(11505, LUT_AMPL_WIDTH - 1),
		29027 => to_unsigned(11502, LUT_AMPL_WIDTH - 1),
		29028 => to_unsigned(11499, LUT_AMPL_WIDTH - 1),
		29029 => to_unsigned(11496, LUT_AMPL_WIDTH - 1),
		29030 => to_unsigned(11493, LUT_AMPL_WIDTH - 1),
		29031 => to_unsigned(11490, LUT_AMPL_WIDTH - 1),
		29032 => to_unsigned(11487, LUT_AMPL_WIDTH - 1),
		29033 => to_unsigned(11484, LUT_AMPL_WIDTH - 1),
		29034 => to_unsigned(11481, LUT_AMPL_WIDTH - 1),
		29035 => to_unsigned(11478, LUT_AMPL_WIDTH - 1),
		29036 => to_unsigned(11476, LUT_AMPL_WIDTH - 1),
		29037 => to_unsigned(11473, LUT_AMPL_WIDTH - 1),
		29038 => to_unsigned(11470, LUT_AMPL_WIDTH - 1),
		29039 => to_unsigned(11467, LUT_AMPL_WIDTH - 1),
		29040 => to_unsigned(11464, LUT_AMPL_WIDTH - 1),
		29041 => to_unsigned(11461, LUT_AMPL_WIDTH - 1),
		29042 => to_unsigned(11458, LUT_AMPL_WIDTH - 1),
		29043 => to_unsigned(11455, LUT_AMPL_WIDTH - 1),
		29044 => to_unsigned(11452, LUT_AMPL_WIDTH - 1),
		29045 => to_unsigned(11449, LUT_AMPL_WIDTH - 1),
		29046 => to_unsigned(11446, LUT_AMPL_WIDTH - 1),
		29047 => to_unsigned(11443, LUT_AMPL_WIDTH - 1),
		29048 => to_unsigned(11440, LUT_AMPL_WIDTH - 1),
		29049 => to_unsigned(11437, LUT_AMPL_WIDTH - 1),
		29050 => to_unsigned(11434, LUT_AMPL_WIDTH - 1),
		29051 => to_unsigned(11431, LUT_AMPL_WIDTH - 1),
		29052 => to_unsigned(11428, LUT_AMPL_WIDTH - 1),
		29053 => to_unsigned(11425, LUT_AMPL_WIDTH - 1),
		29054 => to_unsigned(11423, LUT_AMPL_WIDTH - 1),
		29055 => to_unsigned(11420, LUT_AMPL_WIDTH - 1),
		29056 => to_unsigned(11417, LUT_AMPL_WIDTH - 1),
		29057 => to_unsigned(11414, LUT_AMPL_WIDTH - 1),
		29058 => to_unsigned(11411, LUT_AMPL_WIDTH - 1),
		29059 => to_unsigned(11408, LUT_AMPL_WIDTH - 1),
		29060 => to_unsigned(11405, LUT_AMPL_WIDTH - 1),
		29061 => to_unsigned(11402, LUT_AMPL_WIDTH - 1),
		29062 => to_unsigned(11399, LUT_AMPL_WIDTH - 1),
		29063 => to_unsigned(11396, LUT_AMPL_WIDTH - 1),
		29064 => to_unsigned(11393, LUT_AMPL_WIDTH - 1),
		29065 => to_unsigned(11390, LUT_AMPL_WIDTH - 1),
		29066 => to_unsigned(11387, LUT_AMPL_WIDTH - 1),
		29067 => to_unsigned(11384, LUT_AMPL_WIDTH - 1),
		29068 => to_unsigned(11381, LUT_AMPL_WIDTH - 1),
		29069 => to_unsigned(11378, LUT_AMPL_WIDTH - 1),
		29070 => to_unsigned(11375, LUT_AMPL_WIDTH - 1),
		29071 => to_unsigned(11372, LUT_AMPL_WIDTH - 1),
		29072 => to_unsigned(11370, LUT_AMPL_WIDTH - 1),
		29073 => to_unsigned(11367, LUT_AMPL_WIDTH - 1),
		29074 => to_unsigned(11364, LUT_AMPL_WIDTH - 1),
		29075 => to_unsigned(11361, LUT_AMPL_WIDTH - 1),
		29076 => to_unsigned(11358, LUT_AMPL_WIDTH - 1),
		29077 => to_unsigned(11355, LUT_AMPL_WIDTH - 1),
		29078 => to_unsigned(11352, LUT_AMPL_WIDTH - 1),
		29079 => to_unsigned(11349, LUT_AMPL_WIDTH - 1),
		29080 => to_unsigned(11346, LUT_AMPL_WIDTH - 1),
		29081 => to_unsigned(11343, LUT_AMPL_WIDTH - 1),
		29082 => to_unsigned(11340, LUT_AMPL_WIDTH - 1),
		29083 => to_unsigned(11337, LUT_AMPL_WIDTH - 1),
		29084 => to_unsigned(11334, LUT_AMPL_WIDTH - 1),
		29085 => to_unsigned(11331, LUT_AMPL_WIDTH - 1),
		29086 => to_unsigned(11328, LUT_AMPL_WIDTH - 1),
		29087 => to_unsigned(11325, LUT_AMPL_WIDTH - 1),
		29088 => to_unsigned(11322, LUT_AMPL_WIDTH - 1),
		29089 => to_unsigned(11319, LUT_AMPL_WIDTH - 1),
		29090 => to_unsigned(11316, LUT_AMPL_WIDTH - 1),
		29091 => to_unsigned(11314, LUT_AMPL_WIDTH - 1),
		29092 => to_unsigned(11311, LUT_AMPL_WIDTH - 1),
		29093 => to_unsigned(11308, LUT_AMPL_WIDTH - 1),
		29094 => to_unsigned(11305, LUT_AMPL_WIDTH - 1),
		29095 => to_unsigned(11302, LUT_AMPL_WIDTH - 1),
		29096 => to_unsigned(11299, LUT_AMPL_WIDTH - 1),
		29097 => to_unsigned(11296, LUT_AMPL_WIDTH - 1),
		29098 => to_unsigned(11293, LUT_AMPL_WIDTH - 1),
		29099 => to_unsigned(11290, LUT_AMPL_WIDTH - 1),
		29100 => to_unsigned(11287, LUT_AMPL_WIDTH - 1),
		29101 => to_unsigned(11284, LUT_AMPL_WIDTH - 1),
		29102 => to_unsigned(11281, LUT_AMPL_WIDTH - 1),
		29103 => to_unsigned(11278, LUT_AMPL_WIDTH - 1),
		29104 => to_unsigned(11275, LUT_AMPL_WIDTH - 1),
		29105 => to_unsigned(11272, LUT_AMPL_WIDTH - 1),
		29106 => to_unsigned(11269, LUT_AMPL_WIDTH - 1),
		29107 => to_unsigned(11266, LUT_AMPL_WIDTH - 1),
		29108 => to_unsigned(11263, LUT_AMPL_WIDTH - 1),
		29109 => to_unsigned(11260, LUT_AMPL_WIDTH - 1),
		29110 => to_unsigned(11257, LUT_AMPL_WIDTH - 1),
		29111 => to_unsigned(11255, LUT_AMPL_WIDTH - 1),
		29112 => to_unsigned(11252, LUT_AMPL_WIDTH - 1),
		29113 => to_unsigned(11249, LUT_AMPL_WIDTH - 1),
		29114 => to_unsigned(11246, LUT_AMPL_WIDTH - 1),
		29115 => to_unsigned(11243, LUT_AMPL_WIDTH - 1),
		29116 => to_unsigned(11240, LUT_AMPL_WIDTH - 1),
		29117 => to_unsigned(11237, LUT_AMPL_WIDTH - 1),
		29118 => to_unsigned(11234, LUT_AMPL_WIDTH - 1),
		29119 => to_unsigned(11231, LUT_AMPL_WIDTH - 1),
		29120 => to_unsigned(11228, LUT_AMPL_WIDTH - 1),
		29121 => to_unsigned(11225, LUT_AMPL_WIDTH - 1),
		29122 => to_unsigned(11222, LUT_AMPL_WIDTH - 1),
		29123 => to_unsigned(11219, LUT_AMPL_WIDTH - 1),
		29124 => to_unsigned(11216, LUT_AMPL_WIDTH - 1),
		29125 => to_unsigned(11213, LUT_AMPL_WIDTH - 1),
		29126 => to_unsigned(11210, LUT_AMPL_WIDTH - 1),
		29127 => to_unsigned(11207, LUT_AMPL_WIDTH - 1),
		29128 => to_unsigned(11204, LUT_AMPL_WIDTH - 1),
		29129 => to_unsigned(11201, LUT_AMPL_WIDTH - 1),
		29130 => to_unsigned(11198, LUT_AMPL_WIDTH - 1),
		29131 => to_unsigned(11195, LUT_AMPL_WIDTH - 1),
		29132 => to_unsigned(11193, LUT_AMPL_WIDTH - 1),
		29133 => to_unsigned(11190, LUT_AMPL_WIDTH - 1),
		29134 => to_unsigned(11187, LUT_AMPL_WIDTH - 1),
		29135 => to_unsigned(11184, LUT_AMPL_WIDTH - 1),
		29136 => to_unsigned(11181, LUT_AMPL_WIDTH - 1),
		29137 => to_unsigned(11178, LUT_AMPL_WIDTH - 1),
		29138 => to_unsigned(11175, LUT_AMPL_WIDTH - 1),
		29139 => to_unsigned(11172, LUT_AMPL_WIDTH - 1),
		29140 => to_unsigned(11169, LUT_AMPL_WIDTH - 1),
		29141 => to_unsigned(11166, LUT_AMPL_WIDTH - 1),
		29142 => to_unsigned(11163, LUT_AMPL_WIDTH - 1),
		29143 => to_unsigned(11160, LUT_AMPL_WIDTH - 1),
		29144 => to_unsigned(11157, LUT_AMPL_WIDTH - 1),
		29145 => to_unsigned(11154, LUT_AMPL_WIDTH - 1),
		29146 => to_unsigned(11151, LUT_AMPL_WIDTH - 1),
		29147 => to_unsigned(11148, LUT_AMPL_WIDTH - 1),
		29148 => to_unsigned(11145, LUT_AMPL_WIDTH - 1),
		29149 => to_unsigned(11142, LUT_AMPL_WIDTH - 1),
		29150 => to_unsigned(11139, LUT_AMPL_WIDTH - 1),
		29151 => to_unsigned(11136, LUT_AMPL_WIDTH - 1),
		29152 => to_unsigned(11133, LUT_AMPL_WIDTH - 1),
		29153 => to_unsigned(11131, LUT_AMPL_WIDTH - 1),
		29154 => to_unsigned(11128, LUT_AMPL_WIDTH - 1),
		29155 => to_unsigned(11125, LUT_AMPL_WIDTH - 1),
		29156 => to_unsigned(11122, LUT_AMPL_WIDTH - 1),
		29157 => to_unsigned(11119, LUT_AMPL_WIDTH - 1),
		29158 => to_unsigned(11116, LUT_AMPL_WIDTH - 1),
		29159 => to_unsigned(11113, LUT_AMPL_WIDTH - 1),
		29160 => to_unsigned(11110, LUT_AMPL_WIDTH - 1),
		29161 => to_unsigned(11107, LUT_AMPL_WIDTH - 1),
		29162 => to_unsigned(11104, LUT_AMPL_WIDTH - 1),
		29163 => to_unsigned(11101, LUT_AMPL_WIDTH - 1),
		29164 => to_unsigned(11098, LUT_AMPL_WIDTH - 1),
		29165 => to_unsigned(11095, LUT_AMPL_WIDTH - 1),
		29166 => to_unsigned(11092, LUT_AMPL_WIDTH - 1),
		29167 => to_unsigned(11089, LUT_AMPL_WIDTH - 1),
		29168 => to_unsigned(11086, LUT_AMPL_WIDTH - 1),
		29169 => to_unsigned(11083, LUT_AMPL_WIDTH - 1),
		29170 => to_unsigned(11080, LUT_AMPL_WIDTH - 1),
		29171 => to_unsigned(11077, LUT_AMPL_WIDTH - 1),
		29172 => to_unsigned(11074, LUT_AMPL_WIDTH - 1),
		29173 => to_unsigned(11071, LUT_AMPL_WIDTH - 1),
		29174 => to_unsigned(11068, LUT_AMPL_WIDTH - 1),
		29175 => to_unsigned(11065, LUT_AMPL_WIDTH - 1),
		29176 => to_unsigned(11063, LUT_AMPL_WIDTH - 1),
		29177 => to_unsigned(11060, LUT_AMPL_WIDTH - 1),
		29178 => to_unsigned(11057, LUT_AMPL_WIDTH - 1),
		29179 => to_unsigned(11054, LUT_AMPL_WIDTH - 1),
		29180 => to_unsigned(11051, LUT_AMPL_WIDTH - 1),
		29181 => to_unsigned(11048, LUT_AMPL_WIDTH - 1),
		29182 => to_unsigned(11045, LUT_AMPL_WIDTH - 1),
		29183 => to_unsigned(11042, LUT_AMPL_WIDTH - 1),
		29184 => to_unsigned(11039, LUT_AMPL_WIDTH - 1),
		29185 => to_unsigned(11036, LUT_AMPL_WIDTH - 1),
		29186 => to_unsigned(11033, LUT_AMPL_WIDTH - 1),
		29187 => to_unsigned(11030, LUT_AMPL_WIDTH - 1),
		29188 => to_unsigned(11027, LUT_AMPL_WIDTH - 1),
		29189 => to_unsigned(11024, LUT_AMPL_WIDTH - 1),
		29190 => to_unsigned(11021, LUT_AMPL_WIDTH - 1),
		29191 => to_unsigned(11018, LUT_AMPL_WIDTH - 1),
		29192 => to_unsigned(11015, LUT_AMPL_WIDTH - 1),
		29193 => to_unsigned(11012, LUT_AMPL_WIDTH - 1),
		29194 => to_unsigned(11009, LUT_AMPL_WIDTH - 1),
		29195 => to_unsigned(11006, LUT_AMPL_WIDTH - 1),
		29196 => to_unsigned(11003, LUT_AMPL_WIDTH - 1),
		29197 => to_unsigned(11000, LUT_AMPL_WIDTH - 1),
		29198 => to_unsigned(10997, LUT_AMPL_WIDTH - 1),
		29199 => to_unsigned(10994, LUT_AMPL_WIDTH - 1),
		29200 => to_unsigned(10992, LUT_AMPL_WIDTH - 1),
		29201 => to_unsigned(10989, LUT_AMPL_WIDTH - 1),
		29202 => to_unsigned(10986, LUT_AMPL_WIDTH - 1),
		29203 => to_unsigned(10983, LUT_AMPL_WIDTH - 1),
		29204 => to_unsigned(10980, LUT_AMPL_WIDTH - 1),
		29205 => to_unsigned(10977, LUT_AMPL_WIDTH - 1),
		29206 => to_unsigned(10974, LUT_AMPL_WIDTH - 1),
		29207 => to_unsigned(10971, LUT_AMPL_WIDTH - 1),
		29208 => to_unsigned(10968, LUT_AMPL_WIDTH - 1),
		29209 => to_unsigned(10965, LUT_AMPL_WIDTH - 1),
		29210 => to_unsigned(10962, LUT_AMPL_WIDTH - 1),
		29211 => to_unsigned(10959, LUT_AMPL_WIDTH - 1),
		29212 => to_unsigned(10956, LUT_AMPL_WIDTH - 1),
		29213 => to_unsigned(10953, LUT_AMPL_WIDTH - 1),
		29214 => to_unsigned(10950, LUT_AMPL_WIDTH - 1),
		29215 => to_unsigned(10947, LUT_AMPL_WIDTH - 1),
		29216 => to_unsigned(10944, LUT_AMPL_WIDTH - 1),
		29217 => to_unsigned(10941, LUT_AMPL_WIDTH - 1),
		29218 => to_unsigned(10938, LUT_AMPL_WIDTH - 1),
		29219 => to_unsigned(10935, LUT_AMPL_WIDTH - 1),
		29220 => to_unsigned(10932, LUT_AMPL_WIDTH - 1),
		29221 => to_unsigned(10929, LUT_AMPL_WIDTH - 1),
		29222 => to_unsigned(10926, LUT_AMPL_WIDTH - 1),
		29223 => to_unsigned(10923, LUT_AMPL_WIDTH - 1),
		29224 => to_unsigned(10920, LUT_AMPL_WIDTH - 1),
		29225 => to_unsigned(10918, LUT_AMPL_WIDTH - 1),
		29226 => to_unsigned(10915, LUT_AMPL_WIDTH - 1),
		29227 => to_unsigned(10912, LUT_AMPL_WIDTH - 1),
		29228 => to_unsigned(10909, LUT_AMPL_WIDTH - 1),
		29229 => to_unsigned(10906, LUT_AMPL_WIDTH - 1),
		29230 => to_unsigned(10903, LUT_AMPL_WIDTH - 1),
		29231 => to_unsigned(10900, LUT_AMPL_WIDTH - 1),
		29232 => to_unsigned(10897, LUT_AMPL_WIDTH - 1),
		29233 => to_unsigned(10894, LUT_AMPL_WIDTH - 1),
		29234 => to_unsigned(10891, LUT_AMPL_WIDTH - 1),
		29235 => to_unsigned(10888, LUT_AMPL_WIDTH - 1),
		29236 => to_unsigned(10885, LUT_AMPL_WIDTH - 1),
		29237 => to_unsigned(10882, LUT_AMPL_WIDTH - 1),
		29238 => to_unsigned(10879, LUT_AMPL_WIDTH - 1),
		29239 => to_unsigned(10876, LUT_AMPL_WIDTH - 1),
		29240 => to_unsigned(10873, LUT_AMPL_WIDTH - 1),
		29241 => to_unsigned(10870, LUT_AMPL_WIDTH - 1),
		29242 => to_unsigned(10867, LUT_AMPL_WIDTH - 1),
		29243 => to_unsigned(10864, LUT_AMPL_WIDTH - 1),
		29244 => to_unsigned(10861, LUT_AMPL_WIDTH - 1),
		29245 => to_unsigned(10858, LUT_AMPL_WIDTH - 1),
		29246 => to_unsigned(10855, LUT_AMPL_WIDTH - 1),
		29247 => to_unsigned(10852, LUT_AMPL_WIDTH - 1),
		29248 => to_unsigned(10849, LUT_AMPL_WIDTH - 1),
		29249 => to_unsigned(10846, LUT_AMPL_WIDTH - 1),
		29250 => to_unsigned(10843, LUT_AMPL_WIDTH - 1),
		29251 => to_unsigned(10840, LUT_AMPL_WIDTH - 1),
		29252 => to_unsigned(10838, LUT_AMPL_WIDTH - 1),
		29253 => to_unsigned(10835, LUT_AMPL_WIDTH - 1),
		29254 => to_unsigned(10832, LUT_AMPL_WIDTH - 1),
		29255 => to_unsigned(10829, LUT_AMPL_WIDTH - 1),
		29256 => to_unsigned(10826, LUT_AMPL_WIDTH - 1),
		29257 => to_unsigned(10823, LUT_AMPL_WIDTH - 1),
		29258 => to_unsigned(10820, LUT_AMPL_WIDTH - 1),
		29259 => to_unsigned(10817, LUT_AMPL_WIDTH - 1),
		29260 => to_unsigned(10814, LUT_AMPL_WIDTH - 1),
		29261 => to_unsigned(10811, LUT_AMPL_WIDTH - 1),
		29262 => to_unsigned(10808, LUT_AMPL_WIDTH - 1),
		29263 => to_unsigned(10805, LUT_AMPL_WIDTH - 1),
		29264 => to_unsigned(10802, LUT_AMPL_WIDTH - 1),
		29265 => to_unsigned(10799, LUT_AMPL_WIDTH - 1),
		29266 => to_unsigned(10796, LUT_AMPL_WIDTH - 1),
		29267 => to_unsigned(10793, LUT_AMPL_WIDTH - 1),
		29268 => to_unsigned(10790, LUT_AMPL_WIDTH - 1),
		29269 => to_unsigned(10787, LUT_AMPL_WIDTH - 1),
		29270 => to_unsigned(10784, LUT_AMPL_WIDTH - 1),
		29271 => to_unsigned(10781, LUT_AMPL_WIDTH - 1),
		29272 => to_unsigned(10778, LUT_AMPL_WIDTH - 1),
		29273 => to_unsigned(10775, LUT_AMPL_WIDTH - 1),
		29274 => to_unsigned(10772, LUT_AMPL_WIDTH - 1),
		29275 => to_unsigned(10769, LUT_AMPL_WIDTH - 1),
		29276 => to_unsigned(10766, LUT_AMPL_WIDTH - 1),
		29277 => to_unsigned(10763, LUT_AMPL_WIDTH - 1),
		29278 => to_unsigned(10760, LUT_AMPL_WIDTH - 1),
		29279 => to_unsigned(10757, LUT_AMPL_WIDTH - 1),
		29280 => to_unsigned(10754, LUT_AMPL_WIDTH - 1),
		29281 => to_unsigned(10751, LUT_AMPL_WIDTH - 1),
		29282 => to_unsigned(10749, LUT_AMPL_WIDTH - 1),
		29283 => to_unsigned(10746, LUT_AMPL_WIDTH - 1),
		29284 => to_unsigned(10743, LUT_AMPL_WIDTH - 1),
		29285 => to_unsigned(10740, LUT_AMPL_WIDTH - 1),
		29286 => to_unsigned(10737, LUT_AMPL_WIDTH - 1),
		29287 => to_unsigned(10734, LUT_AMPL_WIDTH - 1),
		29288 => to_unsigned(10731, LUT_AMPL_WIDTH - 1),
		29289 => to_unsigned(10728, LUT_AMPL_WIDTH - 1),
		29290 => to_unsigned(10725, LUT_AMPL_WIDTH - 1),
		29291 => to_unsigned(10722, LUT_AMPL_WIDTH - 1),
		29292 => to_unsigned(10719, LUT_AMPL_WIDTH - 1),
		29293 => to_unsigned(10716, LUT_AMPL_WIDTH - 1),
		29294 => to_unsigned(10713, LUT_AMPL_WIDTH - 1),
		29295 => to_unsigned(10710, LUT_AMPL_WIDTH - 1),
		29296 => to_unsigned(10707, LUT_AMPL_WIDTH - 1),
		29297 => to_unsigned(10704, LUT_AMPL_WIDTH - 1),
		29298 => to_unsigned(10701, LUT_AMPL_WIDTH - 1),
		29299 => to_unsigned(10698, LUT_AMPL_WIDTH - 1),
		29300 => to_unsigned(10695, LUT_AMPL_WIDTH - 1),
		29301 => to_unsigned(10692, LUT_AMPL_WIDTH - 1),
		29302 => to_unsigned(10689, LUT_AMPL_WIDTH - 1),
		29303 => to_unsigned(10686, LUT_AMPL_WIDTH - 1),
		29304 => to_unsigned(10683, LUT_AMPL_WIDTH - 1),
		29305 => to_unsigned(10680, LUT_AMPL_WIDTH - 1),
		29306 => to_unsigned(10677, LUT_AMPL_WIDTH - 1),
		29307 => to_unsigned(10674, LUT_AMPL_WIDTH - 1),
		29308 => to_unsigned(10671, LUT_AMPL_WIDTH - 1),
		29309 => to_unsigned(10668, LUT_AMPL_WIDTH - 1),
		29310 => to_unsigned(10665, LUT_AMPL_WIDTH - 1),
		29311 => to_unsigned(10662, LUT_AMPL_WIDTH - 1),
		29312 => to_unsigned(10659, LUT_AMPL_WIDTH - 1),
		29313 => to_unsigned(10656, LUT_AMPL_WIDTH - 1),
		29314 => to_unsigned(10654, LUT_AMPL_WIDTH - 1),
		29315 => to_unsigned(10651, LUT_AMPL_WIDTH - 1),
		29316 => to_unsigned(10648, LUT_AMPL_WIDTH - 1),
		29317 => to_unsigned(10645, LUT_AMPL_WIDTH - 1),
		29318 => to_unsigned(10642, LUT_AMPL_WIDTH - 1),
		29319 => to_unsigned(10639, LUT_AMPL_WIDTH - 1),
		29320 => to_unsigned(10636, LUT_AMPL_WIDTH - 1),
		29321 => to_unsigned(10633, LUT_AMPL_WIDTH - 1),
		29322 => to_unsigned(10630, LUT_AMPL_WIDTH - 1),
		29323 => to_unsigned(10627, LUT_AMPL_WIDTH - 1),
		29324 => to_unsigned(10624, LUT_AMPL_WIDTH - 1),
		29325 => to_unsigned(10621, LUT_AMPL_WIDTH - 1),
		29326 => to_unsigned(10618, LUT_AMPL_WIDTH - 1),
		29327 => to_unsigned(10615, LUT_AMPL_WIDTH - 1),
		29328 => to_unsigned(10612, LUT_AMPL_WIDTH - 1),
		29329 => to_unsigned(10609, LUT_AMPL_WIDTH - 1),
		29330 => to_unsigned(10606, LUT_AMPL_WIDTH - 1),
		29331 => to_unsigned(10603, LUT_AMPL_WIDTH - 1),
		29332 => to_unsigned(10600, LUT_AMPL_WIDTH - 1),
		29333 => to_unsigned(10597, LUT_AMPL_WIDTH - 1),
		29334 => to_unsigned(10594, LUT_AMPL_WIDTH - 1),
		29335 => to_unsigned(10591, LUT_AMPL_WIDTH - 1),
		29336 => to_unsigned(10588, LUT_AMPL_WIDTH - 1),
		29337 => to_unsigned(10585, LUT_AMPL_WIDTH - 1),
		29338 => to_unsigned(10582, LUT_AMPL_WIDTH - 1),
		29339 => to_unsigned(10579, LUT_AMPL_WIDTH - 1),
		29340 => to_unsigned(10576, LUT_AMPL_WIDTH - 1),
		29341 => to_unsigned(10573, LUT_AMPL_WIDTH - 1),
		29342 => to_unsigned(10570, LUT_AMPL_WIDTH - 1),
		29343 => to_unsigned(10567, LUT_AMPL_WIDTH - 1),
		29344 => to_unsigned(10564, LUT_AMPL_WIDTH - 1),
		29345 => to_unsigned(10561, LUT_AMPL_WIDTH - 1),
		29346 => to_unsigned(10558, LUT_AMPL_WIDTH - 1),
		29347 => to_unsigned(10555, LUT_AMPL_WIDTH - 1),
		29348 => to_unsigned(10552, LUT_AMPL_WIDTH - 1),
		29349 => to_unsigned(10549, LUT_AMPL_WIDTH - 1),
		29350 => to_unsigned(10546, LUT_AMPL_WIDTH - 1),
		29351 => to_unsigned(10544, LUT_AMPL_WIDTH - 1),
		29352 => to_unsigned(10541, LUT_AMPL_WIDTH - 1),
		29353 => to_unsigned(10538, LUT_AMPL_WIDTH - 1),
		29354 => to_unsigned(10535, LUT_AMPL_WIDTH - 1),
		29355 => to_unsigned(10532, LUT_AMPL_WIDTH - 1),
		29356 => to_unsigned(10529, LUT_AMPL_WIDTH - 1),
		29357 => to_unsigned(10526, LUT_AMPL_WIDTH - 1),
		29358 => to_unsigned(10523, LUT_AMPL_WIDTH - 1),
		29359 => to_unsigned(10520, LUT_AMPL_WIDTH - 1),
		29360 => to_unsigned(10517, LUT_AMPL_WIDTH - 1),
		29361 => to_unsigned(10514, LUT_AMPL_WIDTH - 1),
		29362 => to_unsigned(10511, LUT_AMPL_WIDTH - 1),
		29363 => to_unsigned(10508, LUT_AMPL_WIDTH - 1),
		29364 => to_unsigned(10505, LUT_AMPL_WIDTH - 1),
		29365 => to_unsigned(10502, LUT_AMPL_WIDTH - 1),
		29366 => to_unsigned(10499, LUT_AMPL_WIDTH - 1),
		29367 => to_unsigned(10496, LUT_AMPL_WIDTH - 1),
		29368 => to_unsigned(10493, LUT_AMPL_WIDTH - 1),
		29369 => to_unsigned(10490, LUT_AMPL_WIDTH - 1),
		29370 => to_unsigned(10487, LUT_AMPL_WIDTH - 1),
		29371 => to_unsigned(10484, LUT_AMPL_WIDTH - 1),
		29372 => to_unsigned(10481, LUT_AMPL_WIDTH - 1),
		29373 => to_unsigned(10478, LUT_AMPL_WIDTH - 1),
		29374 => to_unsigned(10475, LUT_AMPL_WIDTH - 1),
		29375 => to_unsigned(10472, LUT_AMPL_WIDTH - 1),
		29376 => to_unsigned(10469, LUT_AMPL_WIDTH - 1),
		29377 => to_unsigned(10466, LUT_AMPL_WIDTH - 1),
		29378 => to_unsigned(10463, LUT_AMPL_WIDTH - 1),
		29379 => to_unsigned(10460, LUT_AMPL_WIDTH - 1),
		29380 => to_unsigned(10457, LUT_AMPL_WIDTH - 1),
		29381 => to_unsigned(10454, LUT_AMPL_WIDTH - 1),
		29382 => to_unsigned(10451, LUT_AMPL_WIDTH - 1),
		29383 => to_unsigned(10448, LUT_AMPL_WIDTH - 1),
		29384 => to_unsigned(10445, LUT_AMPL_WIDTH - 1),
		29385 => to_unsigned(10442, LUT_AMPL_WIDTH - 1),
		29386 => to_unsigned(10439, LUT_AMPL_WIDTH - 1),
		29387 => to_unsigned(10436, LUT_AMPL_WIDTH - 1),
		29388 => to_unsigned(10433, LUT_AMPL_WIDTH - 1),
		29389 => to_unsigned(10430, LUT_AMPL_WIDTH - 1),
		29390 => to_unsigned(10427, LUT_AMPL_WIDTH - 1),
		29391 => to_unsigned(10424, LUT_AMPL_WIDTH - 1),
		29392 => to_unsigned(10421, LUT_AMPL_WIDTH - 1),
		29393 => to_unsigned(10419, LUT_AMPL_WIDTH - 1),
		29394 => to_unsigned(10416, LUT_AMPL_WIDTH - 1),
		29395 => to_unsigned(10413, LUT_AMPL_WIDTH - 1),
		29396 => to_unsigned(10410, LUT_AMPL_WIDTH - 1),
		29397 => to_unsigned(10407, LUT_AMPL_WIDTH - 1),
		29398 => to_unsigned(10404, LUT_AMPL_WIDTH - 1),
		29399 => to_unsigned(10401, LUT_AMPL_WIDTH - 1),
		29400 => to_unsigned(10398, LUT_AMPL_WIDTH - 1),
		29401 => to_unsigned(10395, LUT_AMPL_WIDTH - 1),
		29402 => to_unsigned(10392, LUT_AMPL_WIDTH - 1),
		29403 => to_unsigned(10389, LUT_AMPL_WIDTH - 1),
		29404 => to_unsigned(10386, LUT_AMPL_WIDTH - 1),
		29405 => to_unsigned(10383, LUT_AMPL_WIDTH - 1),
		29406 => to_unsigned(10380, LUT_AMPL_WIDTH - 1),
		29407 => to_unsigned(10377, LUT_AMPL_WIDTH - 1),
		29408 => to_unsigned(10374, LUT_AMPL_WIDTH - 1),
		29409 => to_unsigned(10371, LUT_AMPL_WIDTH - 1),
		29410 => to_unsigned(10368, LUT_AMPL_WIDTH - 1),
		29411 => to_unsigned(10365, LUT_AMPL_WIDTH - 1),
		29412 => to_unsigned(10362, LUT_AMPL_WIDTH - 1),
		29413 => to_unsigned(10359, LUT_AMPL_WIDTH - 1),
		29414 => to_unsigned(10356, LUT_AMPL_WIDTH - 1),
		29415 => to_unsigned(10353, LUT_AMPL_WIDTH - 1),
		29416 => to_unsigned(10350, LUT_AMPL_WIDTH - 1),
		29417 => to_unsigned(10347, LUT_AMPL_WIDTH - 1),
		29418 => to_unsigned(10344, LUT_AMPL_WIDTH - 1),
		29419 => to_unsigned(10341, LUT_AMPL_WIDTH - 1),
		29420 => to_unsigned(10338, LUT_AMPL_WIDTH - 1),
		29421 => to_unsigned(10335, LUT_AMPL_WIDTH - 1),
		29422 => to_unsigned(10332, LUT_AMPL_WIDTH - 1),
		29423 => to_unsigned(10329, LUT_AMPL_WIDTH - 1),
		29424 => to_unsigned(10326, LUT_AMPL_WIDTH - 1),
		29425 => to_unsigned(10323, LUT_AMPL_WIDTH - 1),
		29426 => to_unsigned(10320, LUT_AMPL_WIDTH - 1),
		29427 => to_unsigned(10317, LUT_AMPL_WIDTH - 1),
		29428 => to_unsigned(10314, LUT_AMPL_WIDTH - 1),
		29429 => to_unsigned(10311, LUT_AMPL_WIDTH - 1),
		29430 => to_unsigned(10308, LUT_AMPL_WIDTH - 1),
		29431 => to_unsigned(10305, LUT_AMPL_WIDTH - 1),
		29432 => to_unsigned(10302, LUT_AMPL_WIDTH - 1),
		29433 => to_unsigned(10299, LUT_AMPL_WIDTH - 1),
		29434 => to_unsigned(10296, LUT_AMPL_WIDTH - 1),
		29435 => to_unsigned(10293, LUT_AMPL_WIDTH - 1),
		29436 => to_unsigned(10290, LUT_AMPL_WIDTH - 1),
		29437 => to_unsigned(10287, LUT_AMPL_WIDTH - 1),
		29438 => to_unsigned(10284, LUT_AMPL_WIDTH - 1),
		29439 => to_unsigned(10281, LUT_AMPL_WIDTH - 1),
		29440 => to_unsigned(10278, LUT_AMPL_WIDTH - 1),
		29441 => to_unsigned(10275, LUT_AMPL_WIDTH - 1),
		29442 => to_unsigned(10272, LUT_AMPL_WIDTH - 1),
		29443 => to_unsigned(10269, LUT_AMPL_WIDTH - 1),
		29444 => to_unsigned(10266, LUT_AMPL_WIDTH - 1),
		29445 => to_unsigned(10263, LUT_AMPL_WIDTH - 1),
		29446 => to_unsigned(10261, LUT_AMPL_WIDTH - 1),
		29447 => to_unsigned(10258, LUT_AMPL_WIDTH - 1),
		29448 => to_unsigned(10255, LUT_AMPL_WIDTH - 1),
		29449 => to_unsigned(10252, LUT_AMPL_WIDTH - 1),
		29450 => to_unsigned(10249, LUT_AMPL_WIDTH - 1),
		29451 => to_unsigned(10246, LUT_AMPL_WIDTH - 1),
		29452 => to_unsigned(10243, LUT_AMPL_WIDTH - 1),
		29453 => to_unsigned(10240, LUT_AMPL_WIDTH - 1),
		29454 => to_unsigned(10237, LUT_AMPL_WIDTH - 1),
		29455 => to_unsigned(10234, LUT_AMPL_WIDTH - 1),
		29456 => to_unsigned(10231, LUT_AMPL_WIDTH - 1),
		29457 => to_unsigned(10228, LUT_AMPL_WIDTH - 1),
		29458 => to_unsigned(10225, LUT_AMPL_WIDTH - 1),
		29459 => to_unsigned(10222, LUT_AMPL_WIDTH - 1),
		29460 => to_unsigned(10219, LUT_AMPL_WIDTH - 1),
		29461 => to_unsigned(10216, LUT_AMPL_WIDTH - 1),
		29462 => to_unsigned(10213, LUT_AMPL_WIDTH - 1),
		29463 => to_unsigned(10210, LUT_AMPL_WIDTH - 1),
		29464 => to_unsigned(10207, LUT_AMPL_WIDTH - 1),
		29465 => to_unsigned(10204, LUT_AMPL_WIDTH - 1),
		29466 => to_unsigned(10201, LUT_AMPL_WIDTH - 1),
		29467 => to_unsigned(10198, LUT_AMPL_WIDTH - 1),
		29468 => to_unsigned(10195, LUT_AMPL_WIDTH - 1),
		29469 => to_unsigned(10192, LUT_AMPL_WIDTH - 1),
		29470 => to_unsigned(10189, LUT_AMPL_WIDTH - 1),
		29471 => to_unsigned(10186, LUT_AMPL_WIDTH - 1),
		29472 => to_unsigned(10183, LUT_AMPL_WIDTH - 1),
		29473 => to_unsigned(10180, LUT_AMPL_WIDTH - 1),
		29474 => to_unsigned(10177, LUT_AMPL_WIDTH - 1),
		29475 => to_unsigned(10174, LUT_AMPL_WIDTH - 1),
		29476 => to_unsigned(10171, LUT_AMPL_WIDTH - 1),
		29477 => to_unsigned(10168, LUT_AMPL_WIDTH - 1),
		29478 => to_unsigned(10165, LUT_AMPL_WIDTH - 1),
		29479 => to_unsigned(10162, LUT_AMPL_WIDTH - 1),
		29480 => to_unsigned(10159, LUT_AMPL_WIDTH - 1),
		29481 => to_unsigned(10156, LUT_AMPL_WIDTH - 1),
		29482 => to_unsigned(10153, LUT_AMPL_WIDTH - 1),
		29483 => to_unsigned(10150, LUT_AMPL_WIDTH - 1),
		29484 => to_unsigned(10147, LUT_AMPL_WIDTH - 1),
		29485 => to_unsigned(10144, LUT_AMPL_WIDTH - 1),
		29486 => to_unsigned(10141, LUT_AMPL_WIDTH - 1),
		29487 => to_unsigned(10138, LUT_AMPL_WIDTH - 1),
		29488 => to_unsigned(10135, LUT_AMPL_WIDTH - 1),
		29489 => to_unsigned(10132, LUT_AMPL_WIDTH - 1),
		29490 => to_unsigned(10129, LUT_AMPL_WIDTH - 1),
		29491 => to_unsigned(10126, LUT_AMPL_WIDTH - 1),
		29492 => to_unsigned(10123, LUT_AMPL_WIDTH - 1),
		29493 => to_unsigned(10120, LUT_AMPL_WIDTH - 1),
		29494 => to_unsigned(10117, LUT_AMPL_WIDTH - 1),
		29495 => to_unsigned(10114, LUT_AMPL_WIDTH - 1),
		29496 => to_unsigned(10111, LUT_AMPL_WIDTH - 1),
		29497 => to_unsigned(10108, LUT_AMPL_WIDTH - 1),
		29498 => to_unsigned(10105, LUT_AMPL_WIDTH - 1),
		29499 => to_unsigned(10102, LUT_AMPL_WIDTH - 1),
		29500 => to_unsigned(10099, LUT_AMPL_WIDTH - 1),
		29501 => to_unsigned(10096, LUT_AMPL_WIDTH - 1),
		29502 => to_unsigned(10093, LUT_AMPL_WIDTH - 1),
		29503 => to_unsigned(10090, LUT_AMPL_WIDTH - 1),
		29504 => to_unsigned(10087, LUT_AMPL_WIDTH - 1),
		29505 => to_unsigned(10084, LUT_AMPL_WIDTH - 1),
		29506 => to_unsigned(10081, LUT_AMPL_WIDTH - 1),
		29507 => to_unsigned(10078, LUT_AMPL_WIDTH - 1),
		29508 => to_unsigned(10075, LUT_AMPL_WIDTH - 1),
		29509 => to_unsigned(10072, LUT_AMPL_WIDTH - 1),
		29510 => to_unsigned(10069, LUT_AMPL_WIDTH - 1),
		29511 => to_unsigned(10066, LUT_AMPL_WIDTH - 1),
		29512 => to_unsigned(10063, LUT_AMPL_WIDTH - 1),
		29513 => to_unsigned(10060, LUT_AMPL_WIDTH - 1),
		29514 => to_unsigned(10057, LUT_AMPL_WIDTH - 1),
		29515 => to_unsigned(10054, LUT_AMPL_WIDTH - 1),
		29516 => to_unsigned(10051, LUT_AMPL_WIDTH - 1),
		29517 => to_unsigned(10048, LUT_AMPL_WIDTH - 1),
		29518 => to_unsigned(10045, LUT_AMPL_WIDTH - 1),
		29519 => to_unsigned(10042, LUT_AMPL_WIDTH - 1),
		29520 => to_unsigned(10039, LUT_AMPL_WIDTH - 1),
		29521 => to_unsigned(10036, LUT_AMPL_WIDTH - 1),
		29522 => to_unsigned(10033, LUT_AMPL_WIDTH - 1),
		29523 => to_unsigned(10031, LUT_AMPL_WIDTH - 1),
		29524 => to_unsigned(10028, LUT_AMPL_WIDTH - 1),
		29525 => to_unsigned(10025, LUT_AMPL_WIDTH - 1),
		29526 => to_unsigned(10022, LUT_AMPL_WIDTH - 1),
		29527 => to_unsigned(10019, LUT_AMPL_WIDTH - 1),
		29528 => to_unsigned(10016, LUT_AMPL_WIDTH - 1),
		29529 => to_unsigned(10013, LUT_AMPL_WIDTH - 1),
		29530 => to_unsigned(10010, LUT_AMPL_WIDTH - 1),
		29531 => to_unsigned(10007, LUT_AMPL_WIDTH - 1),
		29532 => to_unsigned(10004, LUT_AMPL_WIDTH - 1),
		29533 => to_unsigned(10001, LUT_AMPL_WIDTH - 1),
		29534 => to_unsigned(9998, LUT_AMPL_WIDTH - 1),
		29535 => to_unsigned(9995, LUT_AMPL_WIDTH - 1),
		29536 => to_unsigned(9992, LUT_AMPL_WIDTH - 1),
		29537 => to_unsigned(9989, LUT_AMPL_WIDTH - 1),
		29538 => to_unsigned(9986, LUT_AMPL_WIDTH - 1),
		29539 => to_unsigned(9983, LUT_AMPL_WIDTH - 1),
		29540 => to_unsigned(9980, LUT_AMPL_WIDTH - 1),
		29541 => to_unsigned(9977, LUT_AMPL_WIDTH - 1),
		29542 => to_unsigned(9974, LUT_AMPL_WIDTH - 1),
		29543 => to_unsigned(9971, LUT_AMPL_WIDTH - 1),
		29544 => to_unsigned(9968, LUT_AMPL_WIDTH - 1),
		29545 => to_unsigned(9965, LUT_AMPL_WIDTH - 1),
		29546 => to_unsigned(9962, LUT_AMPL_WIDTH - 1),
		29547 => to_unsigned(9959, LUT_AMPL_WIDTH - 1),
		29548 => to_unsigned(9956, LUT_AMPL_WIDTH - 1),
		29549 => to_unsigned(9953, LUT_AMPL_WIDTH - 1),
		29550 => to_unsigned(9950, LUT_AMPL_WIDTH - 1),
		29551 => to_unsigned(9947, LUT_AMPL_WIDTH - 1),
		29552 => to_unsigned(9944, LUT_AMPL_WIDTH - 1),
		29553 => to_unsigned(9941, LUT_AMPL_WIDTH - 1),
		29554 => to_unsigned(9938, LUT_AMPL_WIDTH - 1),
		29555 => to_unsigned(9935, LUT_AMPL_WIDTH - 1),
		29556 => to_unsigned(9932, LUT_AMPL_WIDTH - 1),
		29557 => to_unsigned(9929, LUT_AMPL_WIDTH - 1),
		29558 => to_unsigned(9926, LUT_AMPL_WIDTH - 1),
		29559 => to_unsigned(9923, LUT_AMPL_WIDTH - 1),
		29560 => to_unsigned(9920, LUT_AMPL_WIDTH - 1),
		29561 => to_unsigned(9917, LUT_AMPL_WIDTH - 1),
		29562 => to_unsigned(9914, LUT_AMPL_WIDTH - 1),
		29563 => to_unsigned(9911, LUT_AMPL_WIDTH - 1),
		29564 => to_unsigned(9908, LUT_AMPL_WIDTH - 1),
		29565 => to_unsigned(9905, LUT_AMPL_WIDTH - 1),
		29566 => to_unsigned(9902, LUT_AMPL_WIDTH - 1),
		29567 => to_unsigned(9899, LUT_AMPL_WIDTH - 1),
		29568 => to_unsigned(9896, LUT_AMPL_WIDTH - 1),
		29569 => to_unsigned(9893, LUT_AMPL_WIDTH - 1),
		29570 => to_unsigned(9890, LUT_AMPL_WIDTH - 1),
		29571 => to_unsigned(9887, LUT_AMPL_WIDTH - 1),
		29572 => to_unsigned(9884, LUT_AMPL_WIDTH - 1),
		29573 => to_unsigned(9881, LUT_AMPL_WIDTH - 1),
		29574 => to_unsigned(9878, LUT_AMPL_WIDTH - 1),
		29575 => to_unsigned(9875, LUT_AMPL_WIDTH - 1),
		29576 => to_unsigned(9872, LUT_AMPL_WIDTH - 1),
		29577 => to_unsigned(9869, LUT_AMPL_WIDTH - 1),
		29578 => to_unsigned(9866, LUT_AMPL_WIDTH - 1),
		29579 => to_unsigned(9863, LUT_AMPL_WIDTH - 1),
		29580 => to_unsigned(9860, LUT_AMPL_WIDTH - 1),
		29581 => to_unsigned(9857, LUT_AMPL_WIDTH - 1),
		29582 => to_unsigned(9854, LUT_AMPL_WIDTH - 1),
		29583 => to_unsigned(9851, LUT_AMPL_WIDTH - 1),
		29584 => to_unsigned(9848, LUT_AMPL_WIDTH - 1),
		29585 => to_unsigned(9845, LUT_AMPL_WIDTH - 1),
		29586 => to_unsigned(9842, LUT_AMPL_WIDTH - 1),
		29587 => to_unsigned(9839, LUT_AMPL_WIDTH - 1),
		29588 => to_unsigned(9836, LUT_AMPL_WIDTH - 1),
		29589 => to_unsigned(9833, LUT_AMPL_WIDTH - 1),
		29590 => to_unsigned(9830, LUT_AMPL_WIDTH - 1),
		29591 => to_unsigned(9827, LUT_AMPL_WIDTH - 1),
		29592 => to_unsigned(9824, LUT_AMPL_WIDTH - 1),
		29593 => to_unsigned(9821, LUT_AMPL_WIDTH - 1),
		29594 => to_unsigned(9818, LUT_AMPL_WIDTH - 1),
		29595 => to_unsigned(9815, LUT_AMPL_WIDTH - 1),
		29596 => to_unsigned(9812, LUT_AMPL_WIDTH - 1),
		29597 => to_unsigned(9809, LUT_AMPL_WIDTH - 1),
		29598 => to_unsigned(9806, LUT_AMPL_WIDTH - 1),
		29599 => to_unsigned(9803, LUT_AMPL_WIDTH - 1),
		29600 => to_unsigned(9800, LUT_AMPL_WIDTH - 1),
		29601 => to_unsigned(9797, LUT_AMPL_WIDTH - 1),
		29602 => to_unsigned(9794, LUT_AMPL_WIDTH - 1),
		29603 => to_unsigned(9791, LUT_AMPL_WIDTH - 1),
		29604 => to_unsigned(9788, LUT_AMPL_WIDTH - 1),
		29605 => to_unsigned(9785, LUT_AMPL_WIDTH - 1),
		29606 => to_unsigned(9782, LUT_AMPL_WIDTH - 1),
		29607 => to_unsigned(9779, LUT_AMPL_WIDTH - 1),
		29608 => to_unsigned(9776, LUT_AMPL_WIDTH - 1),
		29609 => to_unsigned(9773, LUT_AMPL_WIDTH - 1),
		29610 => to_unsigned(9770, LUT_AMPL_WIDTH - 1),
		29611 => to_unsigned(9767, LUT_AMPL_WIDTH - 1),
		29612 => to_unsigned(9764, LUT_AMPL_WIDTH - 1),
		29613 => to_unsigned(9761, LUT_AMPL_WIDTH - 1),
		29614 => to_unsigned(9758, LUT_AMPL_WIDTH - 1),
		29615 => to_unsigned(9755, LUT_AMPL_WIDTH - 1),
		29616 => to_unsigned(9752, LUT_AMPL_WIDTH - 1),
		29617 => to_unsigned(9749, LUT_AMPL_WIDTH - 1),
		29618 => to_unsigned(9746, LUT_AMPL_WIDTH - 1),
		29619 => to_unsigned(9743, LUT_AMPL_WIDTH - 1),
		29620 => to_unsigned(9740, LUT_AMPL_WIDTH - 1),
		29621 => to_unsigned(9737, LUT_AMPL_WIDTH - 1),
		29622 => to_unsigned(9734, LUT_AMPL_WIDTH - 1),
		29623 => to_unsigned(9731, LUT_AMPL_WIDTH - 1),
		29624 => to_unsigned(9728, LUT_AMPL_WIDTH - 1),
		29625 => to_unsigned(9725, LUT_AMPL_WIDTH - 1),
		29626 => to_unsigned(9722, LUT_AMPL_WIDTH - 1),
		29627 => to_unsigned(9719, LUT_AMPL_WIDTH - 1),
		29628 => to_unsigned(9716, LUT_AMPL_WIDTH - 1),
		29629 => to_unsigned(9713, LUT_AMPL_WIDTH - 1),
		29630 => to_unsigned(9710, LUT_AMPL_WIDTH - 1),
		29631 => to_unsigned(9707, LUT_AMPL_WIDTH - 1),
		29632 => to_unsigned(9704, LUT_AMPL_WIDTH - 1),
		29633 => to_unsigned(9701, LUT_AMPL_WIDTH - 1),
		29634 => to_unsigned(9698, LUT_AMPL_WIDTH - 1),
		29635 => to_unsigned(9695, LUT_AMPL_WIDTH - 1),
		29636 => to_unsigned(9692, LUT_AMPL_WIDTH - 1),
		29637 => to_unsigned(9689, LUT_AMPL_WIDTH - 1),
		29638 => to_unsigned(9686, LUT_AMPL_WIDTH - 1),
		29639 => to_unsigned(9683, LUT_AMPL_WIDTH - 1),
		29640 => to_unsigned(9680, LUT_AMPL_WIDTH - 1),
		29641 => to_unsigned(9677, LUT_AMPL_WIDTH - 1),
		29642 => to_unsigned(9674, LUT_AMPL_WIDTH - 1),
		29643 => to_unsigned(9671, LUT_AMPL_WIDTH - 1),
		29644 => to_unsigned(9668, LUT_AMPL_WIDTH - 1),
		29645 => to_unsigned(9665, LUT_AMPL_WIDTH - 1),
		29646 => to_unsigned(9662, LUT_AMPL_WIDTH - 1),
		29647 => to_unsigned(9659, LUT_AMPL_WIDTH - 1),
		29648 => to_unsigned(9656, LUT_AMPL_WIDTH - 1),
		29649 => to_unsigned(9653, LUT_AMPL_WIDTH - 1),
		29650 => to_unsigned(9650, LUT_AMPL_WIDTH - 1),
		29651 => to_unsigned(9647, LUT_AMPL_WIDTH - 1),
		29652 => to_unsigned(9644, LUT_AMPL_WIDTH - 1),
		29653 => to_unsigned(9641, LUT_AMPL_WIDTH - 1),
		29654 => to_unsigned(9638, LUT_AMPL_WIDTH - 1),
		29655 => to_unsigned(9635, LUT_AMPL_WIDTH - 1),
		29656 => to_unsigned(9632, LUT_AMPL_WIDTH - 1),
		29657 => to_unsigned(9629, LUT_AMPL_WIDTH - 1),
		29658 => to_unsigned(9626, LUT_AMPL_WIDTH - 1),
		29659 => to_unsigned(9623, LUT_AMPL_WIDTH - 1),
		29660 => to_unsigned(9620, LUT_AMPL_WIDTH - 1),
		29661 => to_unsigned(9617, LUT_AMPL_WIDTH - 1),
		29662 => to_unsigned(9614, LUT_AMPL_WIDTH - 1),
		29663 => to_unsigned(9611, LUT_AMPL_WIDTH - 1),
		29664 => to_unsigned(9608, LUT_AMPL_WIDTH - 1),
		29665 => to_unsigned(9605, LUT_AMPL_WIDTH - 1),
		29666 => to_unsigned(9602, LUT_AMPL_WIDTH - 1),
		29667 => to_unsigned(9599, LUT_AMPL_WIDTH - 1),
		29668 => to_unsigned(9596, LUT_AMPL_WIDTH - 1),
		29669 => to_unsigned(9593, LUT_AMPL_WIDTH - 1),
		29670 => to_unsigned(9590, LUT_AMPL_WIDTH - 1),
		29671 => to_unsigned(9587, LUT_AMPL_WIDTH - 1),
		29672 => to_unsigned(9584, LUT_AMPL_WIDTH - 1),
		29673 => to_unsigned(9581, LUT_AMPL_WIDTH - 1),
		29674 => to_unsigned(9578, LUT_AMPL_WIDTH - 1),
		29675 => to_unsigned(9575, LUT_AMPL_WIDTH - 1),
		29676 => to_unsigned(9572, LUT_AMPL_WIDTH - 1),
		29677 => to_unsigned(9569, LUT_AMPL_WIDTH - 1),
		29678 => to_unsigned(9566, LUT_AMPL_WIDTH - 1),
		29679 => to_unsigned(9563, LUT_AMPL_WIDTH - 1),
		29680 => to_unsigned(9560, LUT_AMPL_WIDTH - 1),
		29681 => to_unsigned(9557, LUT_AMPL_WIDTH - 1),
		29682 => to_unsigned(9554, LUT_AMPL_WIDTH - 1),
		29683 => to_unsigned(9551, LUT_AMPL_WIDTH - 1),
		29684 => to_unsigned(9548, LUT_AMPL_WIDTH - 1),
		29685 => to_unsigned(9545, LUT_AMPL_WIDTH - 1),
		29686 => to_unsigned(9542, LUT_AMPL_WIDTH - 1),
		29687 => to_unsigned(9539, LUT_AMPL_WIDTH - 1),
		29688 => to_unsigned(9536, LUT_AMPL_WIDTH - 1),
		29689 => to_unsigned(9533, LUT_AMPL_WIDTH - 1),
		29690 => to_unsigned(9530, LUT_AMPL_WIDTH - 1),
		29691 => to_unsigned(9527, LUT_AMPL_WIDTH - 1),
		29692 => to_unsigned(9524, LUT_AMPL_WIDTH - 1),
		29693 => to_unsigned(9521, LUT_AMPL_WIDTH - 1),
		29694 => to_unsigned(9518, LUT_AMPL_WIDTH - 1),
		29695 => to_unsigned(9515, LUT_AMPL_WIDTH - 1),
		29696 => to_unsigned(9512, LUT_AMPL_WIDTH - 1),
		29697 => to_unsigned(9509, LUT_AMPL_WIDTH - 1),
		29698 => to_unsigned(9506, LUT_AMPL_WIDTH - 1),
		29699 => to_unsigned(9503, LUT_AMPL_WIDTH - 1),
		29700 => to_unsigned(9500, LUT_AMPL_WIDTH - 1),
		29701 => to_unsigned(9497, LUT_AMPL_WIDTH - 1),
		29702 => to_unsigned(9494, LUT_AMPL_WIDTH - 1),
		29703 => to_unsigned(9491, LUT_AMPL_WIDTH - 1),
		29704 => to_unsigned(9488, LUT_AMPL_WIDTH - 1),
		29705 => to_unsigned(9485, LUT_AMPL_WIDTH - 1),
		29706 => to_unsigned(9482, LUT_AMPL_WIDTH - 1),
		29707 => to_unsigned(9479, LUT_AMPL_WIDTH - 1),
		29708 => to_unsigned(9476, LUT_AMPL_WIDTH - 1),
		29709 => to_unsigned(9473, LUT_AMPL_WIDTH - 1),
		29710 => to_unsigned(9470, LUT_AMPL_WIDTH - 1),
		29711 => to_unsigned(9467, LUT_AMPL_WIDTH - 1),
		29712 => to_unsigned(9464, LUT_AMPL_WIDTH - 1),
		29713 => to_unsigned(9461, LUT_AMPL_WIDTH - 1),
		29714 => to_unsigned(9458, LUT_AMPL_WIDTH - 1),
		29715 => to_unsigned(9455, LUT_AMPL_WIDTH - 1),
		29716 => to_unsigned(9452, LUT_AMPL_WIDTH - 1),
		29717 => to_unsigned(9449, LUT_AMPL_WIDTH - 1),
		29718 => to_unsigned(9446, LUT_AMPL_WIDTH - 1),
		29719 => to_unsigned(9443, LUT_AMPL_WIDTH - 1),
		29720 => to_unsigned(9440, LUT_AMPL_WIDTH - 1),
		29721 => to_unsigned(9437, LUT_AMPL_WIDTH - 1),
		29722 => to_unsigned(9434, LUT_AMPL_WIDTH - 1),
		29723 => to_unsigned(9431, LUT_AMPL_WIDTH - 1),
		29724 => to_unsigned(9428, LUT_AMPL_WIDTH - 1),
		29725 => to_unsigned(9425, LUT_AMPL_WIDTH - 1),
		29726 => to_unsigned(9422, LUT_AMPL_WIDTH - 1),
		29727 => to_unsigned(9419, LUT_AMPL_WIDTH - 1),
		29728 => to_unsigned(9416, LUT_AMPL_WIDTH - 1),
		29729 => to_unsigned(9413, LUT_AMPL_WIDTH - 1),
		29730 => to_unsigned(9409, LUT_AMPL_WIDTH - 1),
		29731 => to_unsigned(9406, LUT_AMPL_WIDTH - 1),
		29732 => to_unsigned(9403, LUT_AMPL_WIDTH - 1),
		29733 => to_unsigned(9400, LUT_AMPL_WIDTH - 1),
		29734 => to_unsigned(9397, LUT_AMPL_WIDTH - 1),
		29735 => to_unsigned(9394, LUT_AMPL_WIDTH - 1),
		29736 => to_unsigned(9391, LUT_AMPL_WIDTH - 1),
		29737 => to_unsigned(9388, LUT_AMPL_WIDTH - 1),
		29738 => to_unsigned(9385, LUT_AMPL_WIDTH - 1),
		29739 => to_unsigned(9382, LUT_AMPL_WIDTH - 1),
		29740 => to_unsigned(9379, LUT_AMPL_WIDTH - 1),
		29741 => to_unsigned(9376, LUT_AMPL_WIDTH - 1),
		29742 => to_unsigned(9373, LUT_AMPL_WIDTH - 1),
		29743 => to_unsigned(9370, LUT_AMPL_WIDTH - 1),
		29744 => to_unsigned(9367, LUT_AMPL_WIDTH - 1),
		29745 => to_unsigned(9364, LUT_AMPL_WIDTH - 1),
		29746 => to_unsigned(9361, LUT_AMPL_WIDTH - 1),
		29747 => to_unsigned(9358, LUT_AMPL_WIDTH - 1),
		29748 => to_unsigned(9355, LUT_AMPL_WIDTH - 1),
		29749 => to_unsigned(9352, LUT_AMPL_WIDTH - 1),
		29750 => to_unsigned(9349, LUT_AMPL_WIDTH - 1),
		29751 => to_unsigned(9346, LUT_AMPL_WIDTH - 1),
		29752 => to_unsigned(9343, LUT_AMPL_WIDTH - 1),
		29753 => to_unsigned(9340, LUT_AMPL_WIDTH - 1),
		29754 => to_unsigned(9337, LUT_AMPL_WIDTH - 1),
		29755 => to_unsigned(9334, LUT_AMPL_WIDTH - 1),
		29756 => to_unsigned(9331, LUT_AMPL_WIDTH - 1),
		29757 => to_unsigned(9328, LUT_AMPL_WIDTH - 1),
		29758 => to_unsigned(9325, LUT_AMPL_WIDTH - 1),
		29759 => to_unsigned(9322, LUT_AMPL_WIDTH - 1),
		29760 => to_unsigned(9319, LUT_AMPL_WIDTH - 1),
		29761 => to_unsigned(9316, LUT_AMPL_WIDTH - 1),
		29762 => to_unsigned(9313, LUT_AMPL_WIDTH - 1),
		29763 => to_unsigned(9310, LUT_AMPL_WIDTH - 1),
		29764 => to_unsigned(9307, LUT_AMPL_WIDTH - 1),
		29765 => to_unsigned(9304, LUT_AMPL_WIDTH - 1),
		29766 => to_unsigned(9301, LUT_AMPL_WIDTH - 1),
		29767 => to_unsigned(9298, LUT_AMPL_WIDTH - 1),
		29768 => to_unsigned(9295, LUT_AMPL_WIDTH - 1),
		29769 => to_unsigned(9292, LUT_AMPL_WIDTH - 1),
		29770 => to_unsigned(9289, LUT_AMPL_WIDTH - 1),
		29771 => to_unsigned(9286, LUT_AMPL_WIDTH - 1),
		29772 => to_unsigned(9283, LUT_AMPL_WIDTH - 1),
		29773 => to_unsigned(9280, LUT_AMPL_WIDTH - 1),
		29774 => to_unsigned(9277, LUT_AMPL_WIDTH - 1),
		29775 => to_unsigned(9274, LUT_AMPL_WIDTH - 1),
		29776 => to_unsigned(9271, LUT_AMPL_WIDTH - 1),
		29777 => to_unsigned(9268, LUT_AMPL_WIDTH - 1),
		29778 => to_unsigned(9265, LUT_AMPL_WIDTH - 1),
		29779 => to_unsigned(9262, LUT_AMPL_WIDTH - 1),
		29780 => to_unsigned(9259, LUT_AMPL_WIDTH - 1),
		29781 => to_unsigned(9256, LUT_AMPL_WIDTH - 1),
		29782 => to_unsigned(9253, LUT_AMPL_WIDTH - 1),
		29783 => to_unsigned(9250, LUT_AMPL_WIDTH - 1),
		29784 => to_unsigned(9247, LUT_AMPL_WIDTH - 1),
		29785 => to_unsigned(9244, LUT_AMPL_WIDTH - 1),
		29786 => to_unsigned(9241, LUT_AMPL_WIDTH - 1),
		29787 => to_unsigned(9238, LUT_AMPL_WIDTH - 1),
		29788 => to_unsigned(9235, LUT_AMPL_WIDTH - 1),
		29789 => to_unsigned(9232, LUT_AMPL_WIDTH - 1),
		29790 => to_unsigned(9229, LUT_AMPL_WIDTH - 1),
		29791 => to_unsigned(9226, LUT_AMPL_WIDTH - 1),
		29792 => to_unsigned(9223, LUT_AMPL_WIDTH - 1),
		29793 => to_unsigned(9220, LUT_AMPL_WIDTH - 1),
		29794 => to_unsigned(9217, LUT_AMPL_WIDTH - 1),
		29795 => to_unsigned(9214, LUT_AMPL_WIDTH - 1),
		29796 => to_unsigned(9211, LUT_AMPL_WIDTH - 1),
		29797 => to_unsigned(9208, LUT_AMPL_WIDTH - 1),
		29798 => to_unsigned(9205, LUT_AMPL_WIDTH - 1),
		29799 => to_unsigned(9202, LUT_AMPL_WIDTH - 1),
		29800 => to_unsigned(9199, LUT_AMPL_WIDTH - 1),
		29801 => to_unsigned(9196, LUT_AMPL_WIDTH - 1),
		29802 => to_unsigned(9193, LUT_AMPL_WIDTH - 1),
		29803 => to_unsigned(9190, LUT_AMPL_WIDTH - 1),
		29804 => to_unsigned(9187, LUT_AMPL_WIDTH - 1),
		29805 => to_unsigned(9184, LUT_AMPL_WIDTH - 1),
		29806 => to_unsigned(9181, LUT_AMPL_WIDTH - 1),
		29807 => to_unsigned(9178, LUT_AMPL_WIDTH - 1),
		29808 => to_unsigned(9175, LUT_AMPL_WIDTH - 1),
		29809 => to_unsigned(9172, LUT_AMPL_WIDTH - 1),
		29810 => to_unsigned(9168, LUT_AMPL_WIDTH - 1),
		29811 => to_unsigned(9165, LUT_AMPL_WIDTH - 1),
		29812 => to_unsigned(9162, LUT_AMPL_WIDTH - 1),
		29813 => to_unsigned(9159, LUT_AMPL_WIDTH - 1),
		29814 => to_unsigned(9156, LUT_AMPL_WIDTH - 1),
		29815 => to_unsigned(9153, LUT_AMPL_WIDTH - 1),
		29816 => to_unsigned(9150, LUT_AMPL_WIDTH - 1),
		29817 => to_unsigned(9147, LUT_AMPL_WIDTH - 1),
		29818 => to_unsigned(9144, LUT_AMPL_WIDTH - 1),
		29819 => to_unsigned(9141, LUT_AMPL_WIDTH - 1),
		29820 => to_unsigned(9138, LUT_AMPL_WIDTH - 1),
		29821 => to_unsigned(9135, LUT_AMPL_WIDTH - 1),
		29822 => to_unsigned(9132, LUT_AMPL_WIDTH - 1),
		29823 => to_unsigned(9129, LUT_AMPL_WIDTH - 1),
		29824 => to_unsigned(9126, LUT_AMPL_WIDTH - 1),
		29825 => to_unsigned(9123, LUT_AMPL_WIDTH - 1),
		29826 => to_unsigned(9120, LUT_AMPL_WIDTH - 1),
		29827 => to_unsigned(9117, LUT_AMPL_WIDTH - 1),
		29828 => to_unsigned(9114, LUT_AMPL_WIDTH - 1),
		29829 => to_unsigned(9111, LUT_AMPL_WIDTH - 1),
		29830 => to_unsigned(9108, LUT_AMPL_WIDTH - 1),
		29831 => to_unsigned(9105, LUT_AMPL_WIDTH - 1),
		29832 => to_unsigned(9102, LUT_AMPL_WIDTH - 1),
		29833 => to_unsigned(9099, LUT_AMPL_WIDTH - 1),
		29834 => to_unsigned(9096, LUT_AMPL_WIDTH - 1),
		29835 => to_unsigned(9093, LUT_AMPL_WIDTH - 1),
		29836 => to_unsigned(9090, LUT_AMPL_WIDTH - 1),
		29837 => to_unsigned(9087, LUT_AMPL_WIDTH - 1),
		29838 => to_unsigned(9084, LUT_AMPL_WIDTH - 1),
		29839 => to_unsigned(9081, LUT_AMPL_WIDTH - 1),
		29840 => to_unsigned(9078, LUT_AMPL_WIDTH - 1),
		29841 => to_unsigned(9075, LUT_AMPL_WIDTH - 1),
		29842 => to_unsigned(9072, LUT_AMPL_WIDTH - 1),
		29843 => to_unsigned(9069, LUT_AMPL_WIDTH - 1),
		29844 => to_unsigned(9066, LUT_AMPL_WIDTH - 1),
		29845 => to_unsigned(9063, LUT_AMPL_WIDTH - 1),
		29846 => to_unsigned(9060, LUT_AMPL_WIDTH - 1),
		29847 => to_unsigned(9057, LUT_AMPL_WIDTH - 1),
		29848 => to_unsigned(9054, LUT_AMPL_WIDTH - 1),
		29849 => to_unsigned(9051, LUT_AMPL_WIDTH - 1),
		29850 => to_unsigned(9048, LUT_AMPL_WIDTH - 1),
		29851 => to_unsigned(9045, LUT_AMPL_WIDTH - 1),
		29852 => to_unsigned(9042, LUT_AMPL_WIDTH - 1),
		29853 => to_unsigned(9039, LUT_AMPL_WIDTH - 1),
		29854 => to_unsigned(9036, LUT_AMPL_WIDTH - 1),
		29855 => to_unsigned(9033, LUT_AMPL_WIDTH - 1),
		29856 => to_unsigned(9030, LUT_AMPL_WIDTH - 1),
		29857 => to_unsigned(9027, LUT_AMPL_WIDTH - 1),
		29858 => to_unsigned(9024, LUT_AMPL_WIDTH - 1),
		29859 => to_unsigned(9021, LUT_AMPL_WIDTH - 1),
		29860 => to_unsigned(9018, LUT_AMPL_WIDTH - 1),
		29861 => to_unsigned(9015, LUT_AMPL_WIDTH - 1),
		29862 => to_unsigned(9012, LUT_AMPL_WIDTH - 1),
		29863 => to_unsigned(9009, LUT_AMPL_WIDTH - 1),
		29864 => to_unsigned(9006, LUT_AMPL_WIDTH - 1),
		29865 => to_unsigned(9002, LUT_AMPL_WIDTH - 1),
		29866 => to_unsigned(8999, LUT_AMPL_WIDTH - 1),
		29867 => to_unsigned(8996, LUT_AMPL_WIDTH - 1),
		29868 => to_unsigned(8993, LUT_AMPL_WIDTH - 1),
		29869 => to_unsigned(8990, LUT_AMPL_WIDTH - 1),
		29870 => to_unsigned(8987, LUT_AMPL_WIDTH - 1),
		29871 => to_unsigned(8984, LUT_AMPL_WIDTH - 1),
		29872 => to_unsigned(8981, LUT_AMPL_WIDTH - 1),
		29873 => to_unsigned(8978, LUT_AMPL_WIDTH - 1),
		29874 => to_unsigned(8975, LUT_AMPL_WIDTH - 1),
		29875 => to_unsigned(8972, LUT_AMPL_WIDTH - 1),
		29876 => to_unsigned(8969, LUT_AMPL_WIDTH - 1),
		29877 => to_unsigned(8966, LUT_AMPL_WIDTH - 1),
		29878 => to_unsigned(8963, LUT_AMPL_WIDTH - 1),
		29879 => to_unsigned(8960, LUT_AMPL_WIDTH - 1),
		29880 => to_unsigned(8957, LUT_AMPL_WIDTH - 1),
		29881 => to_unsigned(8954, LUT_AMPL_WIDTH - 1),
		29882 => to_unsigned(8951, LUT_AMPL_WIDTH - 1),
		29883 => to_unsigned(8948, LUT_AMPL_WIDTH - 1),
		29884 => to_unsigned(8945, LUT_AMPL_WIDTH - 1),
		29885 => to_unsigned(8942, LUT_AMPL_WIDTH - 1),
		29886 => to_unsigned(8939, LUT_AMPL_WIDTH - 1),
		29887 => to_unsigned(8936, LUT_AMPL_WIDTH - 1),
		29888 => to_unsigned(8933, LUT_AMPL_WIDTH - 1),
		29889 => to_unsigned(8930, LUT_AMPL_WIDTH - 1),
		29890 => to_unsigned(8927, LUT_AMPL_WIDTH - 1),
		29891 => to_unsigned(8924, LUT_AMPL_WIDTH - 1),
		29892 => to_unsigned(8921, LUT_AMPL_WIDTH - 1),
		29893 => to_unsigned(8918, LUT_AMPL_WIDTH - 1),
		29894 => to_unsigned(8915, LUT_AMPL_WIDTH - 1),
		29895 => to_unsigned(8912, LUT_AMPL_WIDTH - 1),
		29896 => to_unsigned(8909, LUT_AMPL_WIDTH - 1),
		29897 => to_unsigned(8906, LUT_AMPL_WIDTH - 1),
		29898 => to_unsigned(8903, LUT_AMPL_WIDTH - 1),
		29899 => to_unsigned(8900, LUT_AMPL_WIDTH - 1),
		29900 => to_unsigned(8897, LUT_AMPL_WIDTH - 1),
		29901 => to_unsigned(8894, LUT_AMPL_WIDTH - 1),
		29902 => to_unsigned(8891, LUT_AMPL_WIDTH - 1),
		29903 => to_unsigned(8888, LUT_AMPL_WIDTH - 1),
		29904 => to_unsigned(8885, LUT_AMPL_WIDTH - 1),
		29905 => to_unsigned(8882, LUT_AMPL_WIDTH - 1),
		29906 => to_unsigned(8879, LUT_AMPL_WIDTH - 1),
		29907 => to_unsigned(8876, LUT_AMPL_WIDTH - 1),
		29908 => to_unsigned(8873, LUT_AMPL_WIDTH - 1),
		29909 => to_unsigned(8869, LUT_AMPL_WIDTH - 1),
		29910 => to_unsigned(8866, LUT_AMPL_WIDTH - 1),
		29911 => to_unsigned(8863, LUT_AMPL_WIDTH - 1),
		29912 => to_unsigned(8860, LUT_AMPL_WIDTH - 1),
		29913 => to_unsigned(8857, LUT_AMPL_WIDTH - 1),
		29914 => to_unsigned(8854, LUT_AMPL_WIDTH - 1),
		29915 => to_unsigned(8851, LUT_AMPL_WIDTH - 1),
		29916 => to_unsigned(8848, LUT_AMPL_WIDTH - 1),
		29917 => to_unsigned(8845, LUT_AMPL_WIDTH - 1),
		29918 => to_unsigned(8842, LUT_AMPL_WIDTH - 1),
		29919 => to_unsigned(8839, LUT_AMPL_WIDTH - 1),
		29920 => to_unsigned(8836, LUT_AMPL_WIDTH - 1),
		29921 => to_unsigned(8833, LUT_AMPL_WIDTH - 1),
		29922 => to_unsigned(8830, LUT_AMPL_WIDTH - 1),
		29923 => to_unsigned(8827, LUT_AMPL_WIDTH - 1),
		29924 => to_unsigned(8824, LUT_AMPL_WIDTH - 1),
		29925 => to_unsigned(8821, LUT_AMPL_WIDTH - 1),
		29926 => to_unsigned(8818, LUT_AMPL_WIDTH - 1),
		29927 => to_unsigned(8815, LUT_AMPL_WIDTH - 1),
		29928 => to_unsigned(8812, LUT_AMPL_WIDTH - 1),
		29929 => to_unsigned(8809, LUT_AMPL_WIDTH - 1),
		29930 => to_unsigned(8806, LUT_AMPL_WIDTH - 1),
		29931 => to_unsigned(8803, LUT_AMPL_WIDTH - 1),
		29932 => to_unsigned(8800, LUT_AMPL_WIDTH - 1),
		29933 => to_unsigned(8797, LUT_AMPL_WIDTH - 1),
		29934 => to_unsigned(8794, LUT_AMPL_WIDTH - 1),
		29935 => to_unsigned(8791, LUT_AMPL_WIDTH - 1),
		29936 => to_unsigned(8788, LUT_AMPL_WIDTH - 1),
		29937 => to_unsigned(8785, LUT_AMPL_WIDTH - 1),
		29938 => to_unsigned(8782, LUT_AMPL_WIDTH - 1),
		29939 => to_unsigned(8779, LUT_AMPL_WIDTH - 1),
		29940 => to_unsigned(8776, LUT_AMPL_WIDTH - 1),
		29941 => to_unsigned(8773, LUT_AMPL_WIDTH - 1),
		29942 => to_unsigned(8770, LUT_AMPL_WIDTH - 1),
		29943 => to_unsigned(8767, LUT_AMPL_WIDTH - 1),
		29944 => to_unsigned(8764, LUT_AMPL_WIDTH - 1),
		29945 => to_unsigned(8761, LUT_AMPL_WIDTH - 1),
		29946 => to_unsigned(8758, LUT_AMPL_WIDTH - 1),
		29947 => to_unsigned(8755, LUT_AMPL_WIDTH - 1),
		29948 => to_unsigned(8751, LUT_AMPL_WIDTH - 1),
		29949 => to_unsigned(8748, LUT_AMPL_WIDTH - 1),
		29950 => to_unsigned(8745, LUT_AMPL_WIDTH - 1),
		29951 => to_unsigned(8742, LUT_AMPL_WIDTH - 1),
		29952 => to_unsigned(8739, LUT_AMPL_WIDTH - 1),
		29953 => to_unsigned(8736, LUT_AMPL_WIDTH - 1),
		29954 => to_unsigned(8733, LUT_AMPL_WIDTH - 1),
		29955 => to_unsigned(8730, LUT_AMPL_WIDTH - 1),
		29956 => to_unsigned(8727, LUT_AMPL_WIDTH - 1),
		29957 => to_unsigned(8724, LUT_AMPL_WIDTH - 1),
		29958 => to_unsigned(8721, LUT_AMPL_WIDTH - 1),
		29959 => to_unsigned(8718, LUT_AMPL_WIDTH - 1),
		29960 => to_unsigned(8715, LUT_AMPL_WIDTH - 1),
		29961 => to_unsigned(8712, LUT_AMPL_WIDTH - 1),
		29962 => to_unsigned(8709, LUT_AMPL_WIDTH - 1),
		29963 => to_unsigned(8706, LUT_AMPL_WIDTH - 1),
		29964 => to_unsigned(8703, LUT_AMPL_WIDTH - 1),
		29965 => to_unsigned(8700, LUT_AMPL_WIDTH - 1),
		29966 => to_unsigned(8697, LUT_AMPL_WIDTH - 1),
		29967 => to_unsigned(8694, LUT_AMPL_WIDTH - 1),
		29968 => to_unsigned(8691, LUT_AMPL_WIDTH - 1),
		29969 => to_unsigned(8688, LUT_AMPL_WIDTH - 1),
		29970 => to_unsigned(8685, LUT_AMPL_WIDTH - 1),
		29971 => to_unsigned(8682, LUT_AMPL_WIDTH - 1),
		29972 => to_unsigned(8679, LUT_AMPL_WIDTH - 1),
		29973 => to_unsigned(8676, LUT_AMPL_WIDTH - 1),
		29974 => to_unsigned(8673, LUT_AMPL_WIDTH - 1),
		29975 => to_unsigned(8670, LUT_AMPL_WIDTH - 1),
		29976 => to_unsigned(8667, LUT_AMPL_WIDTH - 1),
		29977 => to_unsigned(8664, LUT_AMPL_WIDTH - 1),
		29978 => to_unsigned(8661, LUT_AMPL_WIDTH - 1),
		29979 => to_unsigned(8658, LUT_AMPL_WIDTH - 1),
		29980 => to_unsigned(8655, LUT_AMPL_WIDTH - 1),
		29981 => to_unsigned(8652, LUT_AMPL_WIDTH - 1),
		29982 => to_unsigned(8649, LUT_AMPL_WIDTH - 1),
		29983 => to_unsigned(8645, LUT_AMPL_WIDTH - 1),
		29984 => to_unsigned(8642, LUT_AMPL_WIDTH - 1),
		29985 => to_unsigned(8639, LUT_AMPL_WIDTH - 1),
		29986 => to_unsigned(8636, LUT_AMPL_WIDTH - 1),
		29987 => to_unsigned(8633, LUT_AMPL_WIDTH - 1),
		29988 => to_unsigned(8630, LUT_AMPL_WIDTH - 1),
		29989 => to_unsigned(8627, LUT_AMPL_WIDTH - 1),
		29990 => to_unsigned(8624, LUT_AMPL_WIDTH - 1),
		29991 => to_unsigned(8621, LUT_AMPL_WIDTH - 1),
		29992 => to_unsigned(8618, LUT_AMPL_WIDTH - 1),
		29993 => to_unsigned(8615, LUT_AMPL_WIDTH - 1),
		29994 => to_unsigned(8612, LUT_AMPL_WIDTH - 1),
		29995 => to_unsigned(8609, LUT_AMPL_WIDTH - 1),
		29996 => to_unsigned(8606, LUT_AMPL_WIDTH - 1),
		29997 => to_unsigned(8603, LUT_AMPL_WIDTH - 1),
		29998 => to_unsigned(8600, LUT_AMPL_WIDTH - 1),
		29999 => to_unsigned(8597, LUT_AMPL_WIDTH - 1),
		30000 => to_unsigned(8594, LUT_AMPL_WIDTH - 1),
		30001 => to_unsigned(8591, LUT_AMPL_WIDTH - 1),
		30002 => to_unsigned(8588, LUT_AMPL_WIDTH - 1),
		30003 => to_unsigned(8585, LUT_AMPL_WIDTH - 1),
		30004 => to_unsigned(8582, LUT_AMPL_WIDTH - 1),
		30005 => to_unsigned(8579, LUT_AMPL_WIDTH - 1),
		30006 => to_unsigned(8576, LUT_AMPL_WIDTH - 1),
		30007 => to_unsigned(8573, LUT_AMPL_WIDTH - 1),
		30008 => to_unsigned(8570, LUT_AMPL_WIDTH - 1),
		30009 => to_unsigned(8567, LUT_AMPL_WIDTH - 1),
		30010 => to_unsigned(8564, LUT_AMPL_WIDTH - 1),
		30011 => to_unsigned(8561, LUT_AMPL_WIDTH - 1),
		30012 => to_unsigned(8558, LUT_AMPL_WIDTH - 1),
		30013 => to_unsigned(8555, LUT_AMPL_WIDTH - 1),
		30014 => to_unsigned(8552, LUT_AMPL_WIDTH - 1),
		30015 => to_unsigned(8548, LUT_AMPL_WIDTH - 1),
		30016 => to_unsigned(8545, LUT_AMPL_WIDTH - 1),
		30017 => to_unsigned(8542, LUT_AMPL_WIDTH - 1),
		30018 => to_unsigned(8539, LUT_AMPL_WIDTH - 1),
		30019 => to_unsigned(8536, LUT_AMPL_WIDTH - 1),
		30020 => to_unsigned(8533, LUT_AMPL_WIDTH - 1),
		30021 => to_unsigned(8530, LUT_AMPL_WIDTH - 1),
		30022 => to_unsigned(8527, LUT_AMPL_WIDTH - 1),
		30023 => to_unsigned(8524, LUT_AMPL_WIDTH - 1),
		30024 => to_unsigned(8521, LUT_AMPL_WIDTH - 1),
		30025 => to_unsigned(8518, LUT_AMPL_WIDTH - 1),
		30026 => to_unsigned(8515, LUT_AMPL_WIDTH - 1),
		30027 => to_unsigned(8512, LUT_AMPL_WIDTH - 1),
		30028 => to_unsigned(8509, LUT_AMPL_WIDTH - 1),
		30029 => to_unsigned(8506, LUT_AMPL_WIDTH - 1),
		30030 => to_unsigned(8503, LUT_AMPL_WIDTH - 1),
		30031 => to_unsigned(8500, LUT_AMPL_WIDTH - 1),
		30032 => to_unsigned(8497, LUT_AMPL_WIDTH - 1),
		30033 => to_unsigned(8494, LUT_AMPL_WIDTH - 1),
		30034 => to_unsigned(8491, LUT_AMPL_WIDTH - 1),
		30035 => to_unsigned(8488, LUT_AMPL_WIDTH - 1),
		30036 => to_unsigned(8485, LUT_AMPL_WIDTH - 1),
		30037 => to_unsigned(8482, LUT_AMPL_WIDTH - 1),
		30038 => to_unsigned(8479, LUT_AMPL_WIDTH - 1),
		30039 => to_unsigned(8476, LUT_AMPL_WIDTH - 1),
		30040 => to_unsigned(8473, LUT_AMPL_WIDTH - 1),
		30041 => to_unsigned(8470, LUT_AMPL_WIDTH - 1),
		30042 => to_unsigned(8467, LUT_AMPL_WIDTH - 1),
		30043 => to_unsigned(8464, LUT_AMPL_WIDTH - 1),
		30044 => to_unsigned(8460, LUT_AMPL_WIDTH - 1),
		30045 => to_unsigned(8457, LUT_AMPL_WIDTH - 1),
		30046 => to_unsigned(8454, LUT_AMPL_WIDTH - 1),
		30047 => to_unsigned(8451, LUT_AMPL_WIDTH - 1),
		30048 => to_unsigned(8448, LUT_AMPL_WIDTH - 1),
		30049 => to_unsigned(8445, LUT_AMPL_WIDTH - 1),
		30050 => to_unsigned(8442, LUT_AMPL_WIDTH - 1),
		30051 => to_unsigned(8439, LUT_AMPL_WIDTH - 1),
		30052 => to_unsigned(8436, LUT_AMPL_WIDTH - 1),
		30053 => to_unsigned(8433, LUT_AMPL_WIDTH - 1),
		30054 => to_unsigned(8430, LUT_AMPL_WIDTH - 1),
		30055 => to_unsigned(8427, LUT_AMPL_WIDTH - 1),
		30056 => to_unsigned(8424, LUT_AMPL_WIDTH - 1),
		30057 => to_unsigned(8421, LUT_AMPL_WIDTH - 1),
		30058 => to_unsigned(8418, LUT_AMPL_WIDTH - 1),
		30059 => to_unsigned(8415, LUT_AMPL_WIDTH - 1),
		30060 => to_unsigned(8412, LUT_AMPL_WIDTH - 1),
		30061 => to_unsigned(8409, LUT_AMPL_WIDTH - 1),
		30062 => to_unsigned(8406, LUT_AMPL_WIDTH - 1),
		30063 => to_unsigned(8403, LUT_AMPL_WIDTH - 1),
		30064 => to_unsigned(8400, LUT_AMPL_WIDTH - 1),
		30065 => to_unsigned(8397, LUT_AMPL_WIDTH - 1),
		30066 => to_unsigned(8394, LUT_AMPL_WIDTH - 1),
		30067 => to_unsigned(8391, LUT_AMPL_WIDTH - 1),
		30068 => to_unsigned(8388, LUT_AMPL_WIDTH - 1),
		30069 => to_unsigned(8385, LUT_AMPL_WIDTH - 1),
		30070 => to_unsigned(8382, LUT_AMPL_WIDTH - 1),
		30071 => to_unsigned(8379, LUT_AMPL_WIDTH - 1),
		30072 => to_unsigned(8375, LUT_AMPL_WIDTH - 1),
		30073 => to_unsigned(8372, LUT_AMPL_WIDTH - 1),
		30074 => to_unsigned(8369, LUT_AMPL_WIDTH - 1),
		30075 => to_unsigned(8366, LUT_AMPL_WIDTH - 1),
		30076 => to_unsigned(8363, LUT_AMPL_WIDTH - 1),
		30077 => to_unsigned(8360, LUT_AMPL_WIDTH - 1),
		30078 => to_unsigned(8357, LUT_AMPL_WIDTH - 1),
		30079 => to_unsigned(8354, LUT_AMPL_WIDTH - 1),
		30080 => to_unsigned(8351, LUT_AMPL_WIDTH - 1),
		30081 => to_unsigned(8348, LUT_AMPL_WIDTH - 1),
		30082 => to_unsigned(8345, LUT_AMPL_WIDTH - 1),
		30083 => to_unsigned(8342, LUT_AMPL_WIDTH - 1),
		30084 => to_unsigned(8339, LUT_AMPL_WIDTH - 1),
		30085 => to_unsigned(8336, LUT_AMPL_WIDTH - 1),
		30086 => to_unsigned(8333, LUT_AMPL_WIDTH - 1),
		30087 => to_unsigned(8330, LUT_AMPL_WIDTH - 1),
		30088 => to_unsigned(8327, LUT_AMPL_WIDTH - 1),
		30089 => to_unsigned(8324, LUT_AMPL_WIDTH - 1),
		30090 => to_unsigned(8321, LUT_AMPL_WIDTH - 1),
		30091 => to_unsigned(8318, LUT_AMPL_WIDTH - 1),
		30092 => to_unsigned(8315, LUT_AMPL_WIDTH - 1),
		30093 => to_unsigned(8312, LUT_AMPL_WIDTH - 1),
		30094 => to_unsigned(8309, LUT_AMPL_WIDTH - 1),
		30095 => to_unsigned(8306, LUT_AMPL_WIDTH - 1),
		30096 => to_unsigned(8303, LUT_AMPL_WIDTH - 1),
		30097 => to_unsigned(8300, LUT_AMPL_WIDTH - 1),
		30098 => to_unsigned(8296, LUT_AMPL_WIDTH - 1),
		30099 => to_unsigned(8293, LUT_AMPL_WIDTH - 1),
		30100 => to_unsigned(8290, LUT_AMPL_WIDTH - 1),
		30101 => to_unsigned(8287, LUT_AMPL_WIDTH - 1),
		30102 => to_unsigned(8284, LUT_AMPL_WIDTH - 1),
		30103 => to_unsigned(8281, LUT_AMPL_WIDTH - 1),
		30104 => to_unsigned(8278, LUT_AMPL_WIDTH - 1),
		30105 => to_unsigned(8275, LUT_AMPL_WIDTH - 1),
		30106 => to_unsigned(8272, LUT_AMPL_WIDTH - 1),
		30107 => to_unsigned(8269, LUT_AMPL_WIDTH - 1),
		30108 => to_unsigned(8266, LUT_AMPL_WIDTH - 1),
		30109 => to_unsigned(8263, LUT_AMPL_WIDTH - 1),
		30110 => to_unsigned(8260, LUT_AMPL_WIDTH - 1),
		30111 => to_unsigned(8257, LUT_AMPL_WIDTH - 1),
		30112 => to_unsigned(8254, LUT_AMPL_WIDTH - 1),
		30113 => to_unsigned(8251, LUT_AMPL_WIDTH - 1),
		30114 => to_unsigned(8248, LUT_AMPL_WIDTH - 1),
		30115 => to_unsigned(8245, LUT_AMPL_WIDTH - 1),
		30116 => to_unsigned(8242, LUT_AMPL_WIDTH - 1),
		30117 => to_unsigned(8239, LUT_AMPL_WIDTH - 1),
		30118 => to_unsigned(8236, LUT_AMPL_WIDTH - 1),
		30119 => to_unsigned(8233, LUT_AMPL_WIDTH - 1),
		30120 => to_unsigned(8230, LUT_AMPL_WIDTH - 1),
		30121 => to_unsigned(8227, LUT_AMPL_WIDTH - 1),
		30122 => to_unsigned(8224, LUT_AMPL_WIDTH - 1),
		30123 => to_unsigned(8220, LUT_AMPL_WIDTH - 1),
		30124 => to_unsigned(8217, LUT_AMPL_WIDTH - 1),
		30125 => to_unsigned(8214, LUT_AMPL_WIDTH - 1),
		30126 => to_unsigned(8211, LUT_AMPL_WIDTH - 1),
		30127 => to_unsigned(8208, LUT_AMPL_WIDTH - 1),
		30128 => to_unsigned(8205, LUT_AMPL_WIDTH - 1),
		30129 => to_unsigned(8202, LUT_AMPL_WIDTH - 1),
		30130 => to_unsigned(8199, LUT_AMPL_WIDTH - 1),
		30131 => to_unsigned(8196, LUT_AMPL_WIDTH - 1),
		30132 => to_unsigned(8193, LUT_AMPL_WIDTH - 1),
		30133 => to_unsigned(8190, LUT_AMPL_WIDTH - 1),
		30134 => to_unsigned(8187, LUT_AMPL_WIDTH - 1),
		30135 => to_unsigned(8184, LUT_AMPL_WIDTH - 1),
		30136 => to_unsigned(8181, LUT_AMPL_WIDTH - 1),
		30137 => to_unsigned(8178, LUT_AMPL_WIDTH - 1),
		30138 => to_unsigned(8175, LUT_AMPL_WIDTH - 1),
		30139 => to_unsigned(8172, LUT_AMPL_WIDTH - 1),
		30140 => to_unsigned(8169, LUT_AMPL_WIDTH - 1),
		30141 => to_unsigned(8166, LUT_AMPL_WIDTH - 1),
		30142 => to_unsigned(8163, LUT_AMPL_WIDTH - 1),
		30143 => to_unsigned(8160, LUT_AMPL_WIDTH - 1),
		30144 => to_unsigned(8157, LUT_AMPL_WIDTH - 1),
		30145 => to_unsigned(8154, LUT_AMPL_WIDTH - 1),
		30146 => to_unsigned(8151, LUT_AMPL_WIDTH - 1),
		30147 => to_unsigned(8147, LUT_AMPL_WIDTH - 1),
		30148 => to_unsigned(8144, LUT_AMPL_WIDTH - 1),
		30149 => to_unsigned(8141, LUT_AMPL_WIDTH - 1),
		30150 => to_unsigned(8138, LUT_AMPL_WIDTH - 1),
		30151 => to_unsigned(8135, LUT_AMPL_WIDTH - 1),
		30152 => to_unsigned(8132, LUT_AMPL_WIDTH - 1),
		30153 => to_unsigned(8129, LUT_AMPL_WIDTH - 1),
		30154 => to_unsigned(8126, LUT_AMPL_WIDTH - 1),
		30155 => to_unsigned(8123, LUT_AMPL_WIDTH - 1),
		30156 => to_unsigned(8120, LUT_AMPL_WIDTH - 1),
		30157 => to_unsigned(8117, LUT_AMPL_WIDTH - 1),
		30158 => to_unsigned(8114, LUT_AMPL_WIDTH - 1),
		30159 => to_unsigned(8111, LUT_AMPL_WIDTH - 1),
		30160 => to_unsigned(8108, LUT_AMPL_WIDTH - 1),
		30161 => to_unsigned(8105, LUT_AMPL_WIDTH - 1),
		30162 => to_unsigned(8102, LUT_AMPL_WIDTH - 1),
		30163 => to_unsigned(8099, LUT_AMPL_WIDTH - 1),
		30164 => to_unsigned(8096, LUT_AMPL_WIDTH - 1),
		30165 => to_unsigned(8093, LUT_AMPL_WIDTH - 1),
		30166 => to_unsigned(8090, LUT_AMPL_WIDTH - 1),
		30167 => to_unsigned(8087, LUT_AMPL_WIDTH - 1),
		30168 => to_unsigned(8084, LUT_AMPL_WIDTH - 1),
		30169 => to_unsigned(8081, LUT_AMPL_WIDTH - 1),
		30170 => to_unsigned(8077, LUT_AMPL_WIDTH - 1),
		30171 => to_unsigned(8074, LUT_AMPL_WIDTH - 1),
		30172 => to_unsigned(8071, LUT_AMPL_WIDTH - 1),
		30173 => to_unsigned(8068, LUT_AMPL_WIDTH - 1),
		30174 => to_unsigned(8065, LUT_AMPL_WIDTH - 1),
		30175 => to_unsigned(8062, LUT_AMPL_WIDTH - 1),
		30176 => to_unsigned(8059, LUT_AMPL_WIDTH - 1),
		30177 => to_unsigned(8056, LUT_AMPL_WIDTH - 1),
		30178 => to_unsigned(8053, LUT_AMPL_WIDTH - 1),
		30179 => to_unsigned(8050, LUT_AMPL_WIDTH - 1),
		30180 => to_unsigned(8047, LUT_AMPL_WIDTH - 1),
		30181 => to_unsigned(8044, LUT_AMPL_WIDTH - 1),
		30182 => to_unsigned(8041, LUT_AMPL_WIDTH - 1),
		30183 => to_unsigned(8038, LUT_AMPL_WIDTH - 1),
		30184 => to_unsigned(8035, LUT_AMPL_WIDTH - 1),
		30185 => to_unsigned(8032, LUT_AMPL_WIDTH - 1),
		30186 => to_unsigned(8029, LUT_AMPL_WIDTH - 1),
		30187 => to_unsigned(8026, LUT_AMPL_WIDTH - 1),
		30188 => to_unsigned(8023, LUT_AMPL_WIDTH - 1),
		30189 => to_unsigned(8020, LUT_AMPL_WIDTH - 1),
		30190 => to_unsigned(8017, LUT_AMPL_WIDTH - 1),
		30191 => to_unsigned(8014, LUT_AMPL_WIDTH - 1),
		30192 => to_unsigned(8010, LUT_AMPL_WIDTH - 1),
		30193 => to_unsigned(8007, LUT_AMPL_WIDTH - 1),
		30194 => to_unsigned(8004, LUT_AMPL_WIDTH - 1),
		30195 => to_unsigned(8001, LUT_AMPL_WIDTH - 1),
		30196 => to_unsigned(7998, LUT_AMPL_WIDTH - 1),
		30197 => to_unsigned(7995, LUT_AMPL_WIDTH - 1),
		30198 => to_unsigned(7992, LUT_AMPL_WIDTH - 1),
		30199 => to_unsigned(7989, LUT_AMPL_WIDTH - 1),
		30200 => to_unsigned(7986, LUT_AMPL_WIDTH - 1),
		30201 => to_unsigned(7983, LUT_AMPL_WIDTH - 1),
		30202 => to_unsigned(7980, LUT_AMPL_WIDTH - 1),
		30203 => to_unsigned(7977, LUT_AMPL_WIDTH - 1),
		30204 => to_unsigned(7974, LUT_AMPL_WIDTH - 1),
		30205 => to_unsigned(7971, LUT_AMPL_WIDTH - 1),
		30206 => to_unsigned(7968, LUT_AMPL_WIDTH - 1),
		30207 => to_unsigned(7965, LUT_AMPL_WIDTH - 1),
		30208 => to_unsigned(7962, LUT_AMPL_WIDTH - 1),
		30209 => to_unsigned(7959, LUT_AMPL_WIDTH - 1),
		30210 => to_unsigned(7956, LUT_AMPL_WIDTH - 1),
		30211 => to_unsigned(7953, LUT_AMPL_WIDTH - 1),
		30212 => to_unsigned(7950, LUT_AMPL_WIDTH - 1),
		30213 => to_unsigned(7946, LUT_AMPL_WIDTH - 1),
		30214 => to_unsigned(7943, LUT_AMPL_WIDTH - 1),
		30215 => to_unsigned(7940, LUT_AMPL_WIDTH - 1),
		30216 => to_unsigned(7937, LUT_AMPL_WIDTH - 1),
		30217 => to_unsigned(7934, LUT_AMPL_WIDTH - 1),
		30218 => to_unsigned(7931, LUT_AMPL_WIDTH - 1),
		30219 => to_unsigned(7928, LUT_AMPL_WIDTH - 1),
		30220 => to_unsigned(7925, LUT_AMPL_WIDTH - 1),
		30221 => to_unsigned(7922, LUT_AMPL_WIDTH - 1),
		30222 => to_unsigned(7919, LUT_AMPL_WIDTH - 1),
		30223 => to_unsigned(7916, LUT_AMPL_WIDTH - 1),
		30224 => to_unsigned(7913, LUT_AMPL_WIDTH - 1),
		30225 => to_unsigned(7910, LUT_AMPL_WIDTH - 1),
		30226 => to_unsigned(7907, LUT_AMPL_WIDTH - 1),
		30227 => to_unsigned(7904, LUT_AMPL_WIDTH - 1),
		30228 => to_unsigned(7901, LUT_AMPL_WIDTH - 1),
		30229 => to_unsigned(7898, LUT_AMPL_WIDTH - 1),
		30230 => to_unsigned(7895, LUT_AMPL_WIDTH - 1),
		30231 => to_unsigned(7892, LUT_AMPL_WIDTH - 1),
		30232 => to_unsigned(7889, LUT_AMPL_WIDTH - 1),
		30233 => to_unsigned(7886, LUT_AMPL_WIDTH - 1),
		30234 => to_unsigned(7882, LUT_AMPL_WIDTH - 1),
		30235 => to_unsigned(7879, LUT_AMPL_WIDTH - 1),
		30236 => to_unsigned(7876, LUT_AMPL_WIDTH - 1),
		30237 => to_unsigned(7873, LUT_AMPL_WIDTH - 1),
		30238 => to_unsigned(7870, LUT_AMPL_WIDTH - 1),
		30239 => to_unsigned(7867, LUT_AMPL_WIDTH - 1),
		30240 => to_unsigned(7864, LUT_AMPL_WIDTH - 1),
		30241 => to_unsigned(7861, LUT_AMPL_WIDTH - 1),
		30242 => to_unsigned(7858, LUT_AMPL_WIDTH - 1),
		30243 => to_unsigned(7855, LUT_AMPL_WIDTH - 1),
		30244 => to_unsigned(7852, LUT_AMPL_WIDTH - 1),
		30245 => to_unsigned(7849, LUT_AMPL_WIDTH - 1),
		30246 => to_unsigned(7846, LUT_AMPL_WIDTH - 1),
		30247 => to_unsigned(7843, LUT_AMPL_WIDTH - 1),
		30248 => to_unsigned(7840, LUT_AMPL_WIDTH - 1),
		30249 => to_unsigned(7837, LUT_AMPL_WIDTH - 1),
		30250 => to_unsigned(7834, LUT_AMPL_WIDTH - 1),
		30251 => to_unsigned(7831, LUT_AMPL_WIDTH - 1),
		30252 => to_unsigned(7828, LUT_AMPL_WIDTH - 1),
		30253 => to_unsigned(7825, LUT_AMPL_WIDTH - 1),
		30254 => to_unsigned(7821, LUT_AMPL_WIDTH - 1),
		30255 => to_unsigned(7818, LUT_AMPL_WIDTH - 1),
		30256 => to_unsigned(7815, LUT_AMPL_WIDTH - 1),
		30257 => to_unsigned(7812, LUT_AMPL_WIDTH - 1),
		30258 => to_unsigned(7809, LUT_AMPL_WIDTH - 1),
		30259 => to_unsigned(7806, LUT_AMPL_WIDTH - 1),
		30260 => to_unsigned(7803, LUT_AMPL_WIDTH - 1),
		30261 => to_unsigned(7800, LUT_AMPL_WIDTH - 1),
		30262 => to_unsigned(7797, LUT_AMPL_WIDTH - 1),
		30263 => to_unsigned(7794, LUT_AMPL_WIDTH - 1),
		30264 => to_unsigned(7791, LUT_AMPL_WIDTH - 1),
		30265 => to_unsigned(7788, LUT_AMPL_WIDTH - 1),
		30266 => to_unsigned(7785, LUT_AMPL_WIDTH - 1),
		30267 => to_unsigned(7782, LUT_AMPL_WIDTH - 1),
		30268 => to_unsigned(7779, LUT_AMPL_WIDTH - 1),
		30269 => to_unsigned(7776, LUT_AMPL_WIDTH - 1),
		30270 => to_unsigned(7773, LUT_AMPL_WIDTH - 1),
		30271 => to_unsigned(7770, LUT_AMPL_WIDTH - 1),
		30272 => to_unsigned(7767, LUT_AMPL_WIDTH - 1),
		30273 => to_unsigned(7764, LUT_AMPL_WIDTH - 1),
		30274 => to_unsigned(7760, LUT_AMPL_WIDTH - 1),
		30275 => to_unsigned(7757, LUT_AMPL_WIDTH - 1),
		30276 => to_unsigned(7754, LUT_AMPL_WIDTH - 1),
		30277 => to_unsigned(7751, LUT_AMPL_WIDTH - 1),
		30278 => to_unsigned(7748, LUT_AMPL_WIDTH - 1),
		30279 => to_unsigned(7745, LUT_AMPL_WIDTH - 1),
		30280 => to_unsigned(7742, LUT_AMPL_WIDTH - 1),
		30281 => to_unsigned(7739, LUT_AMPL_WIDTH - 1),
		30282 => to_unsigned(7736, LUT_AMPL_WIDTH - 1),
		30283 => to_unsigned(7733, LUT_AMPL_WIDTH - 1),
		30284 => to_unsigned(7730, LUT_AMPL_WIDTH - 1),
		30285 => to_unsigned(7727, LUT_AMPL_WIDTH - 1),
		30286 => to_unsigned(7724, LUT_AMPL_WIDTH - 1),
		30287 => to_unsigned(7721, LUT_AMPL_WIDTH - 1),
		30288 => to_unsigned(7718, LUT_AMPL_WIDTH - 1),
		30289 => to_unsigned(7715, LUT_AMPL_WIDTH - 1),
		30290 => to_unsigned(7712, LUT_AMPL_WIDTH - 1),
		30291 => to_unsigned(7709, LUT_AMPL_WIDTH - 1),
		30292 => to_unsigned(7705, LUT_AMPL_WIDTH - 1),
		30293 => to_unsigned(7702, LUT_AMPL_WIDTH - 1),
		30294 => to_unsigned(7699, LUT_AMPL_WIDTH - 1),
		30295 => to_unsigned(7696, LUT_AMPL_WIDTH - 1),
		30296 => to_unsigned(7693, LUT_AMPL_WIDTH - 1),
		30297 => to_unsigned(7690, LUT_AMPL_WIDTH - 1),
		30298 => to_unsigned(7687, LUT_AMPL_WIDTH - 1),
		30299 => to_unsigned(7684, LUT_AMPL_WIDTH - 1),
		30300 => to_unsigned(7681, LUT_AMPL_WIDTH - 1),
		30301 => to_unsigned(7678, LUT_AMPL_WIDTH - 1),
		30302 => to_unsigned(7675, LUT_AMPL_WIDTH - 1),
		30303 => to_unsigned(7672, LUT_AMPL_WIDTH - 1),
		30304 => to_unsigned(7669, LUT_AMPL_WIDTH - 1),
		30305 => to_unsigned(7666, LUT_AMPL_WIDTH - 1),
		30306 => to_unsigned(7663, LUT_AMPL_WIDTH - 1),
		30307 => to_unsigned(7660, LUT_AMPL_WIDTH - 1),
		30308 => to_unsigned(7657, LUT_AMPL_WIDTH - 1),
		30309 => to_unsigned(7654, LUT_AMPL_WIDTH - 1),
		30310 => to_unsigned(7651, LUT_AMPL_WIDTH - 1),
		30311 => to_unsigned(7647, LUT_AMPL_WIDTH - 1),
		30312 => to_unsigned(7644, LUT_AMPL_WIDTH - 1),
		30313 => to_unsigned(7641, LUT_AMPL_WIDTH - 1),
		30314 => to_unsigned(7638, LUT_AMPL_WIDTH - 1),
		30315 => to_unsigned(7635, LUT_AMPL_WIDTH - 1),
		30316 => to_unsigned(7632, LUT_AMPL_WIDTH - 1),
		30317 => to_unsigned(7629, LUT_AMPL_WIDTH - 1),
		30318 => to_unsigned(7626, LUT_AMPL_WIDTH - 1),
		30319 => to_unsigned(7623, LUT_AMPL_WIDTH - 1),
		30320 => to_unsigned(7620, LUT_AMPL_WIDTH - 1),
		30321 => to_unsigned(7617, LUT_AMPL_WIDTH - 1),
		30322 => to_unsigned(7614, LUT_AMPL_WIDTH - 1),
		30323 => to_unsigned(7611, LUT_AMPL_WIDTH - 1),
		30324 => to_unsigned(7608, LUT_AMPL_WIDTH - 1),
		30325 => to_unsigned(7605, LUT_AMPL_WIDTH - 1),
		30326 => to_unsigned(7602, LUT_AMPL_WIDTH - 1),
		30327 => to_unsigned(7599, LUT_AMPL_WIDTH - 1),
		30328 => to_unsigned(7596, LUT_AMPL_WIDTH - 1),
		30329 => to_unsigned(7592, LUT_AMPL_WIDTH - 1),
		30330 => to_unsigned(7589, LUT_AMPL_WIDTH - 1),
		30331 => to_unsigned(7586, LUT_AMPL_WIDTH - 1),
		30332 => to_unsigned(7583, LUT_AMPL_WIDTH - 1),
		30333 => to_unsigned(7580, LUT_AMPL_WIDTH - 1),
		30334 => to_unsigned(7577, LUT_AMPL_WIDTH - 1),
		30335 => to_unsigned(7574, LUT_AMPL_WIDTH - 1),
		30336 => to_unsigned(7571, LUT_AMPL_WIDTH - 1),
		30337 => to_unsigned(7568, LUT_AMPL_WIDTH - 1),
		30338 => to_unsigned(7565, LUT_AMPL_WIDTH - 1),
		30339 => to_unsigned(7562, LUT_AMPL_WIDTH - 1),
		30340 => to_unsigned(7559, LUT_AMPL_WIDTH - 1),
		30341 => to_unsigned(7556, LUT_AMPL_WIDTH - 1),
		30342 => to_unsigned(7553, LUT_AMPL_WIDTH - 1),
		30343 => to_unsigned(7550, LUT_AMPL_WIDTH - 1),
		30344 => to_unsigned(7547, LUT_AMPL_WIDTH - 1),
		30345 => to_unsigned(7544, LUT_AMPL_WIDTH - 1),
		30346 => to_unsigned(7541, LUT_AMPL_WIDTH - 1),
		30347 => to_unsigned(7537, LUT_AMPL_WIDTH - 1),
		30348 => to_unsigned(7534, LUT_AMPL_WIDTH - 1),
		30349 => to_unsigned(7531, LUT_AMPL_WIDTH - 1),
		30350 => to_unsigned(7528, LUT_AMPL_WIDTH - 1),
		30351 => to_unsigned(7525, LUT_AMPL_WIDTH - 1),
		30352 => to_unsigned(7522, LUT_AMPL_WIDTH - 1),
		30353 => to_unsigned(7519, LUT_AMPL_WIDTH - 1),
		30354 => to_unsigned(7516, LUT_AMPL_WIDTH - 1),
		30355 => to_unsigned(7513, LUT_AMPL_WIDTH - 1),
		30356 => to_unsigned(7510, LUT_AMPL_WIDTH - 1),
		30357 => to_unsigned(7507, LUT_AMPL_WIDTH - 1),
		30358 => to_unsigned(7504, LUT_AMPL_WIDTH - 1),
		30359 => to_unsigned(7501, LUT_AMPL_WIDTH - 1),
		30360 => to_unsigned(7498, LUT_AMPL_WIDTH - 1),
		30361 => to_unsigned(7495, LUT_AMPL_WIDTH - 1),
		30362 => to_unsigned(7492, LUT_AMPL_WIDTH - 1),
		30363 => to_unsigned(7489, LUT_AMPL_WIDTH - 1),
		30364 => to_unsigned(7485, LUT_AMPL_WIDTH - 1),
		30365 => to_unsigned(7482, LUT_AMPL_WIDTH - 1),
		30366 => to_unsigned(7479, LUT_AMPL_WIDTH - 1),
		30367 => to_unsigned(7476, LUT_AMPL_WIDTH - 1),
		30368 => to_unsigned(7473, LUT_AMPL_WIDTH - 1),
		30369 => to_unsigned(7470, LUT_AMPL_WIDTH - 1),
		30370 => to_unsigned(7467, LUT_AMPL_WIDTH - 1),
		30371 => to_unsigned(7464, LUT_AMPL_WIDTH - 1),
		30372 => to_unsigned(7461, LUT_AMPL_WIDTH - 1),
		30373 => to_unsigned(7458, LUT_AMPL_WIDTH - 1),
		30374 => to_unsigned(7455, LUT_AMPL_WIDTH - 1),
		30375 => to_unsigned(7452, LUT_AMPL_WIDTH - 1),
		30376 => to_unsigned(7449, LUT_AMPL_WIDTH - 1),
		30377 => to_unsigned(7446, LUT_AMPL_WIDTH - 1),
		30378 => to_unsigned(7443, LUT_AMPL_WIDTH - 1),
		30379 => to_unsigned(7440, LUT_AMPL_WIDTH - 1),
		30380 => to_unsigned(7437, LUT_AMPL_WIDTH - 1),
		30381 => to_unsigned(7433, LUT_AMPL_WIDTH - 1),
		30382 => to_unsigned(7430, LUT_AMPL_WIDTH - 1),
		30383 => to_unsigned(7427, LUT_AMPL_WIDTH - 1),
		30384 => to_unsigned(7424, LUT_AMPL_WIDTH - 1),
		30385 => to_unsigned(7421, LUT_AMPL_WIDTH - 1),
		30386 => to_unsigned(7418, LUT_AMPL_WIDTH - 1),
		30387 => to_unsigned(7415, LUT_AMPL_WIDTH - 1),
		30388 => to_unsigned(7412, LUT_AMPL_WIDTH - 1),
		30389 => to_unsigned(7409, LUT_AMPL_WIDTH - 1),
		30390 => to_unsigned(7406, LUT_AMPL_WIDTH - 1),
		30391 => to_unsigned(7403, LUT_AMPL_WIDTH - 1),
		30392 => to_unsigned(7400, LUT_AMPL_WIDTH - 1),
		30393 => to_unsigned(7397, LUT_AMPL_WIDTH - 1),
		30394 => to_unsigned(7394, LUT_AMPL_WIDTH - 1),
		30395 => to_unsigned(7391, LUT_AMPL_WIDTH - 1),
		30396 => to_unsigned(7388, LUT_AMPL_WIDTH - 1),
		30397 => to_unsigned(7385, LUT_AMPL_WIDTH - 1),
		30398 => to_unsigned(7381, LUT_AMPL_WIDTH - 1),
		30399 => to_unsigned(7378, LUT_AMPL_WIDTH - 1),
		30400 => to_unsigned(7375, LUT_AMPL_WIDTH - 1),
		30401 => to_unsigned(7372, LUT_AMPL_WIDTH - 1),
		30402 => to_unsigned(7369, LUT_AMPL_WIDTH - 1),
		30403 => to_unsigned(7366, LUT_AMPL_WIDTH - 1),
		30404 => to_unsigned(7363, LUT_AMPL_WIDTH - 1),
		30405 => to_unsigned(7360, LUT_AMPL_WIDTH - 1),
		30406 => to_unsigned(7357, LUT_AMPL_WIDTH - 1),
		30407 => to_unsigned(7354, LUT_AMPL_WIDTH - 1),
		30408 => to_unsigned(7351, LUT_AMPL_WIDTH - 1),
		30409 => to_unsigned(7348, LUT_AMPL_WIDTH - 1),
		30410 => to_unsigned(7345, LUT_AMPL_WIDTH - 1),
		30411 => to_unsigned(7342, LUT_AMPL_WIDTH - 1),
		30412 => to_unsigned(7339, LUT_AMPL_WIDTH - 1),
		30413 => to_unsigned(7336, LUT_AMPL_WIDTH - 1),
		30414 => to_unsigned(7332, LUT_AMPL_WIDTH - 1),
		30415 => to_unsigned(7329, LUT_AMPL_WIDTH - 1),
		30416 => to_unsigned(7326, LUT_AMPL_WIDTH - 1),
		30417 => to_unsigned(7323, LUT_AMPL_WIDTH - 1),
		30418 => to_unsigned(7320, LUT_AMPL_WIDTH - 1),
		30419 => to_unsigned(7317, LUT_AMPL_WIDTH - 1),
		30420 => to_unsigned(7314, LUT_AMPL_WIDTH - 1),
		30421 => to_unsigned(7311, LUT_AMPL_WIDTH - 1),
		30422 => to_unsigned(7308, LUT_AMPL_WIDTH - 1),
		30423 => to_unsigned(7305, LUT_AMPL_WIDTH - 1),
		30424 => to_unsigned(7302, LUT_AMPL_WIDTH - 1),
		30425 => to_unsigned(7299, LUT_AMPL_WIDTH - 1),
		30426 => to_unsigned(7296, LUT_AMPL_WIDTH - 1),
		30427 => to_unsigned(7293, LUT_AMPL_WIDTH - 1),
		30428 => to_unsigned(7290, LUT_AMPL_WIDTH - 1),
		30429 => to_unsigned(7287, LUT_AMPL_WIDTH - 1),
		30430 => to_unsigned(7283, LUT_AMPL_WIDTH - 1),
		30431 => to_unsigned(7280, LUT_AMPL_WIDTH - 1),
		30432 => to_unsigned(7277, LUT_AMPL_WIDTH - 1),
		30433 => to_unsigned(7274, LUT_AMPL_WIDTH - 1),
		30434 => to_unsigned(7271, LUT_AMPL_WIDTH - 1),
		30435 => to_unsigned(7268, LUT_AMPL_WIDTH - 1),
		30436 => to_unsigned(7265, LUT_AMPL_WIDTH - 1),
		30437 => to_unsigned(7262, LUT_AMPL_WIDTH - 1),
		30438 => to_unsigned(7259, LUT_AMPL_WIDTH - 1),
		30439 => to_unsigned(7256, LUT_AMPL_WIDTH - 1),
		30440 => to_unsigned(7253, LUT_AMPL_WIDTH - 1),
		30441 => to_unsigned(7250, LUT_AMPL_WIDTH - 1),
		30442 => to_unsigned(7247, LUT_AMPL_WIDTH - 1),
		30443 => to_unsigned(7244, LUT_AMPL_WIDTH - 1),
		30444 => to_unsigned(7241, LUT_AMPL_WIDTH - 1),
		30445 => to_unsigned(7238, LUT_AMPL_WIDTH - 1),
		30446 => to_unsigned(7234, LUT_AMPL_WIDTH - 1),
		30447 => to_unsigned(7231, LUT_AMPL_WIDTH - 1),
		30448 => to_unsigned(7228, LUT_AMPL_WIDTH - 1),
		30449 => to_unsigned(7225, LUT_AMPL_WIDTH - 1),
		30450 => to_unsigned(7222, LUT_AMPL_WIDTH - 1),
		30451 => to_unsigned(7219, LUT_AMPL_WIDTH - 1),
		30452 => to_unsigned(7216, LUT_AMPL_WIDTH - 1),
		30453 => to_unsigned(7213, LUT_AMPL_WIDTH - 1),
		30454 => to_unsigned(7210, LUT_AMPL_WIDTH - 1),
		30455 => to_unsigned(7207, LUT_AMPL_WIDTH - 1),
		30456 => to_unsigned(7204, LUT_AMPL_WIDTH - 1),
		30457 => to_unsigned(7201, LUT_AMPL_WIDTH - 1),
		30458 => to_unsigned(7198, LUT_AMPL_WIDTH - 1),
		30459 => to_unsigned(7195, LUT_AMPL_WIDTH - 1),
		30460 => to_unsigned(7192, LUT_AMPL_WIDTH - 1),
		30461 => to_unsigned(7188, LUT_AMPL_WIDTH - 1),
		30462 => to_unsigned(7185, LUT_AMPL_WIDTH - 1),
		30463 => to_unsigned(7182, LUT_AMPL_WIDTH - 1),
		30464 => to_unsigned(7179, LUT_AMPL_WIDTH - 1),
		30465 => to_unsigned(7176, LUT_AMPL_WIDTH - 1),
		30466 => to_unsigned(7173, LUT_AMPL_WIDTH - 1),
		30467 => to_unsigned(7170, LUT_AMPL_WIDTH - 1),
		30468 => to_unsigned(7167, LUT_AMPL_WIDTH - 1),
		30469 => to_unsigned(7164, LUT_AMPL_WIDTH - 1),
		30470 => to_unsigned(7161, LUT_AMPL_WIDTH - 1),
		30471 => to_unsigned(7158, LUT_AMPL_WIDTH - 1),
		30472 => to_unsigned(7155, LUT_AMPL_WIDTH - 1),
		30473 => to_unsigned(7152, LUT_AMPL_WIDTH - 1),
		30474 => to_unsigned(7149, LUT_AMPL_WIDTH - 1),
		30475 => to_unsigned(7146, LUT_AMPL_WIDTH - 1),
		30476 => to_unsigned(7143, LUT_AMPL_WIDTH - 1),
		30477 => to_unsigned(7139, LUT_AMPL_WIDTH - 1),
		30478 => to_unsigned(7136, LUT_AMPL_WIDTH - 1),
		30479 => to_unsigned(7133, LUT_AMPL_WIDTH - 1),
		30480 => to_unsigned(7130, LUT_AMPL_WIDTH - 1),
		30481 => to_unsigned(7127, LUT_AMPL_WIDTH - 1),
		30482 => to_unsigned(7124, LUT_AMPL_WIDTH - 1),
		30483 => to_unsigned(7121, LUT_AMPL_WIDTH - 1),
		30484 => to_unsigned(7118, LUT_AMPL_WIDTH - 1),
		30485 => to_unsigned(7115, LUT_AMPL_WIDTH - 1),
		30486 => to_unsigned(7112, LUT_AMPL_WIDTH - 1),
		30487 => to_unsigned(7109, LUT_AMPL_WIDTH - 1),
		30488 => to_unsigned(7106, LUT_AMPL_WIDTH - 1),
		30489 => to_unsigned(7103, LUT_AMPL_WIDTH - 1),
		30490 => to_unsigned(7100, LUT_AMPL_WIDTH - 1),
		30491 => to_unsigned(7097, LUT_AMPL_WIDTH - 1),
		30492 => to_unsigned(7093, LUT_AMPL_WIDTH - 1),
		30493 => to_unsigned(7090, LUT_AMPL_WIDTH - 1),
		30494 => to_unsigned(7087, LUT_AMPL_WIDTH - 1),
		30495 => to_unsigned(7084, LUT_AMPL_WIDTH - 1),
		30496 => to_unsigned(7081, LUT_AMPL_WIDTH - 1),
		30497 => to_unsigned(7078, LUT_AMPL_WIDTH - 1),
		30498 => to_unsigned(7075, LUT_AMPL_WIDTH - 1),
		30499 => to_unsigned(7072, LUT_AMPL_WIDTH - 1),
		30500 => to_unsigned(7069, LUT_AMPL_WIDTH - 1),
		30501 => to_unsigned(7066, LUT_AMPL_WIDTH - 1),
		30502 => to_unsigned(7063, LUT_AMPL_WIDTH - 1),
		30503 => to_unsigned(7060, LUT_AMPL_WIDTH - 1),
		30504 => to_unsigned(7057, LUT_AMPL_WIDTH - 1),
		30505 => to_unsigned(7054, LUT_AMPL_WIDTH - 1),
		30506 => to_unsigned(7050, LUT_AMPL_WIDTH - 1),
		30507 => to_unsigned(7047, LUT_AMPL_WIDTH - 1),
		30508 => to_unsigned(7044, LUT_AMPL_WIDTH - 1),
		30509 => to_unsigned(7041, LUT_AMPL_WIDTH - 1),
		30510 => to_unsigned(7038, LUT_AMPL_WIDTH - 1),
		30511 => to_unsigned(7035, LUT_AMPL_WIDTH - 1),
		30512 => to_unsigned(7032, LUT_AMPL_WIDTH - 1),
		30513 => to_unsigned(7029, LUT_AMPL_WIDTH - 1),
		30514 => to_unsigned(7026, LUT_AMPL_WIDTH - 1),
		30515 => to_unsigned(7023, LUT_AMPL_WIDTH - 1),
		30516 => to_unsigned(7020, LUT_AMPL_WIDTH - 1),
		30517 => to_unsigned(7017, LUT_AMPL_WIDTH - 1),
		30518 => to_unsigned(7014, LUT_AMPL_WIDTH - 1),
		30519 => to_unsigned(7011, LUT_AMPL_WIDTH - 1),
		30520 => to_unsigned(7008, LUT_AMPL_WIDTH - 1),
		30521 => to_unsigned(7004, LUT_AMPL_WIDTH - 1),
		30522 => to_unsigned(7001, LUT_AMPL_WIDTH - 1),
		30523 => to_unsigned(6998, LUT_AMPL_WIDTH - 1),
		30524 => to_unsigned(6995, LUT_AMPL_WIDTH - 1),
		30525 => to_unsigned(6992, LUT_AMPL_WIDTH - 1),
		30526 => to_unsigned(6989, LUT_AMPL_WIDTH - 1),
		30527 => to_unsigned(6986, LUT_AMPL_WIDTH - 1),
		30528 => to_unsigned(6983, LUT_AMPL_WIDTH - 1),
		30529 => to_unsigned(6980, LUT_AMPL_WIDTH - 1),
		30530 => to_unsigned(6977, LUT_AMPL_WIDTH - 1),
		30531 => to_unsigned(6974, LUT_AMPL_WIDTH - 1),
		30532 => to_unsigned(6971, LUT_AMPL_WIDTH - 1),
		30533 => to_unsigned(6968, LUT_AMPL_WIDTH - 1),
		30534 => to_unsigned(6965, LUT_AMPL_WIDTH - 1),
		30535 => to_unsigned(6961, LUT_AMPL_WIDTH - 1),
		30536 => to_unsigned(6958, LUT_AMPL_WIDTH - 1),
		30537 => to_unsigned(6955, LUT_AMPL_WIDTH - 1),
		30538 => to_unsigned(6952, LUT_AMPL_WIDTH - 1),
		30539 => to_unsigned(6949, LUT_AMPL_WIDTH - 1),
		30540 => to_unsigned(6946, LUT_AMPL_WIDTH - 1),
		30541 => to_unsigned(6943, LUT_AMPL_WIDTH - 1),
		30542 => to_unsigned(6940, LUT_AMPL_WIDTH - 1),
		30543 => to_unsigned(6937, LUT_AMPL_WIDTH - 1),
		30544 => to_unsigned(6934, LUT_AMPL_WIDTH - 1),
		30545 => to_unsigned(6931, LUT_AMPL_WIDTH - 1),
		30546 => to_unsigned(6928, LUT_AMPL_WIDTH - 1),
		30547 => to_unsigned(6925, LUT_AMPL_WIDTH - 1),
		30548 => to_unsigned(6922, LUT_AMPL_WIDTH - 1),
		30549 => to_unsigned(6919, LUT_AMPL_WIDTH - 1),
		30550 => to_unsigned(6915, LUT_AMPL_WIDTH - 1),
		30551 => to_unsigned(6912, LUT_AMPL_WIDTH - 1),
		30552 => to_unsigned(6909, LUT_AMPL_WIDTH - 1),
		30553 => to_unsigned(6906, LUT_AMPL_WIDTH - 1),
		30554 => to_unsigned(6903, LUT_AMPL_WIDTH - 1),
		30555 => to_unsigned(6900, LUT_AMPL_WIDTH - 1),
		30556 => to_unsigned(6897, LUT_AMPL_WIDTH - 1),
		30557 => to_unsigned(6894, LUT_AMPL_WIDTH - 1),
		30558 => to_unsigned(6891, LUT_AMPL_WIDTH - 1),
		30559 => to_unsigned(6888, LUT_AMPL_WIDTH - 1),
		30560 => to_unsigned(6885, LUT_AMPL_WIDTH - 1),
		30561 => to_unsigned(6882, LUT_AMPL_WIDTH - 1),
		30562 => to_unsigned(6879, LUT_AMPL_WIDTH - 1),
		30563 => to_unsigned(6876, LUT_AMPL_WIDTH - 1),
		30564 => to_unsigned(6872, LUT_AMPL_WIDTH - 1),
		30565 => to_unsigned(6869, LUT_AMPL_WIDTH - 1),
		30566 => to_unsigned(6866, LUT_AMPL_WIDTH - 1),
		30567 => to_unsigned(6863, LUT_AMPL_WIDTH - 1),
		30568 => to_unsigned(6860, LUT_AMPL_WIDTH - 1),
		30569 => to_unsigned(6857, LUT_AMPL_WIDTH - 1),
		30570 => to_unsigned(6854, LUT_AMPL_WIDTH - 1),
		30571 => to_unsigned(6851, LUT_AMPL_WIDTH - 1),
		30572 => to_unsigned(6848, LUT_AMPL_WIDTH - 1),
		30573 => to_unsigned(6845, LUT_AMPL_WIDTH - 1),
		30574 => to_unsigned(6842, LUT_AMPL_WIDTH - 1),
		30575 => to_unsigned(6839, LUT_AMPL_WIDTH - 1),
		30576 => to_unsigned(6836, LUT_AMPL_WIDTH - 1),
		30577 => to_unsigned(6833, LUT_AMPL_WIDTH - 1),
		30578 => to_unsigned(6829, LUT_AMPL_WIDTH - 1),
		30579 => to_unsigned(6826, LUT_AMPL_WIDTH - 1),
		30580 => to_unsigned(6823, LUT_AMPL_WIDTH - 1),
		30581 => to_unsigned(6820, LUT_AMPL_WIDTH - 1),
		30582 => to_unsigned(6817, LUT_AMPL_WIDTH - 1),
		30583 => to_unsigned(6814, LUT_AMPL_WIDTH - 1),
		30584 => to_unsigned(6811, LUT_AMPL_WIDTH - 1),
		30585 => to_unsigned(6808, LUT_AMPL_WIDTH - 1),
		30586 => to_unsigned(6805, LUT_AMPL_WIDTH - 1),
		30587 => to_unsigned(6802, LUT_AMPL_WIDTH - 1),
		30588 => to_unsigned(6799, LUT_AMPL_WIDTH - 1),
		30589 => to_unsigned(6796, LUT_AMPL_WIDTH - 1),
		30590 => to_unsigned(6793, LUT_AMPL_WIDTH - 1),
		30591 => to_unsigned(6789, LUT_AMPL_WIDTH - 1),
		30592 => to_unsigned(6786, LUT_AMPL_WIDTH - 1),
		30593 => to_unsigned(6783, LUT_AMPL_WIDTH - 1),
		30594 => to_unsigned(6780, LUT_AMPL_WIDTH - 1),
		30595 => to_unsigned(6777, LUT_AMPL_WIDTH - 1),
		30596 => to_unsigned(6774, LUT_AMPL_WIDTH - 1),
		30597 => to_unsigned(6771, LUT_AMPL_WIDTH - 1),
		30598 => to_unsigned(6768, LUT_AMPL_WIDTH - 1),
		30599 => to_unsigned(6765, LUT_AMPL_WIDTH - 1),
		30600 => to_unsigned(6762, LUT_AMPL_WIDTH - 1),
		30601 => to_unsigned(6759, LUT_AMPL_WIDTH - 1),
		30602 => to_unsigned(6756, LUT_AMPL_WIDTH - 1),
		30603 => to_unsigned(6753, LUT_AMPL_WIDTH - 1),
		30604 => to_unsigned(6750, LUT_AMPL_WIDTH - 1),
		30605 => to_unsigned(6746, LUT_AMPL_WIDTH - 1),
		30606 => to_unsigned(6743, LUT_AMPL_WIDTH - 1),
		30607 => to_unsigned(6740, LUT_AMPL_WIDTH - 1),
		30608 => to_unsigned(6737, LUT_AMPL_WIDTH - 1),
		30609 => to_unsigned(6734, LUT_AMPL_WIDTH - 1),
		30610 => to_unsigned(6731, LUT_AMPL_WIDTH - 1),
		30611 => to_unsigned(6728, LUT_AMPL_WIDTH - 1),
		30612 => to_unsigned(6725, LUT_AMPL_WIDTH - 1),
		30613 => to_unsigned(6722, LUT_AMPL_WIDTH - 1),
		30614 => to_unsigned(6719, LUT_AMPL_WIDTH - 1),
		30615 => to_unsigned(6716, LUT_AMPL_WIDTH - 1),
		30616 => to_unsigned(6713, LUT_AMPL_WIDTH - 1),
		30617 => to_unsigned(6710, LUT_AMPL_WIDTH - 1),
		30618 => to_unsigned(6706, LUT_AMPL_WIDTH - 1),
		30619 => to_unsigned(6703, LUT_AMPL_WIDTH - 1),
		30620 => to_unsigned(6700, LUT_AMPL_WIDTH - 1),
		30621 => to_unsigned(6697, LUT_AMPL_WIDTH - 1),
		30622 => to_unsigned(6694, LUT_AMPL_WIDTH - 1),
		30623 => to_unsigned(6691, LUT_AMPL_WIDTH - 1),
		30624 => to_unsigned(6688, LUT_AMPL_WIDTH - 1),
		30625 => to_unsigned(6685, LUT_AMPL_WIDTH - 1),
		30626 => to_unsigned(6682, LUT_AMPL_WIDTH - 1),
		30627 => to_unsigned(6679, LUT_AMPL_WIDTH - 1),
		30628 => to_unsigned(6676, LUT_AMPL_WIDTH - 1),
		30629 => to_unsigned(6673, LUT_AMPL_WIDTH - 1),
		30630 => to_unsigned(6670, LUT_AMPL_WIDTH - 1),
		30631 => to_unsigned(6667, LUT_AMPL_WIDTH - 1),
		30632 => to_unsigned(6663, LUT_AMPL_WIDTH - 1),
		30633 => to_unsigned(6660, LUT_AMPL_WIDTH - 1),
		30634 => to_unsigned(6657, LUT_AMPL_WIDTH - 1),
		30635 => to_unsigned(6654, LUT_AMPL_WIDTH - 1),
		30636 => to_unsigned(6651, LUT_AMPL_WIDTH - 1),
		30637 => to_unsigned(6648, LUT_AMPL_WIDTH - 1),
		30638 => to_unsigned(6645, LUT_AMPL_WIDTH - 1),
		30639 => to_unsigned(6642, LUT_AMPL_WIDTH - 1),
		30640 => to_unsigned(6639, LUT_AMPL_WIDTH - 1),
		30641 => to_unsigned(6636, LUT_AMPL_WIDTH - 1),
		30642 => to_unsigned(6633, LUT_AMPL_WIDTH - 1),
		30643 => to_unsigned(6630, LUT_AMPL_WIDTH - 1),
		30644 => to_unsigned(6627, LUT_AMPL_WIDTH - 1),
		30645 => to_unsigned(6623, LUT_AMPL_WIDTH - 1),
		30646 => to_unsigned(6620, LUT_AMPL_WIDTH - 1),
		30647 => to_unsigned(6617, LUT_AMPL_WIDTH - 1),
		30648 => to_unsigned(6614, LUT_AMPL_WIDTH - 1),
		30649 => to_unsigned(6611, LUT_AMPL_WIDTH - 1),
		30650 => to_unsigned(6608, LUT_AMPL_WIDTH - 1),
		30651 => to_unsigned(6605, LUT_AMPL_WIDTH - 1),
		30652 => to_unsigned(6602, LUT_AMPL_WIDTH - 1),
		30653 => to_unsigned(6599, LUT_AMPL_WIDTH - 1),
		30654 => to_unsigned(6596, LUT_AMPL_WIDTH - 1),
		30655 => to_unsigned(6593, LUT_AMPL_WIDTH - 1),
		30656 => to_unsigned(6590, LUT_AMPL_WIDTH - 1),
		30657 => to_unsigned(6587, LUT_AMPL_WIDTH - 1),
		30658 => to_unsigned(6583, LUT_AMPL_WIDTH - 1),
		30659 => to_unsigned(6580, LUT_AMPL_WIDTH - 1),
		30660 => to_unsigned(6577, LUT_AMPL_WIDTH - 1),
		30661 => to_unsigned(6574, LUT_AMPL_WIDTH - 1),
		30662 => to_unsigned(6571, LUT_AMPL_WIDTH - 1),
		30663 => to_unsigned(6568, LUT_AMPL_WIDTH - 1),
		30664 => to_unsigned(6565, LUT_AMPL_WIDTH - 1),
		30665 => to_unsigned(6562, LUT_AMPL_WIDTH - 1),
		30666 => to_unsigned(6559, LUT_AMPL_WIDTH - 1),
		30667 => to_unsigned(6556, LUT_AMPL_WIDTH - 1),
		30668 => to_unsigned(6553, LUT_AMPL_WIDTH - 1),
		30669 => to_unsigned(6550, LUT_AMPL_WIDTH - 1),
		30670 => to_unsigned(6547, LUT_AMPL_WIDTH - 1),
		30671 => to_unsigned(6543, LUT_AMPL_WIDTH - 1),
		30672 => to_unsigned(6540, LUT_AMPL_WIDTH - 1),
		30673 => to_unsigned(6537, LUT_AMPL_WIDTH - 1),
		30674 => to_unsigned(6534, LUT_AMPL_WIDTH - 1),
		30675 => to_unsigned(6531, LUT_AMPL_WIDTH - 1),
		30676 => to_unsigned(6528, LUT_AMPL_WIDTH - 1),
		30677 => to_unsigned(6525, LUT_AMPL_WIDTH - 1),
		30678 => to_unsigned(6522, LUT_AMPL_WIDTH - 1),
		30679 => to_unsigned(6519, LUT_AMPL_WIDTH - 1),
		30680 => to_unsigned(6516, LUT_AMPL_WIDTH - 1),
		30681 => to_unsigned(6513, LUT_AMPL_WIDTH - 1),
		30682 => to_unsigned(6510, LUT_AMPL_WIDTH - 1),
		30683 => to_unsigned(6506, LUT_AMPL_WIDTH - 1),
		30684 => to_unsigned(6503, LUT_AMPL_WIDTH - 1),
		30685 => to_unsigned(6500, LUT_AMPL_WIDTH - 1),
		30686 => to_unsigned(6497, LUT_AMPL_WIDTH - 1),
		30687 => to_unsigned(6494, LUT_AMPL_WIDTH - 1),
		30688 => to_unsigned(6491, LUT_AMPL_WIDTH - 1),
		30689 => to_unsigned(6488, LUT_AMPL_WIDTH - 1),
		30690 => to_unsigned(6485, LUT_AMPL_WIDTH - 1),
		30691 => to_unsigned(6482, LUT_AMPL_WIDTH - 1),
		30692 => to_unsigned(6479, LUT_AMPL_WIDTH - 1),
		30693 => to_unsigned(6476, LUT_AMPL_WIDTH - 1),
		30694 => to_unsigned(6473, LUT_AMPL_WIDTH - 1),
		30695 => to_unsigned(6470, LUT_AMPL_WIDTH - 1),
		30696 => to_unsigned(6466, LUT_AMPL_WIDTH - 1),
		30697 => to_unsigned(6463, LUT_AMPL_WIDTH - 1),
		30698 => to_unsigned(6460, LUT_AMPL_WIDTH - 1),
		30699 => to_unsigned(6457, LUT_AMPL_WIDTH - 1),
		30700 => to_unsigned(6454, LUT_AMPL_WIDTH - 1),
		30701 => to_unsigned(6451, LUT_AMPL_WIDTH - 1),
		30702 => to_unsigned(6448, LUT_AMPL_WIDTH - 1),
		30703 => to_unsigned(6445, LUT_AMPL_WIDTH - 1),
		30704 => to_unsigned(6442, LUT_AMPL_WIDTH - 1),
		30705 => to_unsigned(6439, LUT_AMPL_WIDTH - 1),
		30706 => to_unsigned(6436, LUT_AMPL_WIDTH - 1),
		30707 => to_unsigned(6433, LUT_AMPL_WIDTH - 1),
		30708 => to_unsigned(6429, LUT_AMPL_WIDTH - 1),
		30709 => to_unsigned(6426, LUT_AMPL_WIDTH - 1),
		30710 => to_unsigned(6423, LUT_AMPL_WIDTH - 1),
		30711 => to_unsigned(6420, LUT_AMPL_WIDTH - 1),
		30712 => to_unsigned(6417, LUT_AMPL_WIDTH - 1),
		30713 => to_unsigned(6414, LUT_AMPL_WIDTH - 1),
		30714 => to_unsigned(6411, LUT_AMPL_WIDTH - 1),
		30715 => to_unsigned(6408, LUT_AMPL_WIDTH - 1),
		30716 => to_unsigned(6405, LUT_AMPL_WIDTH - 1),
		30717 => to_unsigned(6402, LUT_AMPL_WIDTH - 1),
		30718 => to_unsigned(6399, LUT_AMPL_WIDTH - 1),
		30719 => to_unsigned(6396, LUT_AMPL_WIDTH - 1),
		30720 => to_unsigned(6393, LUT_AMPL_WIDTH - 1),
		30721 => to_unsigned(6389, LUT_AMPL_WIDTH - 1),
		30722 => to_unsigned(6386, LUT_AMPL_WIDTH - 1),
		30723 => to_unsigned(6383, LUT_AMPL_WIDTH - 1),
		30724 => to_unsigned(6380, LUT_AMPL_WIDTH - 1),
		30725 => to_unsigned(6377, LUT_AMPL_WIDTH - 1),
		30726 => to_unsigned(6374, LUT_AMPL_WIDTH - 1),
		30727 => to_unsigned(6371, LUT_AMPL_WIDTH - 1),
		30728 => to_unsigned(6368, LUT_AMPL_WIDTH - 1),
		30729 => to_unsigned(6365, LUT_AMPL_WIDTH - 1),
		30730 => to_unsigned(6362, LUT_AMPL_WIDTH - 1),
		30731 => to_unsigned(6359, LUT_AMPL_WIDTH - 1),
		30732 => to_unsigned(6356, LUT_AMPL_WIDTH - 1),
		30733 => to_unsigned(6352, LUT_AMPL_WIDTH - 1),
		30734 => to_unsigned(6349, LUT_AMPL_WIDTH - 1),
		30735 => to_unsigned(6346, LUT_AMPL_WIDTH - 1),
		30736 => to_unsigned(6343, LUT_AMPL_WIDTH - 1),
		30737 => to_unsigned(6340, LUT_AMPL_WIDTH - 1),
		30738 => to_unsigned(6337, LUT_AMPL_WIDTH - 1),
		30739 => to_unsigned(6334, LUT_AMPL_WIDTH - 1),
		30740 => to_unsigned(6331, LUT_AMPL_WIDTH - 1),
		30741 => to_unsigned(6328, LUT_AMPL_WIDTH - 1),
		30742 => to_unsigned(6325, LUT_AMPL_WIDTH - 1),
		30743 => to_unsigned(6322, LUT_AMPL_WIDTH - 1),
		30744 => to_unsigned(6319, LUT_AMPL_WIDTH - 1),
		30745 => to_unsigned(6315, LUT_AMPL_WIDTH - 1),
		30746 => to_unsigned(6312, LUT_AMPL_WIDTH - 1),
		30747 => to_unsigned(6309, LUT_AMPL_WIDTH - 1),
		30748 => to_unsigned(6306, LUT_AMPL_WIDTH - 1),
		30749 => to_unsigned(6303, LUT_AMPL_WIDTH - 1),
		30750 => to_unsigned(6300, LUT_AMPL_WIDTH - 1),
		30751 => to_unsigned(6297, LUT_AMPL_WIDTH - 1),
		30752 => to_unsigned(6294, LUT_AMPL_WIDTH - 1),
		30753 => to_unsigned(6291, LUT_AMPL_WIDTH - 1),
		30754 => to_unsigned(6288, LUT_AMPL_WIDTH - 1),
		30755 => to_unsigned(6285, LUT_AMPL_WIDTH - 1),
		30756 => to_unsigned(6282, LUT_AMPL_WIDTH - 1),
		30757 => to_unsigned(6278, LUT_AMPL_WIDTH - 1),
		30758 => to_unsigned(6275, LUT_AMPL_WIDTH - 1),
		30759 => to_unsigned(6272, LUT_AMPL_WIDTH - 1),
		30760 => to_unsigned(6269, LUT_AMPL_WIDTH - 1),
		30761 => to_unsigned(6266, LUT_AMPL_WIDTH - 1),
		30762 => to_unsigned(6263, LUT_AMPL_WIDTH - 1),
		30763 => to_unsigned(6260, LUT_AMPL_WIDTH - 1),
		30764 => to_unsigned(6257, LUT_AMPL_WIDTH - 1),
		30765 => to_unsigned(6254, LUT_AMPL_WIDTH - 1),
		30766 => to_unsigned(6251, LUT_AMPL_WIDTH - 1),
		30767 => to_unsigned(6248, LUT_AMPL_WIDTH - 1),
		30768 => to_unsigned(6245, LUT_AMPL_WIDTH - 1),
		30769 => to_unsigned(6241, LUT_AMPL_WIDTH - 1),
		30770 => to_unsigned(6238, LUT_AMPL_WIDTH - 1),
		30771 => to_unsigned(6235, LUT_AMPL_WIDTH - 1),
		30772 => to_unsigned(6232, LUT_AMPL_WIDTH - 1),
		30773 => to_unsigned(6229, LUT_AMPL_WIDTH - 1),
		30774 => to_unsigned(6226, LUT_AMPL_WIDTH - 1),
		30775 => to_unsigned(6223, LUT_AMPL_WIDTH - 1),
		30776 => to_unsigned(6220, LUT_AMPL_WIDTH - 1),
		30777 => to_unsigned(6217, LUT_AMPL_WIDTH - 1),
		30778 => to_unsigned(6214, LUT_AMPL_WIDTH - 1),
		30779 => to_unsigned(6211, LUT_AMPL_WIDTH - 1),
		30780 => to_unsigned(6208, LUT_AMPL_WIDTH - 1),
		30781 => to_unsigned(6204, LUT_AMPL_WIDTH - 1),
		30782 => to_unsigned(6201, LUT_AMPL_WIDTH - 1),
		30783 => to_unsigned(6198, LUT_AMPL_WIDTH - 1),
		30784 => to_unsigned(6195, LUT_AMPL_WIDTH - 1),
		30785 => to_unsigned(6192, LUT_AMPL_WIDTH - 1),
		30786 => to_unsigned(6189, LUT_AMPL_WIDTH - 1),
		30787 => to_unsigned(6186, LUT_AMPL_WIDTH - 1),
		30788 => to_unsigned(6183, LUT_AMPL_WIDTH - 1),
		30789 => to_unsigned(6180, LUT_AMPL_WIDTH - 1),
		30790 => to_unsigned(6177, LUT_AMPL_WIDTH - 1),
		30791 => to_unsigned(6174, LUT_AMPL_WIDTH - 1),
		30792 => to_unsigned(6171, LUT_AMPL_WIDTH - 1),
		30793 => to_unsigned(6167, LUT_AMPL_WIDTH - 1),
		30794 => to_unsigned(6164, LUT_AMPL_WIDTH - 1),
		30795 => to_unsigned(6161, LUT_AMPL_WIDTH - 1),
		30796 => to_unsigned(6158, LUT_AMPL_WIDTH - 1),
		30797 => to_unsigned(6155, LUT_AMPL_WIDTH - 1),
		30798 => to_unsigned(6152, LUT_AMPL_WIDTH - 1),
		30799 => to_unsigned(6149, LUT_AMPL_WIDTH - 1),
		30800 => to_unsigned(6146, LUT_AMPL_WIDTH - 1),
		30801 => to_unsigned(6143, LUT_AMPL_WIDTH - 1),
		30802 => to_unsigned(6140, LUT_AMPL_WIDTH - 1),
		30803 => to_unsigned(6137, LUT_AMPL_WIDTH - 1),
		30804 => to_unsigned(6134, LUT_AMPL_WIDTH - 1),
		30805 => to_unsigned(6130, LUT_AMPL_WIDTH - 1),
		30806 => to_unsigned(6127, LUT_AMPL_WIDTH - 1),
		30807 => to_unsigned(6124, LUT_AMPL_WIDTH - 1),
		30808 => to_unsigned(6121, LUT_AMPL_WIDTH - 1),
		30809 => to_unsigned(6118, LUT_AMPL_WIDTH - 1),
		30810 => to_unsigned(6115, LUT_AMPL_WIDTH - 1),
		30811 => to_unsigned(6112, LUT_AMPL_WIDTH - 1),
		30812 => to_unsigned(6109, LUT_AMPL_WIDTH - 1),
		30813 => to_unsigned(6106, LUT_AMPL_WIDTH - 1),
		30814 => to_unsigned(6103, LUT_AMPL_WIDTH - 1),
		30815 => to_unsigned(6100, LUT_AMPL_WIDTH - 1),
		30816 => to_unsigned(6096, LUT_AMPL_WIDTH - 1),
		30817 => to_unsigned(6093, LUT_AMPL_WIDTH - 1),
		30818 => to_unsigned(6090, LUT_AMPL_WIDTH - 1),
		30819 => to_unsigned(6087, LUT_AMPL_WIDTH - 1),
		30820 => to_unsigned(6084, LUT_AMPL_WIDTH - 1),
		30821 => to_unsigned(6081, LUT_AMPL_WIDTH - 1),
		30822 => to_unsigned(6078, LUT_AMPL_WIDTH - 1),
		30823 => to_unsigned(6075, LUT_AMPL_WIDTH - 1),
		30824 => to_unsigned(6072, LUT_AMPL_WIDTH - 1),
		30825 => to_unsigned(6069, LUT_AMPL_WIDTH - 1),
		30826 => to_unsigned(6066, LUT_AMPL_WIDTH - 1),
		30827 => to_unsigned(6063, LUT_AMPL_WIDTH - 1),
		30828 => to_unsigned(6059, LUT_AMPL_WIDTH - 1),
		30829 => to_unsigned(6056, LUT_AMPL_WIDTH - 1),
		30830 => to_unsigned(6053, LUT_AMPL_WIDTH - 1),
		30831 => to_unsigned(6050, LUT_AMPL_WIDTH - 1),
		30832 => to_unsigned(6047, LUT_AMPL_WIDTH - 1),
		30833 => to_unsigned(6044, LUT_AMPL_WIDTH - 1),
		30834 => to_unsigned(6041, LUT_AMPL_WIDTH - 1),
		30835 => to_unsigned(6038, LUT_AMPL_WIDTH - 1),
		30836 => to_unsigned(6035, LUT_AMPL_WIDTH - 1),
		30837 => to_unsigned(6032, LUT_AMPL_WIDTH - 1),
		30838 => to_unsigned(6029, LUT_AMPL_WIDTH - 1),
		30839 => to_unsigned(6025, LUT_AMPL_WIDTH - 1),
		30840 => to_unsigned(6022, LUT_AMPL_WIDTH - 1),
		30841 => to_unsigned(6019, LUT_AMPL_WIDTH - 1),
		30842 => to_unsigned(6016, LUT_AMPL_WIDTH - 1),
		30843 => to_unsigned(6013, LUT_AMPL_WIDTH - 1),
		30844 => to_unsigned(6010, LUT_AMPL_WIDTH - 1),
		30845 => to_unsigned(6007, LUT_AMPL_WIDTH - 1),
		30846 => to_unsigned(6004, LUT_AMPL_WIDTH - 1),
		30847 => to_unsigned(6001, LUT_AMPL_WIDTH - 1),
		30848 => to_unsigned(5998, LUT_AMPL_WIDTH - 1),
		30849 => to_unsigned(5995, LUT_AMPL_WIDTH - 1),
		30850 => to_unsigned(5991, LUT_AMPL_WIDTH - 1),
		30851 => to_unsigned(5988, LUT_AMPL_WIDTH - 1),
		30852 => to_unsigned(5985, LUT_AMPL_WIDTH - 1),
		30853 => to_unsigned(5982, LUT_AMPL_WIDTH - 1),
		30854 => to_unsigned(5979, LUT_AMPL_WIDTH - 1),
		30855 => to_unsigned(5976, LUT_AMPL_WIDTH - 1),
		30856 => to_unsigned(5973, LUT_AMPL_WIDTH - 1),
		30857 => to_unsigned(5970, LUT_AMPL_WIDTH - 1),
		30858 => to_unsigned(5967, LUT_AMPL_WIDTH - 1),
		30859 => to_unsigned(5964, LUT_AMPL_WIDTH - 1),
		30860 => to_unsigned(5961, LUT_AMPL_WIDTH - 1),
		30861 => to_unsigned(5958, LUT_AMPL_WIDTH - 1),
		30862 => to_unsigned(5954, LUT_AMPL_WIDTH - 1),
		30863 => to_unsigned(5951, LUT_AMPL_WIDTH - 1),
		30864 => to_unsigned(5948, LUT_AMPL_WIDTH - 1),
		30865 => to_unsigned(5945, LUT_AMPL_WIDTH - 1),
		30866 => to_unsigned(5942, LUT_AMPL_WIDTH - 1),
		30867 => to_unsigned(5939, LUT_AMPL_WIDTH - 1),
		30868 => to_unsigned(5936, LUT_AMPL_WIDTH - 1),
		30869 => to_unsigned(5933, LUT_AMPL_WIDTH - 1),
		30870 => to_unsigned(5930, LUT_AMPL_WIDTH - 1),
		30871 => to_unsigned(5927, LUT_AMPL_WIDTH - 1),
		30872 => to_unsigned(5924, LUT_AMPL_WIDTH - 1),
		30873 => to_unsigned(5920, LUT_AMPL_WIDTH - 1),
		30874 => to_unsigned(5917, LUT_AMPL_WIDTH - 1),
		30875 => to_unsigned(5914, LUT_AMPL_WIDTH - 1),
		30876 => to_unsigned(5911, LUT_AMPL_WIDTH - 1),
		30877 => to_unsigned(5908, LUT_AMPL_WIDTH - 1),
		30878 => to_unsigned(5905, LUT_AMPL_WIDTH - 1),
		30879 => to_unsigned(5902, LUT_AMPL_WIDTH - 1),
		30880 => to_unsigned(5899, LUT_AMPL_WIDTH - 1),
		30881 => to_unsigned(5896, LUT_AMPL_WIDTH - 1),
		30882 => to_unsigned(5893, LUT_AMPL_WIDTH - 1),
		30883 => to_unsigned(5890, LUT_AMPL_WIDTH - 1),
		30884 => to_unsigned(5886, LUT_AMPL_WIDTH - 1),
		30885 => to_unsigned(5883, LUT_AMPL_WIDTH - 1),
		30886 => to_unsigned(5880, LUT_AMPL_WIDTH - 1),
		30887 => to_unsigned(5877, LUT_AMPL_WIDTH - 1),
		30888 => to_unsigned(5874, LUT_AMPL_WIDTH - 1),
		30889 => to_unsigned(5871, LUT_AMPL_WIDTH - 1),
		30890 => to_unsigned(5868, LUT_AMPL_WIDTH - 1),
		30891 => to_unsigned(5865, LUT_AMPL_WIDTH - 1),
		30892 => to_unsigned(5862, LUT_AMPL_WIDTH - 1),
		30893 => to_unsigned(5859, LUT_AMPL_WIDTH - 1),
		30894 => to_unsigned(5856, LUT_AMPL_WIDTH - 1),
		30895 => to_unsigned(5852, LUT_AMPL_WIDTH - 1),
		30896 => to_unsigned(5849, LUT_AMPL_WIDTH - 1),
		30897 => to_unsigned(5846, LUT_AMPL_WIDTH - 1),
		30898 => to_unsigned(5843, LUT_AMPL_WIDTH - 1),
		30899 => to_unsigned(5840, LUT_AMPL_WIDTH - 1),
		30900 => to_unsigned(5837, LUT_AMPL_WIDTH - 1),
		30901 => to_unsigned(5834, LUT_AMPL_WIDTH - 1),
		30902 => to_unsigned(5831, LUT_AMPL_WIDTH - 1),
		30903 => to_unsigned(5828, LUT_AMPL_WIDTH - 1),
		30904 => to_unsigned(5825, LUT_AMPL_WIDTH - 1),
		30905 => to_unsigned(5822, LUT_AMPL_WIDTH - 1),
		30906 => to_unsigned(5818, LUT_AMPL_WIDTH - 1),
		30907 => to_unsigned(5815, LUT_AMPL_WIDTH - 1),
		30908 => to_unsigned(5812, LUT_AMPL_WIDTH - 1),
		30909 => to_unsigned(5809, LUT_AMPL_WIDTH - 1),
		30910 => to_unsigned(5806, LUT_AMPL_WIDTH - 1),
		30911 => to_unsigned(5803, LUT_AMPL_WIDTH - 1),
		30912 => to_unsigned(5800, LUT_AMPL_WIDTH - 1),
		30913 => to_unsigned(5797, LUT_AMPL_WIDTH - 1),
		30914 => to_unsigned(5794, LUT_AMPL_WIDTH - 1),
		30915 => to_unsigned(5791, LUT_AMPL_WIDTH - 1),
		30916 => to_unsigned(5788, LUT_AMPL_WIDTH - 1),
		30917 => to_unsigned(5784, LUT_AMPL_WIDTH - 1),
		30918 => to_unsigned(5781, LUT_AMPL_WIDTH - 1),
		30919 => to_unsigned(5778, LUT_AMPL_WIDTH - 1),
		30920 => to_unsigned(5775, LUT_AMPL_WIDTH - 1),
		30921 => to_unsigned(5772, LUT_AMPL_WIDTH - 1),
		30922 => to_unsigned(5769, LUT_AMPL_WIDTH - 1),
		30923 => to_unsigned(5766, LUT_AMPL_WIDTH - 1),
		30924 => to_unsigned(5763, LUT_AMPL_WIDTH - 1),
		30925 => to_unsigned(5760, LUT_AMPL_WIDTH - 1),
		30926 => to_unsigned(5757, LUT_AMPL_WIDTH - 1),
		30927 => to_unsigned(5754, LUT_AMPL_WIDTH - 1),
		30928 => to_unsigned(5750, LUT_AMPL_WIDTH - 1),
		30929 => to_unsigned(5747, LUT_AMPL_WIDTH - 1),
		30930 => to_unsigned(5744, LUT_AMPL_WIDTH - 1),
		30931 => to_unsigned(5741, LUT_AMPL_WIDTH - 1),
		30932 => to_unsigned(5738, LUT_AMPL_WIDTH - 1),
		30933 => to_unsigned(5735, LUT_AMPL_WIDTH - 1),
		30934 => to_unsigned(5732, LUT_AMPL_WIDTH - 1),
		30935 => to_unsigned(5729, LUT_AMPL_WIDTH - 1),
		30936 => to_unsigned(5726, LUT_AMPL_WIDTH - 1),
		30937 => to_unsigned(5723, LUT_AMPL_WIDTH - 1),
		30938 => to_unsigned(5719, LUT_AMPL_WIDTH - 1),
		30939 => to_unsigned(5716, LUT_AMPL_WIDTH - 1),
		30940 => to_unsigned(5713, LUT_AMPL_WIDTH - 1),
		30941 => to_unsigned(5710, LUT_AMPL_WIDTH - 1),
		30942 => to_unsigned(5707, LUT_AMPL_WIDTH - 1),
		30943 => to_unsigned(5704, LUT_AMPL_WIDTH - 1),
		30944 => to_unsigned(5701, LUT_AMPL_WIDTH - 1),
		30945 => to_unsigned(5698, LUT_AMPL_WIDTH - 1),
		30946 => to_unsigned(5695, LUT_AMPL_WIDTH - 1),
		30947 => to_unsigned(5692, LUT_AMPL_WIDTH - 1),
		30948 => to_unsigned(5689, LUT_AMPL_WIDTH - 1),
		30949 => to_unsigned(5685, LUT_AMPL_WIDTH - 1),
		30950 => to_unsigned(5682, LUT_AMPL_WIDTH - 1),
		30951 => to_unsigned(5679, LUT_AMPL_WIDTH - 1),
		30952 => to_unsigned(5676, LUT_AMPL_WIDTH - 1),
		30953 => to_unsigned(5673, LUT_AMPL_WIDTH - 1),
		30954 => to_unsigned(5670, LUT_AMPL_WIDTH - 1),
		30955 => to_unsigned(5667, LUT_AMPL_WIDTH - 1),
		30956 => to_unsigned(5664, LUT_AMPL_WIDTH - 1),
		30957 => to_unsigned(5661, LUT_AMPL_WIDTH - 1),
		30958 => to_unsigned(5658, LUT_AMPL_WIDTH - 1),
		30959 => to_unsigned(5655, LUT_AMPL_WIDTH - 1),
		30960 => to_unsigned(5651, LUT_AMPL_WIDTH - 1),
		30961 => to_unsigned(5648, LUT_AMPL_WIDTH - 1),
		30962 => to_unsigned(5645, LUT_AMPL_WIDTH - 1),
		30963 => to_unsigned(5642, LUT_AMPL_WIDTH - 1),
		30964 => to_unsigned(5639, LUT_AMPL_WIDTH - 1),
		30965 => to_unsigned(5636, LUT_AMPL_WIDTH - 1),
		30966 => to_unsigned(5633, LUT_AMPL_WIDTH - 1),
		30967 => to_unsigned(5630, LUT_AMPL_WIDTH - 1),
		30968 => to_unsigned(5627, LUT_AMPL_WIDTH - 1),
		30969 => to_unsigned(5624, LUT_AMPL_WIDTH - 1),
		30970 => to_unsigned(5620, LUT_AMPL_WIDTH - 1),
		30971 => to_unsigned(5617, LUT_AMPL_WIDTH - 1),
		30972 => to_unsigned(5614, LUT_AMPL_WIDTH - 1),
		30973 => to_unsigned(5611, LUT_AMPL_WIDTH - 1),
		30974 => to_unsigned(5608, LUT_AMPL_WIDTH - 1),
		30975 => to_unsigned(5605, LUT_AMPL_WIDTH - 1),
		30976 => to_unsigned(5602, LUT_AMPL_WIDTH - 1),
		30977 => to_unsigned(5599, LUT_AMPL_WIDTH - 1),
		30978 => to_unsigned(5596, LUT_AMPL_WIDTH - 1),
		30979 => to_unsigned(5593, LUT_AMPL_WIDTH - 1),
		30980 => to_unsigned(5590, LUT_AMPL_WIDTH - 1),
		30981 => to_unsigned(5586, LUT_AMPL_WIDTH - 1),
		30982 => to_unsigned(5583, LUT_AMPL_WIDTH - 1),
		30983 => to_unsigned(5580, LUT_AMPL_WIDTH - 1),
		30984 => to_unsigned(5577, LUT_AMPL_WIDTH - 1),
		30985 => to_unsigned(5574, LUT_AMPL_WIDTH - 1),
		30986 => to_unsigned(5571, LUT_AMPL_WIDTH - 1),
		30987 => to_unsigned(5568, LUT_AMPL_WIDTH - 1),
		30988 => to_unsigned(5565, LUT_AMPL_WIDTH - 1),
		30989 => to_unsigned(5562, LUT_AMPL_WIDTH - 1),
		30990 => to_unsigned(5559, LUT_AMPL_WIDTH - 1),
		30991 => to_unsigned(5555, LUT_AMPL_WIDTH - 1),
		30992 => to_unsigned(5552, LUT_AMPL_WIDTH - 1),
		30993 => to_unsigned(5549, LUT_AMPL_WIDTH - 1),
		30994 => to_unsigned(5546, LUT_AMPL_WIDTH - 1),
		30995 => to_unsigned(5543, LUT_AMPL_WIDTH - 1),
		30996 => to_unsigned(5540, LUT_AMPL_WIDTH - 1),
		30997 => to_unsigned(5537, LUT_AMPL_WIDTH - 1),
		30998 => to_unsigned(5534, LUT_AMPL_WIDTH - 1),
		30999 => to_unsigned(5531, LUT_AMPL_WIDTH - 1),
		31000 => to_unsigned(5528, LUT_AMPL_WIDTH - 1),
		31001 => to_unsigned(5525, LUT_AMPL_WIDTH - 1),
		31002 => to_unsigned(5521, LUT_AMPL_WIDTH - 1),
		31003 => to_unsigned(5518, LUT_AMPL_WIDTH - 1),
		31004 => to_unsigned(5515, LUT_AMPL_WIDTH - 1),
		31005 => to_unsigned(5512, LUT_AMPL_WIDTH - 1),
		31006 => to_unsigned(5509, LUT_AMPL_WIDTH - 1),
		31007 => to_unsigned(5506, LUT_AMPL_WIDTH - 1),
		31008 => to_unsigned(5503, LUT_AMPL_WIDTH - 1),
		31009 => to_unsigned(5500, LUT_AMPL_WIDTH - 1),
		31010 => to_unsigned(5497, LUT_AMPL_WIDTH - 1),
		31011 => to_unsigned(5494, LUT_AMPL_WIDTH - 1),
		31012 => to_unsigned(5490, LUT_AMPL_WIDTH - 1),
		31013 => to_unsigned(5487, LUT_AMPL_WIDTH - 1),
		31014 => to_unsigned(5484, LUT_AMPL_WIDTH - 1),
		31015 => to_unsigned(5481, LUT_AMPL_WIDTH - 1),
		31016 => to_unsigned(5478, LUT_AMPL_WIDTH - 1),
		31017 => to_unsigned(5475, LUT_AMPL_WIDTH - 1),
		31018 => to_unsigned(5472, LUT_AMPL_WIDTH - 1),
		31019 => to_unsigned(5469, LUT_AMPL_WIDTH - 1),
		31020 => to_unsigned(5466, LUT_AMPL_WIDTH - 1),
		31021 => to_unsigned(5463, LUT_AMPL_WIDTH - 1),
		31022 => to_unsigned(5459, LUT_AMPL_WIDTH - 1),
		31023 => to_unsigned(5456, LUT_AMPL_WIDTH - 1),
		31024 => to_unsigned(5453, LUT_AMPL_WIDTH - 1),
		31025 => to_unsigned(5450, LUT_AMPL_WIDTH - 1),
		31026 => to_unsigned(5447, LUT_AMPL_WIDTH - 1),
		31027 => to_unsigned(5444, LUT_AMPL_WIDTH - 1),
		31028 => to_unsigned(5441, LUT_AMPL_WIDTH - 1),
		31029 => to_unsigned(5438, LUT_AMPL_WIDTH - 1),
		31030 => to_unsigned(5435, LUT_AMPL_WIDTH - 1),
		31031 => to_unsigned(5432, LUT_AMPL_WIDTH - 1),
		31032 => to_unsigned(5428, LUT_AMPL_WIDTH - 1),
		31033 => to_unsigned(5425, LUT_AMPL_WIDTH - 1),
		31034 => to_unsigned(5422, LUT_AMPL_WIDTH - 1),
		31035 => to_unsigned(5419, LUT_AMPL_WIDTH - 1),
		31036 => to_unsigned(5416, LUT_AMPL_WIDTH - 1),
		31037 => to_unsigned(5413, LUT_AMPL_WIDTH - 1),
		31038 => to_unsigned(5410, LUT_AMPL_WIDTH - 1),
		31039 => to_unsigned(5407, LUT_AMPL_WIDTH - 1),
		31040 => to_unsigned(5404, LUT_AMPL_WIDTH - 1),
		31041 => to_unsigned(5401, LUT_AMPL_WIDTH - 1),
		31042 => to_unsigned(5398, LUT_AMPL_WIDTH - 1),
		31043 => to_unsigned(5394, LUT_AMPL_WIDTH - 1),
		31044 => to_unsigned(5391, LUT_AMPL_WIDTH - 1),
		31045 => to_unsigned(5388, LUT_AMPL_WIDTH - 1),
		31046 => to_unsigned(5385, LUT_AMPL_WIDTH - 1),
		31047 => to_unsigned(5382, LUT_AMPL_WIDTH - 1),
		31048 => to_unsigned(5379, LUT_AMPL_WIDTH - 1),
		31049 => to_unsigned(5376, LUT_AMPL_WIDTH - 1),
		31050 => to_unsigned(5373, LUT_AMPL_WIDTH - 1),
		31051 => to_unsigned(5370, LUT_AMPL_WIDTH - 1),
		31052 => to_unsigned(5367, LUT_AMPL_WIDTH - 1),
		31053 => to_unsigned(5363, LUT_AMPL_WIDTH - 1),
		31054 => to_unsigned(5360, LUT_AMPL_WIDTH - 1),
		31055 => to_unsigned(5357, LUT_AMPL_WIDTH - 1),
		31056 => to_unsigned(5354, LUT_AMPL_WIDTH - 1),
		31057 => to_unsigned(5351, LUT_AMPL_WIDTH - 1),
		31058 => to_unsigned(5348, LUT_AMPL_WIDTH - 1),
		31059 => to_unsigned(5345, LUT_AMPL_WIDTH - 1),
		31060 => to_unsigned(5342, LUT_AMPL_WIDTH - 1),
		31061 => to_unsigned(5339, LUT_AMPL_WIDTH - 1),
		31062 => to_unsigned(5336, LUT_AMPL_WIDTH - 1),
		31063 => to_unsigned(5332, LUT_AMPL_WIDTH - 1),
		31064 => to_unsigned(5329, LUT_AMPL_WIDTH - 1),
		31065 => to_unsigned(5326, LUT_AMPL_WIDTH - 1),
		31066 => to_unsigned(5323, LUT_AMPL_WIDTH - 1),
		31067 => to_unsigned(5320, LUT_AMPL_WIDTH - 1),
		31068 => to_unsigned(5317, LUT_AMPL_WIDTH - 1),
		31069 => to_unsigned(5314, LUT_AMPL_WIDTH - 1),
		31070 => to_unsigned(5311, LUT_AMPL_WIDTH - 1),
		31071 => to_unsigned(5308, LUT_AMPL_WIDTH - 1),
		31072 => to_unsigned(5305, LUT_AMPL_WIDTH - 1),
		31073 => to_unsigned(5301, LUT_AMPL_WIDTH - 1),
		31074 => to_unsigned(5298, LUT_AMPL_WIDTH - 1),
		31075 => to_unsigned(5295, LUT_AMPL_WIDTH - 1),
		31076 => to_unsigned(5292, LUT_AMPL_WIDTH - 1),
		31077 => to_unsigned(5289, LUT_AMPL_WIDTH - 1),
		31078 => to_unsigned(5286, LUT_AMPL_WIDTH - 1),
		31079 => to_unsigned(5283, LUT_AMPL_WIDTH - 1),
		31080 => to_unsigned(5280, LUT_AMPL_WIDTH - 1),
		31081 => to_unsigned(5277, LUT_AMPL_WIDTH - 1),
		31082 => to_unsigned(5274, LUT_AMPL_WIDTH - 1),
		31083 => to_unsigned(5270, LUT_AMPL_WIDTH - 1),
		31084 => to_unsigned(5267, LUT_AMPL_WIDTH - 1),
		31085 => to_unsigned(5264, LUT_AMPL_WIDTH - 1),
		31086 => to_unsigned(5261, LUT_AMPL_WIDTH - 1),
		31087 => to_unsigned(5258, LUT_AMPL_WIDTH - 1),
		31088 => to_unsigned(5255, LUT_AMPL_WIDTH - 1),
		31089 => to_unsigned(5252, LUT_AMPL_WIDTH - 1),
		31090 => to_unsigned(5249, LUT_AMPL_WIDTH - 1),
		31091 => to_unsigned(5246, LUT_AMPL_WIDTH - 1),
		31092 => to_unsigned(5243, LUT_AMPL_WIDTH - 1),
		31093 => to_unsigned(5239, LUT_AMPL_WIDTH - 1),
		31094 => to_unsigned(5236, LUT_AMPL_WIDTH - 1),
		31095 => to_unsigned(5233, LUT_AMPL_WIDTH - 1),
		31096 => to_unsigned(5230, LUT_AMPL_WIDTH - 1),
		31097 => to_unsigned(5227, LUT_AMPL_WIDTH - 1),
		31098 => to_unsigned(5224, LUT_AMPL_WIDTH - 1),
		31099 => to_unsigned(5221, LUT_AMPL_WIDTH - 1),
		31100 => to_unsigned(5218, LUT_AMPL_WIDTH - 1),
		31101 => to_unsigned(5215, LUT_AMPL_WIDTH - 1),
		31102 => to_unsigned(5212, LUT_AMPL_WIDTH - 1),
		31103 => to_unsigned(5208, LUT_AMPL_WIDTH - 1),
		31104 => to_unsigned(5205, LUT_AMPL_WIDTH - 1),
		31105 => to_unsigned(5202, LUT_AMPL_WIDTH - 1),
		31106 => to_unsigned(5199, LUT_AMPL_WIDTH - 1),
		31107 => to_unsigned(5196, LUT_AMPL_WIDTH - 1),
		31108 => to_unsigned(5193, LUT_AMPL_WIDTH - 1),
		31109 => to_unsigned(5190, LUT_AMPL_WIDTH - 1),
		31110 => to_unsigned(5187, LUT_AMPL_WIDTH - 1),
		31111 => to_unsigned(5184, LUT_AMPL_WIDTH - 1),
		31112 => to_unsigned(5180, LUT_AMPL_WIDTH - 1),
		31113 => to_unsigned(5177, LUT_AMPL_WIDTH - 1),
		31114 => to_unsigned(5174, LUT_AMPL_WIDTH - 1),
		31115 => to_unsigned(5171, LUT_AMPL_WIDTH - 1),
		31116 => to_unsigned(5168, LUT_AMPL_WIDTH - 1),
		31117 => to_unsigned(5165, LUT_AMPL_WIDTH - 1),
		31118 => to_unsigned(5162, LUT_AMPL_WIDTH - 1),
		31119 => to_unsigned(5159, LUT_AMPL_WIDTH - 1),
		31120 => to_unsigned(5156, LUT_AMPL_WIDTH - 1),
		31121 => to_unsigned(5153, LUT_AMPL_WIDTH - 1),
		31122 => to_unsigned(5149, LUT_AMPL_WIDTH - 1),
		31123 => to_unsigned(5146, LUT_AMPL_WIDTH - 1),
		31124 => to_unsigned(5143, LUT_AMPL_WIDTH - 1),
		31125 => to_unsigned(5140, LUT_AMPL_WIDTH - 1),
		31126 => to_unsigned(5137, LUT_AMPL_WIDTH - 1),
		31127 => to_unsigned(5134, LUT_AMPL_WIDTH - 1),
		31128 => to_unsigned(5131, LUT_AMPL_WIDTH - 1),
		31129 => to_unsigned(5128, LUT_AMPL_WIDTH - 1),
		31130 => to_unsigned(5125, LUT_AMPL_WIDTH - 1),
		31131 => to_unsigned(5122, LUT_AMPL_WIDTH - 1),
		31132 => to_unsigned(5118, LUT_AMPL_WIDTH - 1),
		31133 => to_unsigned(5115, LUT_AMPL_WIDTH - 1),
		31134 => to_unsigned(5112, LUT_AMPL_WIDTH - 1),
		31135 => to_unsigned(5109, LUT_AMPL_WIDTH - 1),
		31136 => to_unsigned(5106, LUT_AMPL_WIDTH - 1),
		31137 => to_unsigned(5103, LUT_AMPL_WIDTH - 1),
		31138 => to_unsigned(5100, LUT_AMPL_WIDTH - 1),
		31139 => to_unsigned(5097, LUT_AMPL_WIDTH - 1),
		31140 => to_unsigned(5094, LUT_AMPL_WIDTH - 1),
		31141 => to_unsigned(5091, LUT_AMPL_WIDTH - 1),
		31142 => to_unsigned(5087, LUT_AMPL_WIDTH - 1),
		31143 => to_unsigned(5084, LUT_AMPL_WIDTH - 1),
		31144 => to_unsigned(5081, LUT_AMPL_WIDTH - 1),
		31145 => to_unsigned(5078, LUT_AMPL_WIDTH - 1),
		31146 => to_unsigned(5075, LUT_AMPL_WIDTH - 1),
		31147 => to_unsigned(5072, LUT_AMPL_WIDTH - 1),
		31148 => to_unsigned(5069, LUT_AMPL_WIDTH - 1),
		31149 => to_unsigned(5066, LUT_AMPL_WIDTH - 1),
		31150 => to_unsigned(5063, LUT_AMPL_WIDTH - 1),
		31151 => to_unsigned(5059, LUT_AMPL_WIDTH - 1),
		31152 => to_unsigned(5056, LUT_AMPL_WIDTH - 1),
		31153 => to_unsigned(5053, LUT_AMPL_WIDTH - 1),
		31154 => to_unsigned(5050, LUT_AMPL_WIDTH - 1),
		31155 => to_unsigned(5047, LUT_AMPL_WIDTH - 1),
		31156 => to_unsigned(5044, LUT_AMPL_WIDTH - 1),
		31157 => to_unsigned(5041, LUT_AMPL_WIDTH - 1),
		31158 => to_unsigned(5038, LUT_AMPL_WIDTH - 1),
		31159 => to_unsigned(5035, LUT_AMPL_WIDTH - 1),
		31160 => to_unsigned(5032, LUT_AMPL_WIDTH - 1),
		31161 => to_unsigned(5028, LUT_AMPL_WIDTH - 1),
		31162 => to_unsigned(5025, LUT_AMPL_WIDTH - 1),
		31163 => to_unsigned(5022, LUT_AMPL_WIDTH - 1),
		31164 => to_unsigned(5019, LUT_AMPL_WIDTH - 1),
		31165 => to_unsigned(5016, LUT_AMPL_WIDTH - 1),
		31166 => to_unsigned(5013, LUT_AMPL_WIDTH - 1),
		31167 => to_unsigned(5010, LUT_AMPL_WIDTH - 1),
		31168 => to_unsigned(5007, LUT_AMPL_WIDTH - 1),
		31169 => to_unsigned(5004, LUT_AMPL_WIDTH - 1),
		31170 => to_unsigned(5000, LUT_AMPL_WIDTH - 1),
		31171 => to_unsigned(4997, LUT_AMPL_WIDTH - 1),
		31172 => to_unsigned(4994, LUT_AMPL_WIDTH - 1),
		31173 => to_unsigned(4991, LUT_AMPL_WIDTH - 1),
		31174 => to_unsigned(4988, LUT_AMPL_WIDTH - 1),
		31175 => to_unsigned(4985, LUT_AMPL_WIDTH - 1),
		31176 => to_unsigned(4982, LUT_AMPL_WIDTH - 1),
		31177 => to_unsigned(4979, LUT_AMPL_WIDTH - 1),
		31178 => to_unsigned(4976, LUT_AMPL_WIDTH - 1),
		31179 => to_unsigned(4973, LUT_AMPL_WIDTH - 1),
		31180 => to_unsigned(4969, LUT_AMPL_WIDTH - 1),
		31181 => to_unsigned(4966, LUT_AMPL_WIDTH - 1),
		31182 => to_unsigned(4963, LUT_AMPL_WIDTH - 1),
		31183 => to_unsigned(4960, LUT_AMPL_WIDTH - 1),
		31184 => to_unsigned(4957, LUT_AMPL_WIDTH - 1),
		31185 => to_unsigned(4954, LUT_AMPL_WIDTH - 1),
		31186 => to_unsigned(4951, LUT_AMPL_WIDTH - 1),
		31187 => to_unsigned(4948, LUT_AMPL_WIDTH - 1),
		31188 => to_unsigned(4945, LUT_AMPL_WIDTH - 1),
		31189 => to_unsigned(4941, LUT_AMPL_WIDTH - 1),
		31190 => to_unsigned(4938, LUT_AMPL_WIDTH - 1),
		31191 => to_unsigned(4935, LUT_AMPL_WIDTH - 1),
		31192 => to_unsigned(4932, LUT_AMPL_WIDTH - 1),
		31193 => to_unsigned(4929, LUT_AMPL_WIDTH - 1),
		31194 => to_unsigned(4926, LUT_AMPL_WIDTH - 1),
		31195 => to_unsigned(4923, LUT_AMPL_WIDTH - 1),
		31196 => to_unsigned(4920, LUT_AMPL_WIDTH - 1),
		31197 => to_unsigned(4917, LUT_AMPL_WIDTH - 1),
		31198 => to_unsigned(4914, LUT_AMPL_WIDTH - 1),
		31199 => to_unsigned(4910, LUT_AMPL_WIDTH - 1),
		31200 => to_unsigned(4907, LUT_AMPL_WIDTH - 1),
		31201 => to_unsigned(4904, LUT_AMPL_WIDTH - 1),
		31202 => to_unsigned(4901, LUT_AMPL_WIDTH - 1),
		31203 => to_unsigned(4898, LUT_AMPL_WIDTH - 1),
		31204 => to_unsigned(4895, LUT_AMPL_WIDTH - 1),
		31205 => to_unsigned(4892, LUT_AMPL_WIDTH - 1),
		31206 => to_unsigned(4889, LUT_AMPL_WIDTH - 1),
		31207 => to_unsigned(4886, LUT_AMPL_WIDTH - 1),
		31208 => to_unsigned(4882, LUT_AMPL_WIDTH - 1),
		31209 => to_unsigned(4879, LUT_AMPL_WIDTH - 1),
		31210 => to_unsigned(4876, LUT_AMPL_WIDTH - 1),
		31211 => to_unsigned(4873, LUT_AMPL_WIDTH - 1),
		31212 => to_unsigned(4870, LUT_AMPL_WIDTH - 1),
		31213 => to_unsigned(4867, LUT_AMPL_WIDTH - 1),
		31214 => to_unsigned(4864, LUT_AMPL_WIDTH - 1),
		31215 => to_unsigned(4861, LUT_AMPL_WIDTH - 1),
		31216 => to_unsigned(4858, LUT_AMPL_WIDTH - 1),
		31217 => to_unsigned(4855, LUT_AMPL_WIDTH - 1),
		31218 => to_unsigned(4851, LUT_AMPL_WIDTH - 1),
		31219 => to_unsigned(4848, LUT_AMPL_WIDTH - 1),
		31220 => to_unsigned(4845, LUT_AMPL_WIDTH - 1),
		31221 => to_unsigned(4842, LUT_AMPL_WIDTH - 1),
		31222 => to_unsigned(4839, LUT_AMPL_WIDTH - 1),
		31223 => to_unsigned(4836, LUT_AMPL_WIDTH - 1),
		31224 => to_unsigned(4833, LUT_AMPL_WIDTH - 1),
		31225 => to_unsigned(4830, LUT_AMPL_WIDTH - 1),
		31226 => to_unsigned(4827, LUT_AMPL_WIDTH - 1),
		31227 => to_unsigned(4823, LUT_AMPL_WIDTH - 1),
		31228 => to_unsigned(4820, LUT_AMPL_WIDTH - 1),
		31229 => to_unsigned(4817, LUT_AMPL_WIDTH - 1),
		31230 => to_unsigned(4814, LUT_AMPL_WIDTH - 1),
		31231 => to_unsigned(4811, LUT_AMPL_WIDTH - 1),
		31232 => to_unsigned(4808, LUT_AMPL_WIDTH - 1),
		31233 => to_unsigned(4805, LUT_AMPL_WIDTH - 1),
		31234 => to_unsigned(4802, LUT_AMPL_WIDTH - 1),
		31235 => to_unsigned(4799, LUT_AMPL_WIDTH - 1),
		31236 => to_unsigned(4795, LUT_AMPL_WIDTH - 1),
		31237 => to_unsigned(4792, LUT_AMPL_WIDTH - 1),
		31238 => to_unsigned(4789, LUT_AMPL_WIDTH - 1),
		31239 => to_unsigned(4786, LUT_AMPL_WIDTH - 1),
		31240 => to_unsigned(4783, LUT_AMPL_WIDTH - 1),
		31241 => to_unsigned(4780, LUT_AMPL_WIDTH - 1),
		31242 => to_unsigned(4777, LUT_AMPL_WIDTH - 1),
		31243 => to_unsigned(4774, LUT_AMPL_WIDTH - 1),
		31244 => to_unsigned(4771, LUT_AMPL_WIDTH - 1),
		31245 => to_unsigned(4768, LUT_AMPL_WIDTH - 1),
		31246 => to_unsigned(4764, LUT_AMPL_WIDTH - 1),
		31247 => to_unsigned(4761, LUT_AMPL_WIDTH - 1),
		31248 => to_unsigned(4758, LUT_AMPL_WIDTH - 1),
		31249 => to_unsigned(4755, LUT_AMPL_WIDTH - 1),
		31250 => to_unsigned(4752, LUT_AMPL_WIDTH - 1),
		31251 => to_unsigned(4749, LUT_AMPL_WIDTH - 1),
		31252 => to_unsigned(4746, LUT_AMPL_WIDTH - 1),
		31253 => to_unsigned(4743, LUT_AMPL_WIDTH - 1),
		31254 => to_unsigned(4740, LUT_AMPL_WIDTH - 1),
		31255 => to_unsigned(4736, LUT_AMPL_WIDTH - 1),
		31256 => to_unsigned(4733, LUT_AMPL_WIDTH - 1),
		31257 => to_unsigned(4730, LUT_AMPL_WIDTH - 1),
		31258 => to_unsigned(4727, LUT_AMPL_WIDTH - 1),
		31259 => to_unsigned(4724, LUT_AMPL_WIDTH - 1),
		31260 => to_unsigned(4721, LUT_AMPL_WIDTH - 1),
		31261 => to_unsigned(4718, LUT_AMPL_WIDTH - 1),
		31262 => to_unsigned(4715, LUT_AMPL_WIDTH - 1),
		31263 => to_unsigned(4712, LUT_AMPL_WIDTH - 1),
		31264 => to_unsigned(4708, LUT_AMPL_WIDTH - 1),
		31265 => to_unsigned(4705, LUT_AMPL_WIDTH - 1),
		31266 => to_unsigned(4702, LUT_AMPL_WIDTH - 1),
		31267 => to_unsigned(4699, LUT_AMPL_WIDTH - 1),
		31268 => to_unsigned(4696, LUT_AMPL_WIDTH - 1),
		31269 => to_unsigned(4693, LUT_AMPL_WIDTH - 1),
		31270 => to_unsigned(4690, LUT_AMPL_WIDTH - 1),
		31271 => to_unsigned(4687, LUT_AMPL_WIDTH - 1),
		31272 => to_unsigned(4684, LUT_AMPL_WIDTH - 1),
		31273 => to_unsigned(4680, LUT_AMPL_WIDTH - 1),
		31274 => to_unsigned(4677, LUT_AMPL_WIDTH - 1),
		31275 => to_unsigned(4674, LUT_AMPL_WIDTH - 1),
		31276 => to_unsigned(4671, LUT_AMPL_WIDTH - 1),
		31277 => to_unsigned(4668, LUT_AMPL_WIDTH - 1),
		31278 => to_unsigned(4665, LUT_AMPL_WIDTH - 1),
		31279 => to_unsigned(4662, LUT_AMPL_WIDTH - 1),
		31280 => to_unsigned(4659, LUT_AMPL_WIDTH - 1),
		31281 => to_unsigned(4656, LUT_AMPL_WIDTH - 1),
		31282 => to_unsigned(4652, LUT_AMPL_WIDTH - 1),
		31283 => to_unsigned(4649, LUT_AMPL_WIDTH - 1),
		31284 => to_unsigned(4646, LUT_AMPL_WIDTH - 1),
		31285 => to_unsigned(4643, LUT_AMPL_WIDTH - 1),
		31286 => to_unsigned(4640, LUT_AMPL_WIDTH - 1),
		31287 => to_unsigned(4637, LUT_AMPL_WIDTH - 1),
		31288 => to_unsigned(4634, LUT_AMPL_WIDTH - 1),
		31289 => to_unsigned(4631, LUT_AMPL_WIDTH - 1),
		31290 => to_unsigned(4628, LUT_AMPL_WIDTH - 1),
		31291 => to_unsigned(4624, LUT_AMPL_WIDTH - 1),
		31292 => to_unsigned(4621, LUT_AMPL_WIDTH - 1),
		31293 => to_unsigned(4618, LUT_AMPL_WIDTH - 1),
		31294 => to_unsigned(4615, LUT_AMPL_WIDTH - 1),
		31295 => to_unsigned(4612, LUT_AMPL_WIDTH - 1),
		31296 => to_unsigned(4609, LUT_AMPL_WIDTH - 1),
		31297 => to_unsigned(4606, LUT_AMPL_WIDTH - 1),
		31298 => to_unsigned(4603, LUT_AMPL_WIDTH - 1),
		31299 => to_unsigned(4600, LUT_AMPL_WIDTH - 1),
		31300 => to_unsigned(4597, LUT_AMPL_WIDTH - 1),
		31301 => to_unsigned(4593, LUT_AMPL_WIDTH - 1),
		31302 => to_unsigned(4590, LUT_AMPL_WIDTH - 1),
		31303 => to_unsigned(4587, LUT_AMPL_WIDTH - 1),
		31304 => to_unsigned(4584, LUT_AMPL_WIDTH - 1),
		31305 => to_unsigned(4581, LUT_AMPL_WIDTH - 1),
		31306 => to_unsigned(4578, LUT_AMPL_WIDTH - 1),
		31307 => to_unsigned(4575, LUT_AMPL_WIDTH - 1),
		31308 => to_unsigned(4572, LUT_AMPL_WIDTH - 1),
		31309 => to_unsigned(4569, LUT_AMPL_WIDTH - 1),
		31310 => to_unsigned(4565, LUT_AMPL_WIDTH - 1),
		31311 => to_unsigned(4562, LUT_AMPL_WIDTH - 1),
		31312 => to_unsigned(4559, LUT_AMPL_WIDTH - 1),
		31313 => to_unsigned(4556, LUT_AMPL_WIDTH - 1),
		31314 => to_unsigned(4553, LUT_AMPL_WIDTH - 1),
		31315 => to_unsigned(4550, LUT_AMPL_WIDTH - 1),
		31316 => to_unsigned(4547, LUT_AMPL_WIDTH - 1),
		31317 => to_unsigned(4544, LUT_AMPL_WIDTH - 1),
		31318 => to_unsigned(4541, LUT_AMPL_WIDTH - 1),
		31319 => to_unsigned(4537, LUT_AMPL_WIDTH - 1),
		31320 => to_unsigned(4534, LUT_AMPL_WIDTH - 1),
		31321 => to_unsigned(4531, LUT_AMPL_WIDTH - 1),
		31322 => to_unsigned(4528, LUT_AMPL_WIDTH - 1),
		31323 => to_unsigned(4525, LUT_AMPL_WIDTH - 1),
		31324 => to_unsigned(4522, LUT_AMPL_WIDTH - 1),
		31325 => to_unsigned(4519, LUT_AMPL_WIDTH - 1),
		31326 => to_unsigned(4516, LUT_AMPL_WIDTH - 1),
		31327 => to_unsigned(4513, LUT_AMPL_WIDTH - 1),
		31328 => to_unsigned(4509, LUT_AMPL_WIDTH - 1),
		31329 => to_unsigned(4506, LUT_AMPL_WIDTH - 1),
		31330 => to_unsigned(4503, LUT_AMPL_WIDTH - 1),
		31331 => to_unsigned(4500, LUT_AMPL_WIDTH - 1),
		31332 => to_unsigned(4497, LUT_AMPL_WIDTH - 1),
		31333 => to_unsigned(4494, LUT_AMPL_WIDTH - 1),
		31334 => to_unsigned(4491, LUT_AMPL_WIDTH - 1),
		31335 => to_unsigned(4488, LUT_AMPL_WIDTH - 1),
		31336 => to_unsigned(4485, LUT_AMPL_WIDTH - 1),
		31337 => to_unsigned(4481, LUT_AMPL_WIDTH - 1),
		31338 => to_unsigned(4478, LUT_AMPL_WIDTH - 1),
		31339 => to_unsigned(4475, LUT_AMPL_WIDTH - 1),
		31340 => to_unsigned(4472, LUT_AMPL_WIDTH - 1),
		31341 => to_unsigned(4469, LUT_AMPL_WIDTH - 1),
		31342 => to_unsigned(4466, LUT_AMPL_WIDTH - 1),
		31343 => to_unsigned(4463, LUT_AMPL_WIDTH - 1),
		31344 => to_unsigned(4460, LUT_AMPL_WIDTH - 1),
		31345 => to_unsigned(4456, LUT_AMPL_WIDTH - 1),
		31346 => to_unsigned(4453, LUT_AMPL_WIDTH - 1),
		31347 => to_unsigned(4450, LUT_AMPL_WIDTH - 1),
		31348 => to_unsigned(4447, LUT_AMPL_WIDTH - 1),
		31349 => to_unsigned(4444, LUT_AMPL_WIDTH - 1),
		31350 => to_unsigned(4441, LUT_AMPL_WIDTH - 1),
		31351 => to_unsigned(4438, LUT_AMPL_WIDTH - 1),
		31352 => to_unsigned(4435, LUT_AMPL_WIDTH - 1),
		31353 => to_unsigned(4432, LUT_AMPL_WIDTH - 1),
		31354 => to_unsigned(4428, LUT_AMPL_WIDTH - 1),
		31355 => to_unsigned(4425, LUT_AMPL_WIDTH - 1),
		31356 => to_unsigned(4422, LUT_AMPL_WIDTH - 1),
		31357 => to_unsigned(4419, LUT_AMPL_WIDTH - 1),
		31358 => to_unsigned(4416, LUT_AMPL_WIDTH - 1),
		31359 => to_unsigned(4413, LUT_AMPL_WIDTH - 1),
		31360 => to_unsigned(4410, LUT_AMPL_WIDTH - 1),
		31361 => to_unsigned(4407, LUT_AMPL_WIDTH - 1),
		31362 => to_unsigned(4404, LUT_AMPL_WIDTH - 1),
		31363 => to_unsigned(4400, LUT_AMPL_WIDTH - 1),
		31364 => to_unsigned(4397, LUT_AMPL_WIDTH - 1),
		31365 => to_unsigned(4394, LUT_AMPL_WIDTH - 1),
		31366 => to_unsigned(4391, LUT_AMPL_WIDTH - 1),
		31367 => to_unsigned(4388, LUT_AMPL_WIDTH - 1),
		31368 => to_unsigned(4385, LUT_AMPL_WIDTH - 1),
		31369 => to_unsigned(4382, LUT_AMPL_WIDTH - 1),
		31370 => to_unsigned(4379, LUT_AMPL_WIDTH - 1),
		31371 => to_unsigned(4376, LUT_AMPL_WIDTH - 1),
		31372 => to_unsigned(4372, LUT_AMPL_WIDTH - 1),
		31373 => to_unsigned(4369, LUT_AMPL_WIDTH - 1),
		31374 => to_unsigned(4366, LUT_AMPL_WIDTH - 1),
		31375 => to_unsigned(4363, LUT_AMPL_WIDTH - 1),
		31376 => to_unsigned(4360, LUT_AMPL_WIDTH - 1),
		31377 => to_unsigned(4357, LUT_AMPL_WIDTH - 1),
		31378 => to_unsigned(4354, LUT_AMPL_WIDTH - 1),
		31379 => to_unsigned(4351, LUT_AMPL_WIDTH - 1),
		31380 => to_unsigned(4348, LUT_AMPL_WIDTH - 1),
		31381 => to_unsigned(4344, LUT_AMPL_WIDTH - 1),
		31382 => to_unsigned(4341, LUT_AMPL_WIDTH - 1),
		31383 => to_unsigned(4338, LUT_AMPL_WIDTH - 1),
		31384 => to_unsigned(4335, LUT_AMPL_WIDTH - 1),
		31385 => to_unsigned(4332, LUT_AMPL_WIDTH - 1),
		31386 => to_unsigned(4329, LUT_AMPL_WIDTH - 1),
		31387 => to_unsigned(4326, LUT_AMPL_WIDTH - 1),
		31388 => to_unsigned(4323, LUT_AMPL_WIDTH - 1),
		31389 => to_unsigned(4320, LUT_AMPL_WIDTH - 1),
		31390 => to_unsigned(4316, LUT_AMPL_WIDTH - 1),
		31391 => to_unsigned(4313, LUT_AMPL_WIDTH - 1),
		31392 => to_unsigned(4310, LUT_AMPL_WIDTH - 1),
		31393 => to_unsigned(4307, LUT_AMPL_WIDTH - 1),
		31394 => to_unsigned(4304, LUT_AMPL_WIDTH - 1),
		31395 => to_unsigned(4301, LUT_AMPL_WIDTH - 1),
		31396 => to_unsigned(4298, LUT_AMPL_WIDTH - 1),
		31397 => to_unsigned(4295, LUT_AMPL_WIDTH - 1),
		31398 => to_unsigned(4291, LUT_AMPL_WIDTH - 1),
		31399 => to_unsigned(4288, LUT_AMPL_WIDTH - 1),
		31400 => to_unsigned(4285, LUT_AMPL_WIDTH - 1),
		31401 => to_unsigned(4282, LUT_AMPL_WIDTH - 1),
		31402 => to_unsigned(4279, LUT_AMPL_WIDTH - 1),
		31403 => to_unsigned(4276, LUT_AMPL_WIDTH - 1),
		31404 => to_unsigned(4273, LUT_AMPL_WIDTH - 1),
		31405 => to_unsigned(4270, LUT_AMPL_WIDTH - 1),
		31406 => to_unsigned(4267, LUT_AMPL_WIDTH - 1),
		31407 => to_unsigned(4263, LUT_AMPL_WIDTH - 1),
		31408 => to_unsigned(4260, LUT_AMPL_WIDTH - 1),
		31409 => to_unsigned(4257, LUT_AMPL_WIDTH - 1),
		31410 => to_unsigned(4254, LUT_AMPL_WIDTH - 1),
		31411 => to_unsigned(4251, LUT_AMPL_WIDTH - 1),
		31412 => to_unsigned(4248, LUT_AMPL_WIDTH - 1),
		31413 => to_unsigned(4245, LUT_AMPL_WIDTH - 1),
		31414 => to_unsigned(4242, LUT_AMPL_WIDTH - 1),
		31415 => to_unsigned(4239, LUT_AMPL_WIDTH - 1),
		31416 => to_unsigned(4235, LUT_AMPL_WIDTH - 1),
		31417 => to_unsigned(4232, LUT_AMPL_WIDTH - 1),
		31418 => to_unsigned(4229, LUT_AMPL_WIDTH - 1),
		31419 => to_unsigned(4226, LUT_AMPL_WIDTH - 1),
		31420 => to_unsigned(4223, LUT_AMPL_WIDTH - 1),
		31421 => to_unsigned(4220, LUT_AMPL_WIDTH - 1),
		31422 => to_unsigned(4217, LUT_AMPL_WIDTH - 1),
		31423 => to_unsigned(4214, LUT_AMPL_WIDTH - 1),
		31424 => to_unsigned(4210, LUT_AMPL_WIDTH - 1),
		31425 => to_unsigned(4207, LUT_AMPL_WIDTH - 1),
		31426 => to_unsigned(4204, LUT_AMPL_WIDTH - 1),
		31427 => to_unsigned(4201, LUT_AMPL_WIDTH - 1),
		31428 => to_unsigned(4198, LUT_AMPL_WIDTH - 1),
		31429 => to_unsigned(4195, LUT_AMPL_WIDTH - 1),
		31430 => to_unsigned(4192, LUT_AMPL_WIDTH - 1),
		31431 => to_unsigned(4189, LUT_AMPL_WIDTH - 1),
		31432 => to_unsigned(4186, LUT_AMPL_WIDTH - 1),
		31433 => to_unsigned(4182, LUT_AMPL_WIDTH - 1),
		31434 => to_unsigned(4179, LUT_AMPL_WIDTH - 1),
		31435 => to_unsigned(4176, LUT_AMPL_WIDTH - 1),
		31436 => to_unsigned(4173, LUT_AMPL_WIDTH - 1),
		31437 => to_unsigned(4170, LUT_AMPL_WIDTH - 1),
		31438 => to_unsigned(4167, LUT_AMPL_WIDTH - 1),
		31439 => to_unsigned(4164, LUT_AMPL_WIDTH - 1),
		31440 => to_unsigned(4161, LUT_AMPL_WIDTH - 1),
		31441 => to_unsigned(4158, LUT_AMPL_WIDTH - 1),
		31442 => to_unsigned(4154, LUT_AMPL_WIDTH - 1),
		31443 => to_unsigned(4151, LUT_AMPL_WIDTH - 1),
		31444 => to_unsigned(4148, LUT_AMPL_WIDTH - 1),
		31445 => to_unsigned(4145, LUT_AMPL_WIDTH - 1),
		31446 => to_unsigned(4142, LUT_AMPL_WIDTH - 1),
		31447 => to_unsigned(4139, LUT_AMPL_WIDTH - 1),
		31448 => to_unsigned(4136, LUT_AMPL_WIDTH - 1),
		31449 => to_unsigned(4133, LUT_AMPL_WIDTH - 1),
		31450 => to_unsigned(4129, LUT_AMPL_WIDTH - 1),
		31451 => to_unsigned(4126, LUT_AMPL_WIDTH - 1),
		31452 => to_unsigned(4123, LUT_AMPL_WIDTH - 1),
		31453 => to_unsigned(4120, LUT_AMPL_WIDTH - 1),
		31454 => to_unsigned(4117, LUT_AMPL_WIDTH - 1),
		31455 => to_unsigned(4114, LUT_AMPL_WIDTH - 1),
		31456 => to_unsigned(4111, LUT_AMPL_WIDTH - 1),
		31457 => to_unsigned(4108, LUT_AMPL_WIDTH - 1),
		31458 => to_unsigned(4105, LUT_AMPL_WIDTH - 1),
		31459 => to_unsigned(4101, LUT_AMPL_WIDTH - 1),
		31460 => to_unsigned(4098, LUT_AMPL_WIDTH - 1),
		31461 => to_unsigned(4095, LUT_AMPL_WIDTH - 1),
		31462 => to_unsigned(4092, LUT_AMPL_WIDTH - 1),
		31463 => to_unsigned(4089, LUT_AMPL_WIDTH - 1),
		31464 => to_unsigned(4086, LUT_AMPL_WIDTH - 1),
		31465 => to_unsigned(4083, LUT_AMPL_WIDTH - 1),
		31466 => to_unsigned(4080, LUT_AMPL_WIDTH - 1),
		31467 => to_unsigned(4076, LUT_AMPL_WIDTH - 1),
		31468 => to_unsigned(4073, LUT_AMPL_WIDTH - 1),
		31469 => to_unsigned(4070, LUT_AMPL_WIDTH - 1),
		31470 => to_unsigned(4067, LUT_AMPL_WIDTH - 1),
		31471 => to_unsigned(4064, LUT_AMPL_WIDTH - 1),
		31472 => to_unsigned(4061, LUT_AMPL_WIDTH - 1),
		31473 => to_unsigned(4058, LUT_AMPL_WIDTH - 1),
		31474 => to_unsigned(4055, LUT_AMPL_WIDTH - 1),
		31475 => to_unsigned(4052, LUT_AMPL_WIDTH - 1),
		31476 => to_unsigned(4048, LUT_AMPL_WIDTH - 1),
		31477 => to_unsigned(4045, LUT_AMPL_WIDTH - 1),
		31478 => to_unsigned(4042, LUT_AMPL_WIDTH - 1),
		31479 => to_unsigned(4039, LUT_AMPL_WIDTH - 1),
		31480 => to_unsigned(4036, LUT_AMPL_WIDTH - 1),
		31481 => to_unsigned(4033, LUT_AMPL_WIDTH - 1),
		31482 => to_unsigned(4030, LUT_AMPL_WIDTH - 1),
		31483 => to_unsigned(4027, LUT_AMPL_WIDTH - 1),
		31484 => to_unsigned(4024, LUT_AMPL_WIDTH - 1),
		31485 => to_unsigned(4020, LUT_AMPL_WIDTH - 1),
		31486 => to_unsigned(4017, LUT_AMPL_WIDTH - 1),
		31487 => to_unsigned(4014, LUT_AMPL_WIDTH - 1),
		31488 => to_unsigned(4011, LUT_AMPL_WIDTH - 1),
		31489 => to_unsigned(4008, LUT_AMPL_WIDTH - 1),
		31490 => to_unsigned(4005, LUT_AMPL_WIDTH - 1),
		31491 => to_unsigned(4002, LUT_AMPL_WIDTH - 1),
		31492 => to_unsigned(3999, LUT_AMPL_WIDTH - 1),
		31493 => to_unsigned(3995, LUT_AMPL_WIDTH - 1),
		31494 => to_unsigned(3992, LUT_AMPL_WIDTH - 1),
		31495 => to_unsigned(3989, LUT_AMPL_WIDTH - 1),
		31496 => to_unsigned(3986, LUT_AMPL_WIDTH - 1),
		31497 => to_unsigned(3983, LUT_AMPL_WIDTH - 1),
		31498 => to_unsigned(3980, LUT_AMPL_WIDTH - 1),
		31499 => to_unsigned(3977, LUT_AMPL_WIDTH - 1),
		31500 => to_unsigned(3974, LUT_AMPL_WIDTH - 1),
		31501 => to_unsigned(3970, LUT_AMPL_WIDTH - 1),
		31502 => to_unsigned(3967, LUT_AMPL_WIDTH - 1),
		31503 => to_unsigned(3964, LUT_AMPL_WIDTH - 1),
		31504 => to_unsigned(3961, LUT_AMPL_WIDTH - 1),
		31505 => to_unsigned(3958, LUT_AMPL_WIDTH - 1),
		31506 => to_unsigned(3955, LUT_AMPL_WIDTH - 1),
		31507 => to_unsigned(3952, LUT_AMPL_WIDTH - 1),
		31508 => to_unsigned(3949, LUT_AMPL_WIDTH - 1),
		31509 => to_unsigned(3946, LUT_AMPL_WIDTH - 1),
		31510 => to_unsigned(3942, LUT_AMPL_WIDTH - 1),
		31511 => to_unsigned(3939, LUT_AMPL_WIDTH - 1),
		31512 => to_unsigned(3936, LUT_AMPL_WIDTH - 1),
		31513 => to_unsigned(3933, LUT_AMPL_WIDTH - 1),
		31514 => to_unsigned(3930, LUT_AMPL_WIDTH - 1),
		31515 => to_unsigned(3927, LUT_AMPL_WIDTH - 1),
		31516 => to_unsigned(3924, LUT_AMPL_WIDTH - 1),
		31517 => to_unsigned(3921, LUT_AMPL_WIDTH - 1),
		31518 => to_unsigned(3917, LUT_AMPL_WIDTH - 1),
		31519 => to_unsigned(3914, LUT_AMPL_WIDTH - 1),
		31520 => to_unsigned(3911, LUT_AMPL_WIDTH - 1),
		31521 => to_unsigned(3908, LUT_AMPL_WIDTH - 1),
		31522 => to_unsigned(3905, LUT_AMPL_WIDTH - 1),
		31523 => to_unsigned(3902, LUT_AMPL_WIDTH - 1),
		31524 => to_unsigned(3899, LUT_AMPL_WIDTH - 1),
		31525 => to_unsigned(3896, LUT_AMPL_WIDTH - 1),
		31526 => to_unsigned(3893, LUT_AMPL_WIDTH - 1),
		31527 => to_unsigned(3889, LUT_AMPL_WIDTH - 1),
		31528 => to_unsigned(3886, LUT_AMPL_WIDTH - 1),
		31529 => to_unsigned(3883, LUT_AMPL_WIDTH - 1),
		31530 => to_unsigned(3880, LUT_AMPL_WIDTH - 1),
		31531 => to_unsigned(3877, LUT_AMPL_WIDTH - 1),
		31532 => to_unsigned(3874, LUT_AMPL_WIDTH - 1),
		31533 => to_unsigned(3871, LUT_AMPL_WIDTH - 1),
		31534 => to_unsigned(3868, LUT_AMPL_WIDTH - 1),
		31535 => to_unsigned(3864, LUT_AMPL_WIDTH - 1),
		31536 => to_unsigned(3861, LUT_AMPL_WIDTH - 1),
		31537 => to_unsigned(3858, LUT_AMPL_WIDTH - 1),
		31538 => to_unsigned(3855, LUT_AMPL_WIDTH - 1),
		31539 => to_unsigned(3852, LUT_AMPL_WIDTH - 1),
		31540 => to_unsigned(3849, LUT_AMPL_WIDTH - 1),
		31541 => to_unsigned(3846, LUT_AMPL_WIDTH - 1),
		31542 => to_unsigned(3843, LUT_AMPL_WIDTH - 1),
		31543 => to_unsigned(3839, LUT_AMPL_WIDTH - 1),
		31544 => to_unsigned(3836, LUT_AMPL_WIDTH - 1),
		31545 => to_unsigned(3833, LUT_AMPL_WIDTH - 1),
		31546 => to_unsigned(3830, LUT_AMPL_WIDTH - 1),
		31547 => to_unsigned(3827, LUT_AMPL_WIDTH - 1),
		31548 => to_unsigned(3824, LUT_AMPL_WIDTH - 1),
		31549 => to_unsigned(3821, LUT_AMPL_WIDTH - 1),
		31550 => to_unsigned(3818, LUT_AMPL_WIDTH - 1),
		31551 => to_unsigned(3815, LUT_AMPL_WIDTH - 1),
		31552 => to_unsigned(3811, LUT_AMPL_WIDTH - 1),
		31553 => to_unsigned(3808, LUT_AMPL_WIDTH - 1),
		31554 => to_unsigned(3805, LUT_AMPL_WIDTH - 1),
		31555 => to_unsigned(3802, LUT_AMPL_WIDTH - 1),
		31556 => to_unsigned(3799, LUT_AMPL_WIDTH - 1),
		31557 => to_unsigned(3796, LUT_AMPL_WIDTH - 1),
		31558 => to_unsigned(3793, LUT_AMPL_WIDTH - 1),
		31559 => to_unsigned(3790, LUT_AMPL_WIDTH - 1),
		31560 => to_unsigned(3786, LUT_AMPL_WIDTH - 1),
		31561 => to_unsigned(3783, LUT_AMPL_WIDTH - 1),
		31562 => to_unsigned(3780, LUT_AMPL_WIDTH - 1),
		31563 => to_unsigned(3777, LUT_AMPL_WIDTH - 1),
		31564 => to_unsigned(3774, LUT_AMPL_WIDTH - 1),
		31565 => to_unsigned(3771, LUT_AMPL_WIDTH - 1),
		31566 => to_unsigned(3768, LUT_AMPL_WIDTH - 1),
		31567 => to_unsigned(3765, LUT_AMPL_WIDTH - 1),
		31568 => to_unsigned(3761, LUT_AMPL_WIDTH - 1),
		31569 => to_unsigned(3758, LUT_AMPL_WIDTH - 1),
		31570 => to_unsigned(3755, LUT_AMPL_WIDTH - 1),
		31571 => to_unsigned(3752, LUT_AMPL_WIDTH - 1),
		31572 => to_unsigned(3749, LUT_AMPL_WIDTH - 1),
		31573 => to_unsigned(3746, LUT_AMPL_WIDTH - 1),
		31574 => to_unsigned(3743, LUT_AMPL_WIDTH - 1),
		31575 => to_unsigned(3740, LUT_AMPL_WIDTH - 1),
		31576 => to_unsigned(3737, LUT_AMPL_WIDTH - 1),
		31577 => to_unsigned(3733, LUT_AMPL_WIDTH - 1),
		31578 => to_unsigned(3730, LUT_AMPL_WIDTH - 1),
		31579 => to_unsigned(3727, LUT_AMPL_WIDTH - 1),
		31580 => to_unsigned(3724, LUT_AMPL_WIDTH - 1),
		31581 => to_unsigned(3721, LUT_AMPL_WIDTH - 1),
		31582 => to_unsigned(3718, LUT_AMPL_WIDTH - 1),
		31583 => to_unsigned(3715, LUT_AMPL_WIDTH - 1),
		31584 => to_unsigned(3712, LUT_AMPL_WIDTH - 1),
		31585 => to_unsigned(3708, LUT_AMPL_WIDTH - 1),
		31586 => to_unsigned(3705, LUT_AMPL_WIDTH - 1),
		31587 => to_unsigned(3702, LUT_AMPL_WIDTH - 1),
		31588 => to_unsigned(3699, LUT_AMPL_WIDTH - 1),
		31589 => to_unsigned(3696, LUT_AMPL_WIDTH - 1),
		31590 => to_unsigned(3693, LUT_AMPL_WIDTH - 1),
		31591 => to_unsigned(3690, LUT_AMPL_WIDTH - 1),
		31592 => to_unsigned(3687, LUT_AMPL_WIDTH - 1),
		31593 => to_unsigned(3683, LUT_AMPL_WIDTH - 1),
		31594 => to_unsigned(3680, LUT_AMPL_WIDTH - 1),
		31595 => to_unsigned(3677, LUT_AMPL_WIDTH - 1),
		31596 => to_unsigned(3674, LUT_AMPL_WIDTH - 1),
		31597 => to_unsigned(3671, LUT_AMPL_WIDTH - 1),
		31598 => to_unsigned(3668, LUT_AMPL_WIDTH - 1),
		31599 => to_unsigned(3665, LUT_AMPL_WIDTH - 1),
		31600 => to_unsigned(3662, LUT_AMPL_WIDTH - 1),
		31601 => to_unsigned(3658, LUT_AMPL_WIDTH - 1),
		31602 => to_unsigned(3655, LUT_AMPL_WIDTH - 1),
		31603 => to_unsigned(3652, LUT_AMPL_WIDTH - 1),
		31604 => to_unsigned(3649, LUT_AMPL_WIDTH - 1),
		31605 => to_unsigned(3646, LUT_AMPL_WIDTH - 1),
		31606 => to_unsigned(3643, LUT_AMPL_WIDTH - 1),
		31607 => to_unsigned(3640, LUT_AMPL_WIDTH - 1),
		31608 => to_unsigned(3637, LUT_AMPL_WIDTH - 1),
		31609 => to_unsigned(3634, LUT_AMPL_WIDTH - 1),
		31610 => to_unsigned(3630, LUT_AMPL_WIDTH - 1),
		31611 => to_unsigned(3627, LUT_AMPL_WIDTH - 1),
		31612 => to_unsigned(3624, LUT_AMPL_WIDTH - 1),
		31613 => to_unsigned(3621, LUT_AMPL_WIDTH - 1),
		31614 => to_unsigned(3618, LUT_AMPL_WIDTH - 1),
		31615 => to_unsigned(3615, LUT_AMPL_WIDTH - 1),
		31616 => to_unsigned(3612, LUT_AMPL_WIDTH - 1),
		31617 => to_unsigned(3609, LUT_AMPL_WIDTH - 1),
		31618 => to_unsigned(3605, LUT_AMPL_WIDTH - 1),
		31619 => to_unsigned(3602, LUT_AMPL_WIDTH - 1),
		31620 => to_unsigned(3599, LUT_AMPL_WIDTH - 1),
		31621 => to_unsigned(3596, LUT_AMPL_WIDTH - 1),
		31622 => to_unsigned(3593, LUT_AMPL_WIDTH - 1),
		31623 => to_unsigned(3590, LUT_AMPL_WIDTH - 1),
		31624 => to_unsigned(3587, LUT_AMPL_WIDTH - 1),
		31625 => to_unsigned(3584, LUT_AMPL_WIDTH - 1),
		31626 => to_unsigned(3580, LUT_AMPL_WIDTH - 1),
		31627 => to_unsigned(3577, LUT_AMPL_WIDTH - 1),
		31628 => to_unsigned(3574, LUT_AMPL_WIDTH - 1),
		31629 => to_unsigned(3571, LUT_AMPL_WIDTH - 1),
		31630 => to_unsigned(3568, LUT_AMPL_WIDTH - 1),
		31631 => to_unsigned(3565, LUT_AMPL_WIDTH - 1),
		31632 => to_unsigned(3562, LUT_AMPL_WIDTH - 1),
		31633 => to_unsigned(3559, LUT_AMPL_WIDTH - 1),
		31634 => to_unsigned(3555, LUT_AMPL_WIDTH - 1),
		31635 => to_unsigned(3552, LUT_AMPL_WIDTH - 1),
		31636 => to_unsigned(3549, LUT_AMPL_WIDTH - 1),
		31637 => to_unsigned(3546, LUT_AMPL_WIDTH - 1),
		31638 => to_unsigned(3543, LUT_AMPL_WIDTH - 1),
		31639 => to_unsigned(3540, LUT_AMPL_WIDTH - 1),
		31640 => to_unsigned(3537, LUT_AMPL_WIDTH - 1),
		31641 => to_unsigned(3534, LUT_AMPL_WIDTH - 1),
		31642 => to_unsigned(3530, LUT_AMPL_WIDTH - 1),
		31643 => to_unsigned(3527, LUT_AMPL_WIDTH - 1),
		31644 => to_unsigned(3524, LUT_AMPL_WIDTH - 1),
		31645 => to_unsigned(3521, LUT_AMPL_WIDTH - 1),
		31646 => to_unsigned(3518, LUT_AMPL_WIDTH - 1),
		31647 => to_unsigned(3515, LUT_AMPL_WIDTH - 1),
		31648 => to_unsigned(3512, LUT_AMPL_WIDTH - 1),
		31649 => to_unsigned(3509, LUT_AMPL_WIDTH - 1),
		31650 => to_unsigned(3505, LUT_AMPL_WIDTH - 1),
		31651 => to_unsigned(3502, LUT_AMPL_WIDTH - 1),
		31652 => to_unsigned(3499, LUT_AMPL_WIDTH - 1),
		31653 => to_unsigned(3496, LUT_AMPL_WIDTH - 1),
		31654 => to_unsigned(3493, LUT_AMPL_WIDTH - 1),
		31655 => to_unsigned(3490, LUT_AMPL_WIDTH - 1),
		31656 => to_unsigned(3487, LUT_AMPL_WIDTH - 1),
		31657 => to_unsigned(3484, LUT_AMPL_WIDTH - 1),
		31658 => to_unsigned(3480, LUT_AMPL_WIDTH - 1),
		31659 => to_unsigned(3477, LUT_AMPL_WIDTH - 1),
		31660 => to_unsigned(3474, LUT_AMPL_WIDTH - 1),
		31661 => to_unsigned(3471, LUT_AMPL_WIDTH - 1),
		31662 => to_unsigned(3468, LUT_AMPL_WIDTH - 1),
		31663 => to_unsigned(3465, LUT_AMPL_WIDTH - 1),
		31664 => to_unsigned(3462, LUT_AMPL_WIDTH - 1),
		31665 => to_unsigned(3459, LUT_AMPL_WIDTH - 1),
		31666 => to_unsigned(3455, LUT_AMPL_WIDTH - 1),
		31667 => to_unsigned(3452, LUT_AMPL_WIDTH - 1),
		31668 => to_unsigned(3449, LUT_AMPL_WIDTH - 1),
		31669 => to_unsigned(3446, LUT_AMPL_WIDTH - 1),
		31670 => to_unsigned(3443, LUT_AMPL_WIDTH - 1),
		31671 => to_unsigned(3440, LUT_AMPL_WIDTH - 1),
		31672 => to_unsigned(3437, LUT_AMPL_WIDTH - 1),
		31673 => to_unsigned(3434, LUT_AMPL_WIDTH - 1),
		31674 => to_unsigned(3430, LUT_AMPL_WIDTH - 1),
		31675 => to_unsigned(3427, LUT_AMPL_WIDTH - 1),
		31676 => to_unsigned(3424, LUT_AMPL_WIDTH - 1),
		31677 => to_unsigned(3421, LUT_AMPL_WIDTH - 1),
		31678 => to_unsigned(3418, LUT_AMPL_WIDTH - 1),
		31679 => to_unsigned(3415, LUT_AMPL_WIDTH - 1),
		31680 => to_unsigned(3412, LUT_AMPL_WIDTH - 1),
		31681 => to_unsigned(3409, LUT_AMPL_WIDTH - 1),
		31682 => to_unsigned(3406, LUT_AMPL_WIDTH - 1),
		31683 => to_unsigned(3402, LUT_AMPL_WIDTH - 1),
		31684 => to_unsigned(3399, LUT_AMPL_WIDTH - 1),
		31685 => to_unsigned(3396, LUT_AMPL_WIDTH - 1),
		31686 => to_unsigned(3393, LUT_AMPL_WIDTH - 1),
		31687 => to_unsigned(3390, LUT_AMPL_WIDTH - 1),
		31688 => to_unsigned(3387, LUT_AMPL_WIDTH - 1),
		31689 => to_unsigned(3384, LUT_AMPL_WIDTH - 1),
		31690 => to_unsigned(3381, LUT_AMPL_WIDTH - 1),
		31691 => to_unsigned(3377, LUT_AMPL_WIDTH - 1),
		31692 => to_unsigned(3374, LUT_AMPL_WIDTH - 1),
		31693 => to_unsigned(3371, LUT_AMPL_WIDTH - 1),
		31694 => to_unsigned(3368, LUT_AMPL_WIDTH - 1),
		31695 => to_unsigned(3365, LUT_AMPL_WIDTH - 1),
		31696 => to_unsigned(3362, LUT_AMPL_WIDTH - 1),
		31697 => to_unsigned(3359, LUT_AMPL_WIDTH - 1),
		31698 => to_unsigned(3356, LUT_AMPL_WIDTH - 1),
		31699 => to_unsigned(3352, LUT_AMPL_WIDTH - 1),
		31700 => to_unsigned(3349, LUT_AMPL_WIDTH - 1),
		31701 => to_unsigned(3346, LUT_AMPL_WIDTH - 1),
		31702 => to_unsigned(3343, LUT_AMPL_WIDTH - 1),
		31703 => to_unsigned(3340, LUT_AMPL_WIDTH - 1),
		31704 => to_unsigned(3337, LUT_AMPL_WIDTH - 1),
		31705 => to_unsigned(3334, LUT_AMPL_WIDTH - 1),
		31706 => to_unsigned(3331, LUT_AMPL_WIDTH - 1),
		31707 => to_unsigned(3327, LUT_AMPL_WIDTH - 1),
		31708 => to_unsigned(3324, LUT_AMPL_WIDTH - 1),
		31709 => to_unsigned(3321, LUT_AMPL_WIDTH - 1),
		31710 => to_unsigned(3318, LUT_AMPL_WIDTH - 1),
		31711 => to_unsigned(3315, LUT_AMPL_WIDTH - 1),
		31712 => to_unsigned(3312, LUT_AMPL_WIDTH - 1),
		31713 => to_unsigned(3309, LUT_AMPL_WIDTH - 1),
		31714 => to_unsigned(3306, LUT_AMPL_WIDTH - 1),
		31715 => to_unsigned(3302, LUT_AMPL_WIDTH - 1),
		31716 => to_unsigned(3299, LUT_AMPL_WIDTH - 1),
		31717 => to_unsigned(3296, LUT_AMPL_WIDTH - 1),
		31718 => to_unsigned(3293, LUT_AMPL_WIDTH - 1),
		31719 => to_unsigned(3290, LUT_AMPL_WIDTH - 1),
		31720 => to_unsigned(3287, LUT_AMPL_WIDTH - 1),
		31721 => to_unsigned(3284, LUT_AMPL_WIDTH - 1),
		31722 => to_unsigned(3281, LUT_AMPL_WIDTH - 1),
		31723 => to_unsigned(3277, LUT_AMPL_WIDTH - 1),
		31724 => to_unsigned(3274, LUT_AMPL_WIDTH - 1),
		31725 => to_unsigned(3271, LUT_AMPL_WIDTH - 1),
		31726 => to_unsigned(3268, LUT_AMPL_WIDTH - 1),
		31727 => to_unsigned(3265, LUT_AMPL_WIDTH - 1),
		31728 => to_unsigned(3262, LUT_AMPL_WIDTH - 1),
		31729 => to_unsigned(3259, LUT_AMPL_WIDTH - 1),
		31730 => to_unsigned(3255, LUT_AMPL_WIDTH - 1),
		31731 => to_unsigned(3252, LUT_AMPL_WIDTH - 1),
		31732 => to_unsigned(3249, LUT_AMPL_WIDTH - 1),
		31733 => to_unsigned(3246, LUT_AMPL_WIDTH - 1),
		31734 => to_unsigned(3243, LUT_AMPL_WIDTH - 1),
		31735 => to_unsigned(3240, LUT_AMPL_WIDTH - 1),
		31736 => to_unsigned(3237, LUT_AMPL_WIDTH - 1),
		31737 => to_unsigned(3234, LUT_AMPL_WIDTH - 1),
		31738 => to_unsigned(3230, LUT_AMPL_WIDTH - 1),
		31739 => to_unsigned(3227, LUT_AMPL_WIDTH - 1),
		31740 => to_unsigned(3224, LUT_AMPL_WIDTH - 1),
		31741 => to_unsigned(3221, LUT_AMPL_WIDTH - 1),
		31742 => to_unsigned(3218, LUT_AMPL_WIDTH - 1),
		31743 => to_unsigned(3215, LUT_AMPL_WIDTH - 1),
		31744 => to_unsigned(3212, LUT_AMPL_WIDTH - 1),
		31745 => to_unsigned(3209, LUT_AMPL_WIDTH - 1),
		31746 => to_unsigned(3205, LUT_AMPL_WIDTH - 1),
		31747 => to_unsigned(3202, LUT_AMPL_WIDTH - 1),
		31748 => to_unsigned(3199, LUT_AMPL_WIDTH - 1),
		31749 => to_unsigned(3196, LUT_AMPL_WIDTH - 1),
		31750 => to_unsigned(3193, LUT_AMPL_WIDTH - 1),
		31751 => to_unsigned(3190, LUT_AMPL_WIDTH - 1),
		31752 => to_unsigned(3187, LUT_AMPL_WIDTH - 1),
		31753 => to_unsigned(3184, LUT_AMPL_WIDTH - 1),
		31754 => to_unsigned(3180, LUT_AMPL_WIDTH - 1),
		31755 => to_unsigned(3177, LUT_AMPL_WIDTH - 1),
		31756 => to_unsigned(3174, LUT_AMPL_WIDTH - 1),
		31757 => to_unsigned(3171, LUT_AMPL_WIDTH - 1),
		31758 => to_unsigned(3168, LUT_AMPL_WIDTH - 1),
		31759 => to_unsigned(3165, LUT_AMPL_WIDTH - 1),
		31760 => to_unsigned(3162, LUT_AMPL_WIDTH - 1),
		31761 => to_unsigned(3159, LUT_AMPL_WIDTH - 1),
		31762 => to_unsigned(3155, LUT_AMPL_WIDTH - 1),
		31763 => to_unsigned(3152, LUT_AMPL_WIDTH - 1),
		31764 => to_unsigned(3149, LUT_AMPL_WIDTH - 1),
		31765 => to_unsigned(3146, LUT_AMPL_WIDTH - 1),
		31766 => to_unsigned(3143, LUT_AMPL_WIDTH - 1),
		31767 => to_unsigned(3140, LUT_AMPL_WIDTH - 1),
		31768 => to_unsigned(3137, LUT_AMPL_WIDTH - 1),
		31769 => to_unsigned(3134, LUT_AMPL_WIDTH - 1),
		31770 => to_unsigned(3130, LUT_AMPL_WIDTH - 1),
		31771 => to_unsigned(3127, LUT_AMPL_WIDTH - 1),
		31772 => to_unsigned(3124, LUT_AMPL_WIDTH - 1),
		31773 => to_unsigned(3121, LUT_AMPL_WIDTH - 1),
		31774 => to_unsigned(3118, LUT_AMPL_WIDTH - 1),
		31775 => to_unsigned(3115, LUT_AMPL_WIDTH - 1),
		31776 => to_unsigned(3112, LUT_AMPL_WIDTH - 1),
		31777 => to_unsigned(3109, LUT_AMPL_WIDTH - 1),
		31778 => to_unsigned(3105, LUT_AMPL_WIDTH - 1),
		31779 => to_unsigned(3102, LUT_AMPL_WIDTH - 1),
		31780 => to_unsigned(3099, LUT_AMPL_WIDTH - 1),
		31781 => to_unsigned(3096, LUT_AMPL_WIDTH - 1),
		31782 => to_unsigned(3093, LUT_AMPL_WIDTH - 1),
		31783 => to_unsigned(3090, LUT_AMPL_WIDTH - 1),
		31784 => to_unsigned(3087, LUT_AMPL_WIDTH - 1),
		31785 => to_unsigned(3084, LUT_AMPL_WIDTH - 1),
		31786 => to_unsigned(3080, LUT_AMPL_WIDTH - 1),
		31787 => to_unsigned(3077, LUT_AMPL_WIDTH - 1),
		31788 => to_unsigned(3074, LUT_AMPL_WIDTH - 1),
		31789 => to_unsigned(3071, LUT_AMPL_WIDTH - 1),
		31790 => to_unsigned(3068, LUT_AMPL_WIDTH - 1),
		31791 => to_unsigned(3065, LUT_AMPL_WIDTH - 1),
		31792 => to_unsigned(3062, LUT_AMPL_WIDTH - 1),
		31793 => to_unsigned(3059, LUT_AMPL_WIDTH - 1),
		31794 => to_unsigned(3055, LUT_AMPL_WIDTH - 1),
		31795 => to_unsigned(3052, LUT_AMPL_WIDTH - 1),
		31796 => to_unsigned(3049, LUT_AMPL_WIDTH - 1),
		31797 => to_unsigned(3046, LUT_AMPL_WIDTH - 1),
		31798 => to_unsigned(3043, LUT_AMPL_WIDTH - 1),
		31799 => to_unsigned(3040, LUT_AMPL_WIDTH - 1),
		31800 => to_unsigned(3037, LUT_AMPL_WIDTH - 1),
		31801 => to_unsigned(3033, LUT_AMPL_WIDTH - 1),
		31802 => to_unsigned(3030, LUT_AMPL_WIDTH - 1),
		31803 => to_unsigned(3027, LUT_AMPL_WIDTH - 1),
		31804 => to_unsigned(3024, LUT_AMPL_WIDTH - 1),
		31805 => to_unsigned(3021, LUT_AMPL_WIDTH - 1),
		31806 => to_unsigned(3018, LUT_AMPL_WIDTH - 1),
		31807 => to_unsigned(3015, LUT_AMPL_WIDTH - 1),
		31808 => to_unsigned(3012, LUT_AMPL_WIDTH - 1),
		31809 => to_unsigned(3008, LUT_AMPL_WIDTH - 1),
		31810 => to_unsigned(3005, LUT_AMPL_WIDTH - 1),
		31811 => to_unsigned(3002, LUT_AMPL_WIDTH - 1),
		31812 => to_unsigned(2999, LUT_AMPL_WIDTH - 1),
		31813 => to_unsigned(2996, LUT_AMPL_WIDTH - 1),
		31814 => to_unsigned(2993, LUT_AMPL_WIDTH - 1),
		31815 => to_unsigned(2990, LUT_AMPL_WIDTH - 1),
		31816 => to_unsigned(2987, LUT_AMPL_WIDTH - 1),
		31817 => to_unsigned(2983, LUT_AMPL_WIDTH - 1),
		31818 => to_unsigned(2980, LUT_AMPL_WIDTH - 1),
		31819 => to_unsigned(2977, LUT_AMPL_WIDTH - 1),
		31820 => to_unsigned(2974, LUT_AMPL_WIDTH - 1),
		31821 => to_unsigned(2971, LUT_AMPL_WIDTH - 1),
		31822 => to_unsigned(2968, LUT_AMPL_WIDTH - 1),
		31823 => to_unsigned(2965, LUT_AMPL_WIDTH - 1),
		31824 => to_unsigned(2962, LUT_AMPL_WIDTH - 1),
		31825 => to_unsigned(2958, LUT_AMPL_WIDTH - 1),
		31826 => to_unsigned(2955, LUT_AMPL_WIDTH - 1),
		31827 => to_unsigned(2952, LUT_AMPL_WIDTH - 1),
		31828 => to_unsigned(2949, LUT_AMPL_WIDTH - 1),
		31829 => to_unsigned(2946, LUT_AMPL_WIDTH - 1),
		31830 => to_unsigned(2943, LUT_AMPL_WIDTH - 1),
		31831 => to_unsigned(2940, LUT_AMPL_WIDTH - 1),
		31832 => to_unsigned(2936, LUT_AMPL_WIDTH - 1),
		31833 => to_unsigned(2933, LUT_AMPL_WIDTH - 1),
		31834 => to_unsigned(2930, LUT_AMPL_WIDTH - 1),
		31835 => to_unsigned(2927, LUT_AMPL_WIDTH - 1),
		31836 => to_unsigned(2924, LUT_AMPL_WIDTH - 1),
		31837 => to_unsigned(2921, LUT_AMPL_WIDTH - 1),
		31838 => to_unsigned(2918, LUT_AMPL_WIDTH - 1),
		31839 => to_unsigned(2915, LUT_AMPL_WIDTH - 1),
		31840 => to_unsigned(2911, LUT_AMPL_WIDTH - 1),
		31841 => to_unsigned(2908, LUT_AMPL_WIDTH - 1),
		31842 => to_unsigned(2905, LUT_AMPL_WIDTH - 1),
		31843 => to_unsigned(2902, LUT_AMPL_WIDTH - 1),
		31844 => to_unsigned(2899, LUT_AMPL_WIDTH - 1),
		31845 => to_unsigned(2896, LUT_AMPL_WIDTH - 1),
		31846 => to_unsigned(2893, LUT_AMPL_WIDTH - 1),
		31847 => to_unsigned(2890, LUT_AMPL_WIDTH - 1),
		31848 => to_unsigned(2886, LUT_AMPL_WIDTH - 1),
		31849 => to_unsigned(2883, LUT_AMPL_WIDTH - 1),
		31850 => to_unsigned(2880, LUT_AMPL_WIDTH - 1),
		31851 => to_unsigned(2877, LUT_AMPL_WIDTH - 1),
		31852 => to_unsigned(2874, LUT_AMPL_WIDTH - 1),
		31853 => to_unsigned(2871, LUT_AMPL_WIDTH - 1),
		31854 => to_unsigned(2868, LUT_AMPL_WIDTH - 1),
		31855 => to_unsigned(2865, LUT_AMPL_WIDTH - 1),
		31856 => to_unsigned(2861, LUT_AMPL_WIDTH - 1),
		31857 => to_unsigned(2858, LUT_AMPL_WIDTH - 1),
		31858 => to_unsigned(2855, LUT_AMPL_WIDTH - 1),
		31859 => to_unsigned(2852, LUT_AMPL_WIDTH - 1),
		31860 => to_unsigned(2849, LUT_AMPL_WIDTH - 1),
		31861 => to_unsigned(2846, LUT_AMPL_WIDTH - 1),
		31862 => to_unsigned(2843, LUT_AMPL_WIDTH - 1),
		31863 => to_unsigned(2839, LUT_AMPL_WIDTH - 1),
		31864 => to_unsigned(2836, LUT_AMPL_WIDTH - 1),
		31865 => to_unsigned(2833, LUT_AMPL_WIDTH - 1),
		31866 => to_unsigned(2830, LUT_AMPL_WIDTH - 1),
		31867 => to_unsigned(2827, LUT_AMPL_WIDTH - 1),
		31868 => to_unsigned(2824, LUT_AMPL_WIDTH - 1),
		31869 => to_unsigned(2821, LUT_AMPL_WIDTH - 1),
		31870 => to_unsigned(2818, LUT_AMPL_WIDTH - 1),
		31871 => to_unsigned(2814, LUT_AMPL_WIDTH - 1),
		31872 => to_unsigned(2811, LUT_AMPL_WIDTH - 1),
		31873 => to_unsigned(2808, LUT_AMPL_WIDTH - 1),
		31874 => to_unsigned(2805, LUT_AMPL_WIDTH - 1),
		31875 => to_unsigned(2802, LUT_AMPL_WIDTH - 1),
		31876 => to_unsigned(2799, LUT_AMPL_WIDTH - 1),
		31877 => to_unsigned(2796, LUT_AMPL_WIDTH - 1),
		31878 => to_unsigned(2793, LUT_AMPL_WIDTH - 1),
		31879 => to_unsigned(2789, LUT_AMPL_WIDTH - 1),
		31880 => to_unsigned(2786, LUT_AMPL_WIDTH - 1),
		31881 => to_unsigned(2783, LUT_AMPL_WIDTH - 1),
		31882 => to_unsigned(2780, LUT_AMPL_WIDTH - 1),
		31883 => to_unsigned(2777, LUT_AMPL_WIDTH - 1),
		31884 => to_unsigned(2774, LUT_AMPL_WIDTH - 1),
		31885 => to_unsigned(2771, LUT_AMPL_WIDTH - 1),
		31886 => to_unsigned(2767, LUT_AMPL_WIDTH - 1),
		31887 => to_unsigned(2764, LUT_AMPL_WIDTH - 1),
		31888 => to_unsigned(2761, LUT_AMPL_WIDTH - 1),
		31889 => to_unsigned(2758, LUT_AMPL_WIDTH - 1),
		31890 => to_unsigned(2755, LUT_AMPL_WIDTH - 1),
		31891 => to_unsigned(2752, LUT_AMPL_WIDTH - 1),
		31892 => to_unsigned(2749, LUT_AMPL_WIDTH - 1),
		31893 => to_unsigned(2746, LUT_AMPL_WIDTH - 1),
		31894 => to_unsigned(2742, LUT_AMPL_WIDTH - 1),
		31895 => to_unsigned(2739, LUT_AMPL_WIDTH - 1),
		31896 => to_unsigned(2736, LUT_AMPL_WIDTH - 1),
		31897 => to_unsigned(2733, LUT_AMPL_WIDTH - 1),
		31898 => to_unsigned(2730, LUT_AMPL_WIDTH - 1),
		31899 => to_unsigned(2727, LUT_AMPL_WIDTH - 1),
		31900 => to_unsigned(2724, LUT_AMPL_WIDTH - 1),
		31901 => to_unsigned(2721, LUT_AMPL_WIDTH - 1),
		31902 => to_unsigned(2717, LUT_AMPL_WIDTH - 1),
		31903 => to_unsigned(2714, LUT_AMPL_WIDTH - 1),
		31904 => to_unsigned(2711, LUT_AMPL_WIDTH - 1),
		31905 => to_unsigned(2708, LUT_AMPL_WIDTH - 1),
		31906 => to_unsigned(2705, LUT_AMPL_WIDTH - 1),
		31907 => to_unsigned(2702, LUT_AMPL_WIDTH - 1),
		31908 => to_unsigned(2699, LUT_AMPL_WIDTH - 1),
		31909 => to_unsigned(2695, LUT_AMPL_WIDTH - 1),
		31910 => to_unsigned(2692, LUT_AMPL_WIDTH - 1),
		31911 => to_unsigned(2689, LUT_AMPL_WIDTH - 1),
		31912 => to_unsigned(2686, LUT_AMPL_WIDTH - 1),
		31913 => to_unsigned(2683, LUT_AMPL_WIDTH - 1),
		31914 => to_unsigned(2680, LUT_AMPL_WIDTH - 1),
		31915 => to_unsigned(2677, LUT_AMPL_WIDTH - 1),
		31916 => to_unsigned(2674, LUT_AMPL_WIDTH - 1),
		31917 => to_unsigned(2670, LUT_AMPL_WIDTH - 1),
		31918 => to_unsigned(2667, LUT_AMPL_WIDTH - 1),
		31919 => to_unsigned(2664, LUT_AMPL_WIDTH - 1),
		31920 => to_unsigned(2661, LUT_AMPL_WIDTH - 1),
		31921 => to_unsigned(2658, LUT_AMPL_WIDTH - 1),
		31922 => to_unsigned(2655, LUT_AMPL_WIDTH - 1),
		31923 => to_unsigned(2652, LUT_AMPL_WIDTH - 1),
		31924 => to_unsigned(2649, LUT_AMPL_WIDTH - 1),
		31925 => to_unsigned(2645, LUT_AMPL_WIDTH - 1),
		31926 => to_unsigned(2642, LUT_AMPL_WIDTH - 1),
		31927 => to_unsigned(2639, LUT_AMPL_WIDTH - 1),
		31928 => to_unsigned(2636, LUT_AMPL_WIDTH - 1),
		31929 => to_unsigned(2633, LUT_AMPL_WIDTH - 1),
		31930 => to_unsigned(2630, LUT_AMPL_WIDTH - 1),
		31931 => to_unsigned(2627, LUT_AMPL_WIDTH - 1),
		31932 => to_unsigned(2623, LUT_AMPL_WIDTH - 1),
		31933 => to_unsigned(2620, LUT_AMPL_WIDTH - 1),
		31934 => to_unsigned(2617, LUT_AMPL_WIDTH - 1),
		31935 => to_unsigned(2614, LUT_AMPL_WIDTH - 1),
		31936 => to_unsigned(2611, LUT_AMPL_WIDTH - 1),
		31937 => to_unsigned(2608, LUT_AMPL_WIDTH - 1),
		31938 => to_unsigned(2605, LUT_AMPL_WIDTH - 1),
		31939 => to_unsigned(2602, LUT_AMPL_WIDTH - 1),
		31940 => to_unsigned(2598, LUT_AMPL_WIDTH - 1),
		31941 => to_unsigned(2595, LUT_AMPL_WIDTH - 1),
		31942 => to_unsigned(2592, LUT_AMPL_WIDTH - 1),
		31943 => to_unsigned(2589, LUT_AMPL_WIDTH - 1),
		31944 => to_unsigned(2586, LUT_AMPL_WIDTH - 1),
		31945 => to_unsigned(2583, LUT_AMPL_WIDTH - 1),
		31946 => to_unsigned(2580, LUT_AMPL_WIDTH - 1),
		31947 => to_unsigned(2577, LUT_AMPL_WIDTH - 1),
		31948 => to_unsigned(2573, LUT_AMPL_WIDTH - 1),
		31949 => to_unsigned(2570, LUT_AMPL_WIDTH - 1),
		31950 => to_unsigned(2567, LUT_AMPL_WIDTH - 1),
		31951 => to_unsigned(2564, LUT_AMPL_WIDTH - 1),
		31952 => to_unsigned(2561, LUT_AMPL_WIDTH - 1),
		31953 => to_unsigned(2558, LUT_AMPL_WIDTH - 1),
		31954 => to_unsigned(2555, LUT_AMPL_WIDTH - 1),
		31955 => to_unsigned(2551, LUT_AMPL_WIDTH - 1),
		31956 => to_unsigned(2548, LUT_AMPL_WIDTH - 1),
		31957 => to_unsigned(2545, LUT_AMPL_WIDTH - 1),
		31958 => to_unsigned(2542, LUT_AMPL_WIDTH - 1),
		31959 => to_unsigned(2539, LUT_AMPL_WIDTH - 1),
		31960 => to_unsigned(2536, LUT_AMPL_WIDTH - 1),
		31961 => to_unsigned(2533, LUT_AMPL_WIDTH - 1),
		31962 => to_unsigned(2530, LUT_AMPL_WIDTH - 1),
		31963 => to_unsigned(2526, LUT_AMPL_WIDTH - 1),
		31964 => to_unsigned(2523, LUT_AMPL_WIDTH - 1),
		31965 => to_unsigned(2520, LUT_AMPL_WIDTH - 1),
		31966 => to_unsigned(2517, LUT_AMPL_WIDTH - 1),
		31967 => to_unsigned(2514, LUT_AMPL_WIDTH - 1),
		31968 => to_unsigned(2511, LUT_AMPL_WIDTH - 1),
		31969 => to_unsigned(2508, LUT_AMPL_WIDTH - 1),
		31970 => to_unsigned(2504, LUT_AMPL_WIDTH - 1),
		31971 => to_unsigned(2501, LUT_AMPL_WIDTH - 1),
		31972 => to_unsigned(2498, LUT_AMPL_WIDTH - 1),
		31973 => to_unsigned(2495, LUT_AMPL_WIDTH - 1),
		31974 => to_unsigned(2492, LUT_AMPL_WIDTH - 1),
		31975 => to_unsigned(2489, LUT_AMPL_WIDTH - 1),
		31976 => to_unsigned(2486, LUT_AMPL_WIDTH - 1),
		31977 => to_unsigned(2483, LUT_AMPL_WIDTH - 1),
		31978 => to_unsigned(2479, LUT_AMPL_WIDTH - 1),
		31979 => to_unsigned(2476, LUT_AMPL_WIDTH - 1),
		31980 => to_unsigned(2473, LUT_AMPL_WIDTH - 1),
		31981 => to_unsigned(2470, LUT_AMPL_WIDTH - 1),
		31982 => to_unsigned(2467, LUT_AMPL_WIDTH - 1),
		31983 => to_unsigned(2464, LUT_AMPL_WIDTH - 1),
		31984 => to_unsigned(2461, LUT_AMPL_WIDTH - 1),
		31985 => to_unsigned(2457, LUT_AMPL_WIDTH - 1),
		31986 => to_unsigned(2454, LUT_AMPL_WIDTH - 1),
		31987 => to_unsigned(2451, LUT_AMPL_WIDTH - 1),
		31988 => to_unsigned(2448, LUT_AMPL_WIDTH - 1),
		31989 => to_unsigned(2445, LUT_AMPL_WIDTH - 1),
		31990 => to_unsigned(2442, LUT_AMPL_WIDTH - 1),
		31991 => to_unsigned(2439, LUT_AMPL_WIDTH - 1),
		31992 => to_unsigned(2436, LUT_AMPL_WIDTH - 1),
		31993 => to_unsigned(2432, LUT_AMPL_WIDTH - 1),
		31994 => to_unsigned(2429, LUT_AMPL_WIDTH - 1),
		31995 => to_unsigned(2426, LUT_AMPL_WIDTH - 1),
		31996 => to_unsigned(2423, LUT_AMPL_WIDTH - 1),
		31997 => to_unsigned(2420, LUT_AMPL_WIDTH - 1),
		31998 => to_unsigned(2417, LUT_AMPL_WIDTH - 1),
		31999 => to_unsigned(2414, LUT_AMPL_WIDTH - 1),
		32000 => to_unsigned(2410, LUT_AMPL_WIDTH - 1),
		32001 => to_unsigned(2407, LUT_AMPL_WIDTH - 1),
		32002 => to_unsigned(2404, LUT_AMPL_WIDTH - 1),
		32003 => to_unsigned(2401, LUT_AMPL_WIDTH - 1),
		32004 => to_unsigned(2398, LUT_AMPL_WIDTH - 1),
		32005 => to_unsigned(2395, LUT_AMPL_WIDTH - 1),
		32006 => to_unsigned(2392, LUT_AMPL_WIDTH - 1),
		32007 => to_unsigned(2389, LUT_AMPL_WIDTH - 1),
		32008 => to_unsigned(2385, LUT_AMPL_WIDTH - 1),
		32009 => to_unsigned(2382, LUT_AMPL_WIDTH - 1),
		32010 => to_unsigned(2379, LUT_AMPL_WIDTH - 1),
		32011 => to_unsigned(2376, LUT_AMPL_WIDTH - 1),
		32012 => to_unsigned(2373, LUT_AMPL_WIDTH - 1),
		32013 => to_unsigned(2370, LUT_AMPL_WIDTH - 1),
		32014 => to_unsigned(2367, LUT_AMPL_WIDTH - 1),
		32015 => to_unsigned(2363, LUT_AMPL_WIDTH - 1),
		32016 => to_unsigned(2360, LUT_AMPL_WIDTH - 1),
		32017 => to_unsigned(2357, LUT_AMPL_WIDTH - 1),
		32018 => to_unsigned(2354, LUT_AMPL_WIDTH - 1),
		32019 => to_unsigned(2351, LUT_AMPL_WIDTH - 1),
		32020 => to_unsigned(2348, LUT_AMPL_WIDTH - 1),
		32021 => to_unsigned(2345, LUT_AMPL_WIDTH - 1),
		32022 => to_unsigned(2342, LUT_AMPL_WIDTH - 1),
		32023 => to_unsigned(2338, LUT_AMPL_WIDTH - 1),
		32024 => to_unsigned(2335, LUT_AMPL_WIDTH - 1),
		32025 => to_unsigned(2332, LUT_AMPL_WIDTH - 1),
		32026 => to_unsigned(2329, LUT_AMPL_WIDTH - 1),
		32027 => to_unsigned(2326, LUT_AMPL_WIDTH - 1),
		32028 => to_unsigned(2323, LUT_AMPL_WIDTH - 1),
		32029 => to_unsigned(2320, LUT_AMPL_WIDTH - 1),
		32030 => to_unsigned(2316, LUT_AMPL_WIDTH - 1),
		32031 => to_unsigned(2313, LUT_AMPL_WIDTH - 1),
		32032 => to_unsigned(2310, LUT_AMPL_WIDTH - 1),
		32033 => to_unsigned(2307, LUT_AMPL_WIDTH - 1),
		32034 => to_unsigned(2304, LUT_AMPL_WIDTH - 1),
		32035 => to_unsigned(2301, LUT_AMPL_WIDTH - 1),
		32036 => to_unsigned(2298, LUT_AMPL_WIDTH - 1),
		32037 => to_unsigned(2295, LUT_AMPL_WIDTH - 1),
		32038 => to_unsigned(2291, LUT_AMPL_WIDTH - 1),
		32039 => to_unsigned(2288, LUT_AMPL_WIDTH - 1),
		32040 => to_unsigned(2285, LUT_AMPL_WIDTH - 1),
		32041 => to_unsigned(2282, LUT_AMPL_WIDTH - 1),
		32042 => to_unsigned(2279, LUT_AMPL_WIDTH - 1),
		32043 => to_unsigned(2276, LUT_AMPL_WIDTH - 1),
		32044 => to_unsigned(2273, LUT_AMPL_WIDTH - 1),
		32045 => to_unsigned(2269, LUT_AMPL_WIDTH - 1),
		32046 => to_unsigned(2266, LUT_AMPL_WIDTH - 1),
		32047 => to_unsigned(2263, LUT_AMPL_WIDTH - 1),
		32048 => to_unsigned(2260, LUT_AMPL_WIDTH - 1),
		32049 => to_unsigned(2257, LUT_AMPL_WIDTH - 1),
		32050 => to_unsigned(2254, LUT_AMPL_WIDTH - 1),
		32051 => to_unsigned(2251, LUT_AMPL_WIDTH - 1),
		32052 => to_unsigned(2248, LUT_AMPL_WIDTH - 1),
		32053 => to_unsigned(2244, LUT_AMPL_WIDTH - 1),
		32054 => to_unsigned(2241, LUT_AMPL_WIDTH - 1),
		32055 => to_unsigned(2238, LUT_AMPL_WIDTH - 1),
		32056 => to_unsigned(2235, LUT_AMPL_WIDTH - 1),
		32057 => to_unsigned(2232, LUT_AMPL_WIDTH - 1),
		32058 => to_unsigned(2229, LUT_AMPL_WIDTH - 1),
		32059 => to_unsigned(2226, LUT_AMPL_WIDTH - 1),
		32060 => to_unsigned(2222, LUT_AMPL_WIDTH - 1),
		32061 => to_unsigned(2219, LUT_AMPL_WIDTH - 1),
		32062 => to_unsigned(2216, LUT_AMPL_WIDTH - 1),
		32063 => to_unsigned(2213, LUT_AMPL_WIDTH - 1),
		32064 => to_unsigned(2210, LUT_AMPL_WIDTH - 1),
		32065 => to_unsigned(2207, LUT_AMPL_WIDTH - 1),
		32066 => to_unsigned(2204, LUT_AMPL_WIDTH - 1),
		32067 => to_unsigned(2201, LUT_AMPL_WIDTH - 1),
		32068 => to_unsigned(2197, LUT_AMPL_WIDTH - 1),
		32069 => to_unsigned(2194, LUT_AMPL_WIDTH - 1),
		32070 => to_unsigned(2191, LUT_AMPL_WIDTH - 1),
		32071 => to_unsigned(2188, LUT_AMPL_WIDTH - 1),
		32072 => to_unsigned(2185, LUT_AMPL_WIDTH - 1),
		32073 => to_unsigned(2182, LUT_AMPL_WIDTH - 1),
		32074 => to_unsigned(2179, LUT_AMPL_WIDTH - 1),
		32075 => to_unsigned(2175, LUT_AMPL_WIDTH - 1),
		32076 => to_unsigned(2172, LUT_AMPL_WIDTH - 1),
		32077 => to_unsigned(2169, LUT_AMPL_WIDTH - 1),
		32078 => to_unsigned(2166, LUT_AMPL_WIDTH - 1),
		32079 => to_unsigned(2163, LUT_AMPL_WIDTH - 1),
		32080 => to_unsigned(2160, LUT_AMPL_WIDTH - 1),
		32081 => to_unsigned(2157, LUT_AMPL_WIDTH - 1),
		32082 => to_unsigned(2154, LUT_AMPL_WIDTH - 1),
		32083 => to_unsigned(2150, LUT_AMPL_WIDTH - 1),
		32084 => to_unsigned(2147, LUT_AMPL_WIDTH - 1),
		32085 => to_unsigned(2144, LUT_AMPL_WIDTH - 1),
		32086 => to_unsigned(2141, LUT_AMPL_WIDTH - 1),
		32087 => to_unsigned(2138, LUT_AMPL_WIDTH - 1),
		32088 => to_unsigned(2135, LUT_AMPL_WIDTH - 1),
		32089 => to_unsigned(2132, LUT_AMPL_WIDTH - 1),
		32090 => to_unsigned(2128, LUT_AMPL_WIDTH - 1),
		32091 => to_unsigned(2125, LUT_AMPL_WIDTH - 1),
		32092 => to_unsigned(2122, LUT_AMPL_WIDTH - 1),
		32093 => to_unsigned(2119, LUT_AMPL_WIDTH - 1),
		32094 => to_unsigned(2116, LUT_AMPL_WIDTH - 1),
		32095 => to_unsigned(2113, LUT_AMPL_WIDTH - 1),
		32096 => to_unsigned(2110, LUT_AMPL_WIDTH - 1),
		32097 => to_unsigned(2106, LUT_AMPL_WIDTH - 1),
		32098 => to_unsigned(2103, LUT_AMPL_WIDTH - 1),
		32099 => to_unsigned(2100, LUT_AMPL_WIDTH - 1),
		32100 => to_unsigned(2097, LUT_AMPL_WIDTH - 1),
		32101 => to_unsigned(2094, LUT_AMPL_WIDTH - 1),
		32102 => to_unsigned(2091, LUT_AMPL_WIDTH - 1),
		32103 => to_unsigned(2088, LUT_AMPL_WIDTH - 1),
		32104 => to_unsigned(2085, LUT_AMPL_WIDTH - 1),
		32105 => to_unsigned(2081, LUT_AMPL_WIDTH - 1),
		32106 => to_unsigned(2078, LUT_AMPL_WIDTH - 1),
		32107 => to_unsigned(2075, LUT_AMPL_WIDTH - 1),
		32108 => to_unsigned(2072, LUT_AMPL_WIDTH - 1),
		32109 => to_unsigned(2069, LUT_AMPL_WIDTH - 1),
		32110 => to_unsigned(2066, LUT_AMPL_WIDTH - 1),
		32111 => to_unsigned(2063, LUT_AMPL_WIDTH - 1),
		32112 => to_unsigned(2059, LUT_AMPL_WIDTH - 1),
		32113 => to_unsigned(2056, LUT_AMPL_WIDTH - 1),
		32114 => to_unsigned(2053, LUT_AMPL_WIDTH - 1),
		32115 => to_unsigned(2050, LUT_AMPL_WIDTH - 1),
		32116 => to_unsigned(2047, LUT_AMPL_WIDTH - 1),
		32117 => to_unsigned(2044, LUT_AMPL_WIDTH - 1),
		32118 => to_unsigned(2041, LUT_AMPL_WIDTH - 1),
		32119 => to_unsigned(2038, LUT_AMPL_WIDTH - 1),
		32120 => to_unsigned(2034, LUT_AMPL_WIDTH - 1),
		32121 => to_unsigned(2031, LUT_AMPL_WIDTH - 1),
		32122 => to_unsigned(2028, LUT_AMPL_WIDTH - 1),
		32123 => to_unsigned(2025, LUT_AMPL_WIDTH - 1),
		32124 => to_unsigned(2022, LUT_AMPL_WIDTH - 1),
		32125 => to_unsigned(2019, LUT_AMPL_WIDTH - 1),
		32126 => to_unsigned(2016, LUT_AMPL_WIDTH - 1),
		32127 => to_unsigned(2012, LUT_AMPL_WIDTH - 1),
		32128 => to_unsigned(2009, LUT_AMPL_WIDTH - 1),
		32129 => to_unsigned(2006, LUT_AMPL_WIDTH - 1),
		32130 => to_unsigned(2003, LUT_AMPL_WIDTH - 1),
		32131 => to_unsigned(2000, LUT_AMPL_WIDTH - 1),
		32132 => to_unsigned(1997, LUT_AMPL_WIDTH - 1),
		32133 => to_unsigned(1994, LUT_AMPL_WIDTH - 1),
		32134 => to_unsigned(1990, LUT_AMPL_WIDTH - 1),
		32135 => to_unsigned(1987, LUT_AMPL_WIDTH - 1),
		32136 => to_unsigned(1984, LUT_AMPL_WIDTH - 1),
		32137 => to_unsigned(1981, LUT_AMPL_WIDTH - 1),
		32138 => to_unsigned(1978, LUT_AMPL_WIDTH - 1),
		32139 => to_unsigned(1975, LUT_AMPL_WIDTH - 1),
		32140 => to_unsigned(1972, LUT_AMPL_WIDTH - 1),
		32141 => to_unsigned(1969, LUT_AMPL_WIDTH - 1),
		32142 => to_unsigned(1965, LUT_AMPL_WIDTH - 1),
		32143 => to_unsigned(1962, LUT_AMPL_WIDTH - 1),
		32144 => to_unsigned(1959, LUT_AMPL_WIDTH - 1),
		32145 => to_unsigned(1956, LUT_AMPL_WIDTH - 1),
		32146 => to_unsigned(1953, LUT_AMPL_WIDTH - 1),
		32147 => to_unsigned(1950, LUT_AMPL_WIDTH - 1),
		32148 => to_unsigned(1947, LUT_AMPL_WIDTH - 1),
		32149 => to_unsigned(1943, LUT_AMPL_WIDTH - 1),
		32150 => to_unsigned(1940, LUT_AMPL_WIDTH - 1),
		32151 => to_unsigned(1937, LUT_AMPL_WIDTH - 1),
		32152 => to_unsigned(1934, LUT_AMPL_WIDTH - 1),
		32153 => to_unsigned(1931, LUT_AMPL_WIDTH - 1),
		32154 => to_unsigned(1928, LUT_AMPL_WIDTH - 1),
		32155 => to_unsigned(1925, LUT_AMPL_WIDTH - 1),
		32156 => to_unsigned(1921, LUT_AMPL_WIDTH - 1),
		32157 => to_unsigned(1918, LUT_AMPL_WIDTH - 1),
		32158 => to_unsigned(1915, LUT_AMPL_WIDTH - 1),
		32159 => to_unsigned(1912, LUT_AMPL_WIDTH - 1),
		32160 => to_unsigned(1909, LUT_AMPL_WIDTH - 1),
		32161 => to_unsigned(1906, LUT_AMPL_WIDTH - 1),
		32162 => to_unsigned(1903, LUT_AMPL_WIDTH - 1),
		32163 => to_unsigned(1900, LUT_AMPL_WIDTH - 1),
		32164 => to_unsigned(1896, LUT_AMPL_WIDTH - 1),
		32165 => to_unsigned(1893, LUT_AMPL_WIDTH - 1),
		32166 => to_unsigned(1890, LUT_AMPL_WIDTH - 1),
		32167 => to_unsigned(1887, LUT_AMPL_WIDTH - 1),
		32168 => to_unsigned(1884, LUT_AMPL_WIDTH - 1),
		32169 => to_unsigned(1881, LUT_AMPL_WIDTH - 1),
		32170 => to_unsigned(1878, LUT_AMPL_WIDTH - 1),
		32171 => to_unsigned(1874, LUT_AMPL_WIDTH - 1),
		32172 => to_unsigned(1871, LUT_AMPL_WIDTH - 1),
		32173 => to_unsigned(1868, LUT_AMPL_WIDTH - 1),
		32174 => to_unsigned(1865, LUT_AMPL_WIDTH - 1),
		32175 => to_unsigned(1862, LUT_AMPL_WIDTH - 1),
		32176 => to_unsigned(1859, LUT_AMPL_WIDTH - 1),
		32177 => to_unsigned(1856, LUT_AMPL_WIDTH - 1),
		32178 => to_unsigned(1852, LUT_AMPL_WIDTH - 1),
		32179 => to_unsigned(1849, LUT_AMPL_WIDTH - 1),
		32180 => to_unsigned(1846, LUT_AMPL_WIDTH - 1),
		32181 => to_unsigned(1843, LUT_AMPL_WIDTH - 1),
		32182 => to_unsigned(1840, LUT_AMPL_WIDTH - 1),
		32183 => to_unsigned(1837, LUT_AMPL_WIDTH - 1),
		32184 => to_unsigned(1834, LUT_AMPL_WIDTH - 1),
		32185 => to_unsigned(1831, LUT_AMPL_WIDTH - 1),
		32186 => to_unsigned(1827, LUT_AMPL_WIDTH - 1),
		32187 => to_unsigned(1824, LUT_AMPL_WIDTH - 1),
		32188 => to_unsigned(1821, LUT_AMPL_WIDTH - 1),
		32189 => to_unsigned(1818, LUT_AMPL_WIDTH - 1),
		32190 => to_unsigned(1815, LUT_AMPL_WIDTH - 1),
		32191 => to_unsigned(1812, LUT_AMPL_WIDTH - 1),
		32192 => to_unsigned(1809, LUT_AMPL_WIDTH - 1),
		32193 => to_unsigned(1805, LUT_AMPL_WIDTH - 1),
		32194 => to_unsigned(1802, LUT_AMPL_WIDTH - 1),
		32195 => to_unsigned(1799, LUT_AMPL_WIDTH - 1),
		32196 => to_unsigned(1796, LUT_AMPL_WIDTH - 1),
		32197 => to_unsigned(1793, LUT_AMPL_WIDTH - 1),
		32198 => to_unsigned(1790, LUT_AMPL_WIDTH - 1),
		32199 => to_unsigned(1787, LUT_AMPL_WIDTH - 1),
		32200 => to_unsigned(1783, LUT_AMPL_WIDTH - 1),
		32201 => to_unsigned(1780, LUT_AMPL_WIDTH - 1),
		32202 => to_unsigned(1777, LUT_AMPL_WIDTH - 1),
		32203 => to_unsigned(1774, LUT_AMPL_WIDTH - 1),
		32204 => to_unsigned(1771, LUT_AMPL_WIDTH - 1),
		32205 => to_unsigned(1768, LUT_AMPL_WIDTH - 1),
		32206 => to_unsigned(1765, LUT_AMPL_WIDTH - 1),
		32207 => to_unsigned(1762, LUT_AMPL_WIDTH - 1),
		32208 => to_unsigned(1758, LUT_AMPL_WIDTH - 1),
		32209 => to_unsigned(1755, LUT_AMPL_WIDTH - 1),
		32210 => to_unsigned(1752, LUT_AMPL_WIDTH - 1),
		32211 => to_unsigned(1749, LUT_AMPL_WIDTH - 1),
		32212 => to_unsigned(1746, LUT_AMPL_WIDTH - 1),
		32213 => to_unsigned(1743, LUT_AMPL_WIDTH - 1),
		32214 => to_unsigned(1740, LUT_AMPL_WIDTH - 1),
		32215 => to_unsigned(1736, LUT_AMPL_WIDTH - 1),
		32216 => to_unsigned(1733, LUT_AMPL_WIDTH - 1),
		32217 => to_unsigned(1730, LUT_AMPL_WIDTH - 1),
		32218 => to_unsigned(1727, LUT_AMPL_WIDTH - 1),
		32219 => to_unsigned(1724, LUT_AMPL_WIDTH - 1),
		32220 => to_unsigned(1721, LUT_AMPL_WIDTH - 1),
		32221 => to_unsigned(1718, LUT_AMPL_WIDTH - 1),
		32222 => to_unsigned(1714, LUT_AMPL_WIDTH - 1),
		32223 => to_unsigned(1711, LUT_AMPL_WIDTH - 1),
		32224 => to_unsigned(1708, LUT_AMPL_WIDTH - 1),
		32225 => to_unsigned(1705, LUT_AMPL_WIDTH - 1),
		32226 => to_unsigned(1702, LUT_AMPL_WIDTH - 1),
		32227 => to_unsigned(1699, LUT_AMPL_WIDTH - 1),
		32228 => to_unsigned(1696, LUT_AMPL_WIDTH - 1),
		32229 => to_unsigned(1693, LUT_AMPL_WIDTH - 1),
		32230 => to_unsigned(1689, LUT_AMPL_WIDTH - 1),
		32231 => to_unsigned(1686, LUT_AMPL_WIDTH - 1),
		32232 => to_unsigned(1683, LUT_AMPL_WIDTH - 1),
		32233 => to_unsigned(1680, LUT_AMPL_WIDTH - 1),
		32234 => to_unsigned(1677, LUT_AMPL_WIDTH - 1),
		32235 => to_unsigned(1674, LUT_AMPL_WIDTH - 1),
		32236 => to_unsigned(1671, LUT_AMPL_WIDTH - 1),
		32237 => to_unsigned(1667, LUT_AMPL_WIDTH - 1),
		32238 => to_unsigned(1664, LUT_AMPL_WIDTH - 1),
		32239 => to_unsigned(1661, LUT_AMPL_WIDTH - 1),
		32240 => to_unsigned(1658, LUT_AMPL_WIDTH - 1),
		32241 => to_unsigned(1655, LUT_AMPL_WIDTH - 1),
		32242 => to_unsigned(1652, LUT_AMPL_WIDTH - 1),
		32243 => to_unsigned(1649, LUT_AMPL_WIDTH - 1),
		32244 => to_unsigned(1645, LUT_AMPL_WIDTH - 1),
		32245 => to_unsigned(1642, LUT_AMPL_WIDTH - 1),
		32246 => to_unsigned(1639, LUT_AMPL_WIDTH - 1),
		32247 => to_unsigned(1636, LUT_AMPL_WIDTH - 1),
		32248 => to_unsigned(1633, LUT_AMPL_WIDTH - 1),
		32249 => to_unsigned(1630, LUT_AMPL_WIDTH - 1),
		32250 => to_unsigned(1627, LUT_AMPL_WIDTH - 1),
		32251 => to_unsigned(1623, LUT_AMPL_WIDTH - 1),
		32252 => to_unsigned(1620, LUT_AMPL_WIDTH - 1),
		32253 => to_unsigned(1617, LUT_AMPL_WIDTH - 1),
		32254 => to_unsigned(1614, LUT_AMPL_WIDTH - 1),
		32255 => to_unsigned(1611, LUT_AMPL_WIDTH - 1),
		32256 => to_unsigned(1608, LUT_AMPL_WIDTH - 1),
		32257 => to_unsigned(1605, LUT_AMPL_WIDTH - 1),
		32258 => to_unsigned(1602, LUT_AMPL_WIDTH - 1),
		32259 => to_unsigned(1598, LUT_AMPL_WIDTH - 1),
		32260 => to_unsigned(1595, LUT_AMPL_WIDTH - 1),
		32261 => to_unsigned(1592, LUT_AMPL_WIDTH - 1),
		32262 => to_unsigned(1589, LUT_AMPL_WIDTH - 1),
		32263 => to_unsigned(1586, LUT_AMPL_WIDTH - 1),
		32264 => to_unsigned(1583, LUT_AMPL_WIDTH - 1),
		32265 => to_unsigned(1580, LUT_AMPL_WIDTH - 1),
		32266 => to_unsigned(1576, LUT_AMPL_WIDTH - 1),
		32267 => to_unsigned(1573, LUT_AMPL_WIDTH - 1),
		32268 => to_unsigned(1570, LUT_AMPL_WIDTH - 1),
		32269 => to_unsigned(1567, LUT_AMPL_WIDTH - 1),
		32270 => to_unsigned(1564, LUT_AMPL_WIDTH - 1),
		32271 => to_unsigned(1561, LUT_AMPL_WIDTH - 1),
		32272 => to_unsigned(1558, LUT_AMPL_WIDTH - 1),
		32273 => to_unsigned(1554, LUT_AMPL_WIDTH - 1),
		32274 => to_unsigned(1551, LUT_AMPL_WIDTH - 1),
		32275 => to_unsigned(1548, LUT_AMPL_WIDTH - 1),
		32276 => to_unsigned(1545, LUT_AMPL_WIDTH - 1),
		32277 => to_unsigned(1542, LUT_AMPL_WIDTH - 1),
		32278 => to_unsigned(1539, LUT_AMPL_WIDTH - 1),
		32279 => to_unsigned(1536, LUT_AMPL_WIDTH - 1),
		32280 => to_unsigned(1532, LUT_AMPL_WIDTH - 1),
		32281 => to_unsigned(1529, LUT_AMPL_WIDTH - 1),
		32282 => to_unsigned(1526, LUT_AMPL_WIDTH - 1),
		32283 => to_unsigned(1523, LUT_AMPL_WIDTH - 1),
		32284 => to_unsigned(1520, LUT_AMPL_WIDTH - 1),
		32285 => to_unsigned(1517, LUT_AMPL_WIDTH - 1),
		32286 => to_unsigned(1514, LUT_AMPL_WIDTH - 1),
		32287 => to_unsigned(1511, LUT_AMPL_WIDTH - 1),
		32288 => to_unsigned(1507, LUT_AMPL_WIDTH - 1),
		32289 => to_unsigned(1504, LUT_AMPL_WIDTH - 1),
		32290 => to_unsigned(1501, LUT_AMPL_WIDTH - 1),
		32291 => to_unsigned(1498, LUT_AMPL_WIDTH - 1),
		32292 => to_unsigned(1495, LUT_AMPL_WIDTH - 1),
		32293 => to_unsigned(1492, LUT_AMPL_WIDTH - 1),
		32294 => to_unsigned(1489, LUT_AMPL_WIDTH - 1),
		32295 => to_unsigned(1485, LUT_AMPL_WIDTH - 1),
		32296 => to_unsigned(1482, LUT_AMPL_WIDTH - 1),
		32297 => to_unsigned(1479, LUT_AMPL_WIDTH - 1),
		32298 => to_unsigned(1476, LUT_AMPL_WIDTH - 1),
		32299 => to_unsigned(1473, LUT_AMPL_WIDTH - 1),
		32300 => to_unsigned(1470, LUT_AMPL_WIDTH - 1),
		32301 => to_unsigned(1467, LUT_AMPL_WIDTH - 1),
		32302 => to_unsigned(1463, LUT_AMPL_WIDTH - 1),
		32303 => to_unsigned(1460, LUT_AMPL_WIDTH - 1),
		32304 => to_unsigned(1457, LUT_AMPL_WIDTH - 1),
		32305 => to_unsigned(1454, LUT_AMPL_WIDTH - 1),
		32306 => to_unsigned(1451, LUT_AMPL_WIDTH - 1),
		32307 => to_unsigned(1448, LUT_AMPL_WIDTH - 1),
		32308 => to_unsigned(1445, LUT_AMPL_WIDTH - 1),
		32309 => to_unsigned(1441, LUT_AMPL_WIDTH - 1),
		32310 => to_unsigned(1438, LUT_AMPL_WIDTH - 1),
		32311 => to_unsigned(1435, LUT_AMPL_WIDTH - 1),
		32312 => to_unsigned(1432, LUT_AMPL_WIDTH - 1),
		32313 => to_unsigned(1429, LUT_AMPL_WIDTH - 1),
		32314 => to_unsigned(1426, LUT_AMPL_WIDTH - 1),
		32315 => to_unsigned(1423, LUT_AMPL_WIDTH - 1),
		32316 => to_unsigned(1420, LUT_AMPL_WIDTH - 1),
		32317 => to_unsigned(1416, LUT_AMPL_WIDTH - 1),
		32318 => to_unsigned(1413, LUT_AMPL_WIDTH - 1),
		32319 => to_unsigned(1410, LUT_AMPL_WIDTH - 1),
		32320 => to_unsigned(1407, LUT_AMPL_WIDTH - 1),
		32321 => to_unsigned(1404, LUT_AMPL_WIDTH - 1),
		32322 => to_unsigned(1401, LUT_AMPL_WIDTH - 1),
		32323 => to_unsigned(1398, LUT_AMPL_WIDTH - 1),
		32324 => to_unsigned(1394, LUT_AMPL_WIDTH - 1),
		32325 => to_unsigned(1391, LUT_AMPL_WIDTH - 1),
		32326 => to_unsigned(1388, LUT_AMPL_WIDTH - 1),
		32327 => to_unsigned(1385, LUT_AMPL_WIDTH - 1),
		32328 => to_unsigned(1382, LUT_AMPL_WIDTH - 1),
		32329 => to_unsigned(1379, LUT_AMPL_WIDTH - 1),
		32330 => to_unsigned(1376, LUT_AMPL_WIDTH - 1),
		32331 => to_unsigned(1372, LUT_AMPL_WIDTH - 1),
		32332 => to_unsigned(1369, LUT_AMPL_WIDTH - 1),
		32333 => to_unsigned(1366, LUT_AMPL_WIDTH - 1),
		32334 => to_unsigned(1363, LUT_AMPL_WIDTH - 1),
		32335 => to_unsigned(1360, LUT_AMPL_WIDTH - 1),
		32336 => to_unsigned(1357, LUT_AMPL_WIDTH - 1),
		32337 => to_unsigned(1354, LUT_AMPL_WIDTH - 1),
		32338 => to_unsigned(1350, LUT_AMPL_WIDTH - 1),
		32339 => to_unsigned(1347, LUT_AMPL_WIDTH - 1),
		32340 => to_unsigned(1344, LUT_AMPL_WIDTH - 1),
		32341 => to_unsigned(1341, LUT_AMPL_WIDTH - 1),
		32342 => to_unsigned(1338, LUT_AMPL_WIDTH - 1),
		32343 => to_unsigned(1335, LUT_AMPL_WIDTH - 1),
		32344 => to_unsigned(1332, LUT_AMPL_WIDTH - 1),
		32345 => to_unsigned(1328, LUT_AMPL_WIDTH - 1),
		32346 => to_unsigned(1325, LUT_AMPL_WIDTH - 1),
		32347 => to_unsigned(1322, LUT_AMPL_WIDTH - 1),
		32348 => to_unsigned(1319, LUT_AMPL_WIDTH - 1),
		32349 => to_unsigned(1316, LUT_AMPL_WIDTH - 1),
		32350 => to_unsigned(1313, LUT_AMPL_WIDTH - 1),
		32351 => to_unsigned(1310, LUT_AMPL_WIDTH - 1),
		32352 => to_unsigned(1307, LUT_AMPL_WIDTH - 1),
		32353 => to_unsigned(1303, LUT_AMPL_WIDTH - 1),
		32354 => to_unsigned(1300, LUT_AMPL_WIDTH - 1),
		32355 => to_unsigned(1297, LUT_AMPL_WIDTH - 1),
		32356 => to_unsigned(1294, LUT_AMPL_WIDTH - 1),
		32357 => to_unsigned(1291, LUT_AMPL_WIDTH - 1),
		32358 => to_unsigned(1288, LUT_AMPL_WIDTH - 1),
		32359 => to_unsigned(1285, LUT_AMPL_WIDTH - 1),
		32360 => to_unsigned(1281, LUT_AMPL_WIDTH - 1),
		32361 => to_unsigned(1278, LUT_AMPL_WIDTH - 1),
		32362 => to_unsigned(1275, LUT_AMPL_WIDTH - 1),
		32363 => to_unsigned(1272, LUT_AMPL_WIDTH - 1),
		32364 => to_unsigned(1269, LUT_AMPL_WIDTH - 1),
		32365 => to_unsigned(1266, LUT_AMPL_WIDTH - 1),
		32366 => to_unsigned(1263, LUT_AMPL_WIDTH - 1),
		32367 => to_unsigned(1259, LUT_AMPL_WIDTH - 1),
		32368 => to_unsigned(1256, LUT_AMPL_WIDTH - 1),
		32369 => to_unsigned(1253, LUT_AMPL_WIDTH - 1),
		32370 => to_unsigned(1250, LUT_AMPL_WIDTH - 1),
		32371 => to_unsigned(1247, LUT_AMPL_WIDTH - 1),
		32372 => to_unsigned(1244, LUT_AMPL_WIDTH - 1),
		32373 => to_unsigned(1241, LUT_AMPL_WIDTH - 1),
		32374 => to_unsigned(1237, LUT_AMPL_WIDTH - 1),
		32375 => to_unsigned(1234, LUT_AMPL_WIDTH - 1),
		32376 => to_unsigned(1231, LUT_AMPL_WIDTH - 1),
		32377 => to_unsigned(1228, LUT_AMPL_WIDTH - 1),
		32378 => to_unsigned(1225, LUT_AMPL_WIDTH - 1),
		32379 => to_unsigned(1222, LUT_AMPL_WIDTH - 1),
		32380 => to_unsigned(1219, LUT_AMPL_WIDTH - 1),
		32381 => to_unsigned(1215, LUT_AMPL_WIDTH - 1),
		32382 => to_unsigned(1212, LUT_AMPL_WIDTH - 1),
		32383 => to_unsigned(1209, LUT_AMPL_WIDTH - 1),
		32384 => to_unsigned(1206, LUT_AMPL_WIDTH - 1),
		32385 => to_unsigned(1203, LUT_AMPL_WIDTH - 1),
		32386 => to_unsigned(1200, LUT_AMPL_WIDTH - 1),
		32387 => to_unsigned(1197, LUT_AMPL_WIDTH - 1),
		32388 => to_unsigned(1194, LUT_AMPL_WIDTH - 1),
		32389 => to_unsigned(1190, LUT_AMPL_WIDTH - 1),
		32390 => to_unsigned(1187, LUT_AMPL_WIDTH - 1),
		32391 => to_unsigned(1184, LUT_AMPL_WIDTH - 1),
		32392 => to_unsigned(1181, LUT_AMPL_WIDTH - 1),
		32393 => to_unsigned(1178, LUT_AMPL_WIDTH - 1),
		32394 => to_unsigned(1175, LUT_AMPL_WIDTH - 1),
		32395 => to_unsigned(1172, LUT_AMPL_WIDTH - 1),
		32396 => to_unsigned(1168, LUT_AMPL_WIDTH - 1),
		32397 => to_unsigned(1165, LUT_AMPL_WIDTH - 1),
		32398 => to_unsigned(1162, LUT_AMPL_WIDTH - 1),
		32399 => to_unsigned(1159, LUT_AMPL_WIDTH - 1),
		32400 => to_unsigned(1156, LUT_AMPL_WIDTH - 1),
		32401 => to_unsigned(1153, LUT_AMPL_WIDTH - 1),
		32402 => to_unsigned(1150, LUT_AMPL_WIDTH - 1),
		32403 => to_unsigned(1146, LUT_AMPL_WIDTH - 1),
		32404 => to_unsigned(1143, LUT_AMPL_WIDTH - 1),
		32405 => to_unsigned(1140, LUT_AMPL_WIDTH - 1),
		32406 => to_unsigned(1137, LUT_AMPL_WIDTH - 1),
		32407 => to_unsigned(1134, LUT_AMPL_WIDTH - 1),
		32408 => to_unsigned(1131, LUT_AMPL_WIDTH - 1),
		32409 => to_unsigned(1128, LUT_AMPL_WIDTH - 1),
		32410 => to_unsigned(1124, LUT_AMPL_WIDTH - 1),
		32411 => to_unsigned(1121, LUT_AMPL_WIDTH - 1),
		32412 => to_unsigned(1118, LUT_AMPL_WIDTH - 1),
		32413 => to_unsigned(1115, LUT_AMPL_WIDTH - 1),
		32414 => to_unsigned(1112, LUT_AMPL_WIDTH - 1),
		32415 => to_unsigned(1109, LUT_AMPL_WIDTH - 1),
		32416 => to_unsigned(1106, LUT_AMPL_WIDTH - 1),
		32417 => to_unsigned(1102, LUT_AMPL_WIDTH - 1),
		32418 => to_unsigned(1099, LUT_AMPL_WIDTH - 1),
		32419 => to_unsigned(1096, LUT_AMPL_WIDTH - 1),
		32420 => to_unsigned(1093, LUT_AMPL_WIDTH - 1),
		32421 => to_unsigned(1090, LUT_AMPL_WIDTH - 1),
		32422 => to_unsigned(1087, LUT_AMPL_WIDTH - 1),
		32423 => to_unsigned(1084, LUT_AMPL_WIDTH - 1),
		32424 => to_unsigned(1080, LUT_AMPL_WIDTH - 1),
		32425 => to_unsigned(1077, LUT_AMPL_WIDTH - 1),
		32426 => to_unsigned(1074, LUT_AMPL_WIDTH - 1),
		32427 => to_unsigned(1071, LUT_AMPL_WIDTH - 1),
		32428 => to_unsigned(1068, LUT_AMPL_WIDTH - 1),
		32429 => to_unsigned(1065, LUT_AMPL_WIDTH - 1),
		32430 => to_unsigned(1062, LUT_AMPL_WIDTH - 1),
		32431 => to_unsigned(1059, LUT_AMPL_WIDTH - 1),
		32432 => to_unsigned(1055, LUT_AMPL_WIDTH - 1),
		32433 => to_unsigned(1052, LUT_AMPL_WIDTH - 1),
		32434 => to_unsigned(1049, LUT_AMPL_WIDTH - 1),
		32435 => to_unsigned(1046, LUT_AMPL_WIDTH - 1),
		32436 => to_unsigned(1043, LUT_AMPL_WIDTH - 1),
		32437 => to_unsigned(1040, LUT_AMPL_WIDTH - 1),
		32438 => to_unsigned(1037, LUT_AMPL_WIDTH - 1),
		32439 => to_unsigned(1033, LUT_AMPL_WIDTH - 1),
		32440 => to_unsigned(1030, LUT_AMPL_WIDTH - 1),
		32441 => to_unsigned(1027, LUT_AMPL_WIDTH - 1),
		32442 => to_unsigned(1024, LUT_AMPL_WIDTH - 1),
		32443 => to_unsigned(1021, LUT_AMPL_WIDTH - 1),
		32444 => to_unsigned(1018, LUT_AMPL_WIDTH - 1),
		32445 => to_unsigned(1015, LUT_AMPL_WIDTH - 1),
		32446 => to_unsigned(1011, LUT_AMPL_WIDTH - 1),
		32447 => to_unsigned(1008, LUT_AMPL_WIDTH - 1),
		32448 => to_unsigned(1005, LUT_AMPL_WIDTH - 1),
		32449 => to_unsigned(1002, LUT_AMPL_WIDTH - 1),
		32450 => to_unsigned(999, LUT_AMPL_WIDTH - 1),
		32451 => to_unsigned(996, LUT_AMPL_WIDTH - 1),
		32452 => to_unsigned(993, LUT_AMPL_WIDTH - 1),
		32453 => to_unsigned(989, LUT_AMPL_WIDTH - 1),
		32454 => to_unsigned(986, LUT_AMPL_WIDTH - 1),
		32455 => to_unsigned(983, LUT_AMPL_WIDTH - 1),
		32456 => to_unsigned(980, LUT_AMPL_WIDTH - 1),
		32457 => to_unsigned(977, LUT_AMPL_WIDTH - 1),
		32458 => to_unsigned(974, LUT_AMPL_WIDTH - 1),
		32459 => to_unsigned(971, LUT_AMPL_WIDTH - 1),
		32460 => to_unsigned(967, LUT_AMPL_WIDTH - 1),
		32461 => to_unsigned(964, LUT_AMPL_WIDTH - 1),
		32462 => to_unsigned(961, LUT_AMPL_WIDTH - 1),
		32463 => to_unsigned(958, LUT_AMPL_WIDTH - 1),
		32464 => to_unsigned(955, LUT_AMPL_WIDTH - 1),
		32465 => to_unsigned(952, LUT_AMPL_WIDTH - 1),
		32466 => to_unsigned(949, LUT_AMPL_WIDTH - 1),
		32467 => to_unsigned(945, LUT_AMPL_WIDTH - 1),
		32468 => to_unsigned(942, LUT_AMPL_WIDTH - 1),
		32469 => to_unsigned(939, LUT_AMPL_WIDTH - 1),
		32470 => to_unsigned(936, LUT_AMPL_WIDTH - 1),
		32471 => to_unsigned(933, LUT_AMPL_WIDTH - 1),
		32472 => to_unsigned(930, LUT_AMPL_WIDTH - 1),
		32473 => to_unsigned(927, LUT_AMPL_WIDTH - 1),
		32474 => to_unsigned(923, LUT_AMPL_WIDTH - 1),
		32475 => to_unsigned(920, LUT_AMPL_WIDTH - 1),
		32476 => to_unsigned(917, LUT_AMPL_WIDTH - 1),
		32477 => to_unsigned(914, LUT_AMPL_WIDTH - 1),
		32478 => to_unsigned(911, LUT_AMPL_WIDTH - 1),
		32479 => to_unsigned(908, LUT_AMPL_WIDTH - 1),
		32480 => to_unsigned(905, LUT_AMPL_WIDTH - 1),
		32481 => to_unsigned(901, LUT_AMPL_WIDTH - 1),
		32482 => to_unsigned(898, LUT_AMPL_WIDTH - 1),
		32483 => to_unsigned(895, LUT_AMPL_WIDTH - 1),
		32484 => to_unsigned(892, LUT_AMPL_WIDTH - 1),
		32485 => to_unsigned(889, LUT_AMPL_WIDTH - 1),
		32486 => to_unsigned(886, LUT_AMPL_WIDTH - 1),
		32487 => to_unsigned(883, LUT_AMPL_WIDTH - 1),
		32488 => to_unsigned(880, LUT_AMPL_WIDTH - 1),
		32489 => to_unsigned(876, LUT_AMPL_WIDTH - 1),
		32490 => to_unsigned(873, LUT_AMPL_WIDTH - 1),
		32491 => to_unsigned(870, LUT_AMPL_WIDTH - 1),
		32492 => to_unsigned(867, LUT_AMPL_WIDTH - 1),
		32493 => to_unsigned(864, LUT_AMPL_WIDTH - 1),
		32494 => to_unsigned(861, LUT_AMPL_WIDTH - 1),
		32495 => to_unsigned(858, LUT_AMPL_WIDTH - 1),
		32496 => to_unsigned(854, LUT_AMPL_WIDTH - 1),
		32497 => to_unsigned(851, LUT_AMPL_WIDTH - 1),
		32498 => to_unsigned(848, LUT_AMPL_WIDTH - 1),
		32499 => to_unsigned(845, LUT_AMPL_WIDTH - 1),
		32500 => to_unsigned(842, LUT_AMPL_WIDTH - 1),
		32501 => to_unsigned(839, LUT_AMPL_WIDTH - 1),
		32502 => to_unsigned(836, LUT_AMPL_WIDTH - 1),
		32503 => to_unsigned(832, LUT_AMPL_WIDTH - 1),
		32504 => to_unsigned(829, LUT_AMPL_WIDTH - 1),
		32505 => to_unsigned(826, LUT_AMPL_WIDTH - 1),
		32506 => to_unsigned(823, LUT_AMPL_WIDTH - 1),
		32507 => to_unsigned(820, LUT_AMPL_WIDTH - 1),
		32508 => to_unsigned(817, LUT_AMPL_WIDTH - 1),
		32509 => to_unsigned(814, LUT_AMPL_WIDTH - 1),
		32510 => to_unsigned(810, LUT_AMPL_WIDTH - 1),
		32511 => to_unsigned(807, LUT_AMPL_WIDTH - 1),
		32512 => to_unsigned(804, LUT_AMPL_WIDTH - 1),
		32513 => to_unsigned(801, LUT_AMPL_WIDTH - 1),
		32514 => to_unsigned(798, LUT_AMPL_WIDTH - 1),
		32515 => to_unsigned(795, LUT_AMPL_WIDTH - 1),
		32516 => to_unsigned(792, LUT_AMPL_WIDTH - 1),
		32517 => to_unsigned(788, LUT_AMPL_WIDTH - 1),
		32518 => to_unsigned(785, LUT_AMPL_WIDTH - 1),
		32519 => to_unsigned(782, LUT_AMPL_WIDTH - 1),
		32520 => to_unsigned(779, LUT_AMPL_WIDTH - 1),
		32521 => to_unsigned(776, LUT_AMPL_WIDTH - 1),
		32522 => to_unsigned(773, LUT_AMPL_WIDTH - 1),
		32523 => to_unsigned(770, LUT_AMPL_WIDTH - 1),
		32524 => to_unsigned(766, LUT_AMPL_WIDTH - 1),
		32525 => to_unsigned(763, LUT_AMPL_WIDTH - 1),
		32526 => to_unsigned(760, LUT_AMPL_WIDTH - 1),
		32527 => to_unsigned(757, LUT_AMPL_WIDTH - 1),
		32528 => to_unsigned(754, LUT_AMPL_WIDTH - 1),
		32529 => to_unsigned(751, LUT_AMPL_WIDTH - 1),
		32530 => to_unsigned(748, LUT_AMPL_WIDTH - 1),
		32531 => to_unsigned(744, LUT_AMPL_WIDTH - 1),
		32532 => to_unsigned(741, LUT_AMPL_WIDTH - 1),
		32533 => to_unsigned(738, LUT_AMPL_WIDTH - 1),
		32534 => to_unsigned(735, LUT_AMPL_WIDTH - 1),
		32535 => to_unsigned(732, LUT_AMPL_WIDTH - 1),
		32536 => to_unsigned(729, LUT_AMPL_WIDTH - 1),
		32537 => to_unsigned(726, LUT_AMPL_WIDTH - 1),
		32538 => to_unsigned(722, LUT_AMPL_WIDTH - 1),
		32539 => to_unsigned(719, LUT_AMPL_WIDTH - 1),
		32540 => to_unsigned(716, LUT_AMPL_WIDTH - 1),
		32541 => to_unsigned(713, LUT_AMPL_WIDTH - 1),
		32542 => to_unsigned(710, LUT_AMPL_WIDTH - 1),
		32543 => to_unsigned(707, LUT_AMPL_WIDTH - 1),
		32544 => to_unsigned(704, LUT_AMPL_WIDTH - 1),
		32545 => to_unsigned(701, LUT_AMPL_WIDTH - 1),
		32546 => to_unsigned(697, LUT_AMPL_WIDTH - 1),
		32547 => to_unsigned(694, LUT_AMPL_WIDTH - 1),
		32548 => to_unsigned(691, LUT_AMPL_WIDTH - 1),
		32549 => to_unsigned(688, LUT_AMPL_WIDTH - 1),
		32550 => to_unsigned(685, LUT_AMPL_WIDTH - 1),
		32551 => to_unsigned(682, LUT_AMPL_WIDTH - 1),
		32552 => to_unsigned(679, LUT_AMPL_WIDTH - 1),
		32553 => to_unsigned(675, LUT_AMPL_WIDTH - 1),
		32554 => to_unsigned(672, LUT_AMPL_WIDTH - 1),
		32555 => to_unsigned(669, LUT_AMPL_WIDTH - 1),
		32556 => to_unsigned(666, LUT_AMPL_WIDTH - 1),
		32557 => to_unsigned(663, LUT_AMPL_WIDTH - 1),
		32558 => to_unsigned(660, LUT_AMPL_WIDTH - 1),
		32559 => to_unsigned(657, LUT_AMPL_WIDTH - 1),
		32560 => to_unsigned(653, LUT_AMPL_WIDTH - 1),
		32561 => to_unsigned(650, LUT_AMPL_WIDTH - 1),
		32562 => to_unsigned(647, LUT_AMPL_WIDTH - 1),
		32563 => to_unsigned(644, LUT_AMPL_WIDTH - 1),
		32564 => to_unsigned(641, LUT_AMPL_WIDTH - 1),
		32565 => to_unsigned(638, LUT_AMPL_WIDTH - 1),
		32566 => to_unsigned(635, LUT_AMPL_WIDTH - 1),
		32567 => to_unsigned(631, LUT_AMPL_WIDTH - 1),
		32568 => to_unsigned(628, LUT_AMPL_WIDTH - 1),
		32569 => to_unsigned(625, LUT_AMPL_WIDTH - 1),
		32570 => to_unsigned(622, LUT_AMPL_WIDTH - 1),
		32571 => to_unsigned(619, LUT_AMPL_WIDTH - 1),
		32572 => to_unsigned(616, LUT_AMPL_WIDTH - 1),
		32573 => to_unsigned(613, LUT_AMPL_WIDTH - 1),
		32574 => to_unsigned(609, LUT_AMPL_WIDTH - 1),
		32575 => to_unsigned(606, LUT_AMPL_WIDTH - 1),
		32576 => to_unsigned(603, LUT_AMPL_WIDTH - 1),
		32577 => to_unsigned(600, LUT_AMPL_WIDTH - 1),
		32578 => to_unsigned(597, LUT_AMPL_WIDTH - 1),
		32579 => to_unsigned(594, LUT_AMPL_WIDTH - 1),
		32580 => to_unsigned(591, LUT_AMPL_WIDTH - 1),
		32581 => to_unsigned(587, LUT_AMPL_WIDTH - 1),
		32582 => to_unsigned(584, LUT_AMPL_WIDTH - 1),
		32583 => to_unsigned(581, LUT_AMPL_WIDTH - 1),
		32584 => to_unsigned(578, LUT_AMPL_WIDTH - 1),
		32585 => to_unsigned(575, LUT_AMPL_WIDTH - 1),
		32586 => to_unsigned(572, LUT_AMPL_WIDTH - 1),
		32587 => to_unsigned(569, LUT_AMPL_WIDTH - 1),
		32588 => to_unsigned(565, LUT_AMPL_WIDTH - 1),
		32589 => to_unsigned(562, LUT_AMPL_WIDTH - 1),
		32590 => to_unsigned(559, LUT_AMPL_WIDTH - 1),
		32591 => to_unsigned(556, LUT_AMPL_WIDTH - 1),
		32592 => to_unsigned(553, LUT_AMPL_WIDTH - 1),
		32593 => to_unsigned(550, LUT_AMPL_WIDTH - 1),
		32594 => to_unsigned(547, LUT_AMPL_WIDTH - 1),
		32595 => to_unsigned(543, LUT_AMPL_WIDTH - 1),
		32596 => to_unsigned(540, LUT_AMPL_WIDTH - 1),
		32597 => to_unsigned(537, LUT_AMPL_WIDTH - 1),
		32598 => to_unsigned(534, LUT_AMPL_WIDTH - 1),
		32599 => to_unsigned(531, LUT_AMPL_WIDTH - 1),
		32600 => to_unsigned(528, LUT_AMPL_WIDTH - 1),
		32601 => to_unsigned(525, LUT_AMPL_WIDTH - 1),
		32602 => to_unsigned(521, LUT_AMPL_WIDTH - 1),
		32603 => to_unsigned(518, LUT_AMPL_WIDTH - 1),
		32604 => to_unsigned(515, LUT_AMPL_WIDTH - 1),
		32605 => to_unsigned(512, LUT_AMPL_WIDTH - 1),
		32606 => to_unsigned(509, LUT_AMPL_WIDTH - 1),
		32607 => to_unsigned(506, LUT_AMPL_WIDTH - 1),
		32608 => to_unsigned(503, LUT_AMPL_WIDTH - 1),
		32609 => to_unsigned(499, LUT_AMPL_WIDTH - 1),
		32610 => to_unsigned(496, LUT_AMPL_WIDTH - 1),
		32611 => to_unsigned(493, LUT_AMPL_WIDTH - 1),
		32612 => to_unsigned(490, LUT_AMPL_WIDTH - 1),
		32613 => to_unsigned(487, LUT_AMPL_WIDTH - 1),
		32614 => to_unsigned(484, LUT_AMPL_WIDTH - 1),
		32615 => to_unsigned(481, LUT_AMPL_WIDTH - 1),
		32616 => to_unsigned(477, LUT_AMPL_WIDTH - 1),
		32617 => to_unsigned(474, LUT_AMPL_WIDTH - 1),
		32618 => to_unsigned(471, LUT_AMPL_WIDTH - 1),
		32619 => to_unsigned(468, LUT_AMPL_WIDTH - 1),
		32620 => to_unsigned(465, LUT_AMPL_WIDTH - 1),
		32621 => to_unsigned(462, LUT_AMPL_WIDTH - 1),
		32622 => to_unsigned(459, LUT_AMPL_WIDTH - 1),
		32623 => to_unsigned(456, LUT_AMPL_WIDTH - 1),
		32624 => to_unsigned(452, LUT_AMPL_WIDTH - 1),
		32625 => to_unsigned(449, LUT_AMPL_WIDTH - 1),
		32626 => to_unsigned(446, LUT_AMPL_WIDTH - 1),
		32627 => to_unsigned(443, LUT_AMPL_WIDTH - 1),
		32628 => to_unsigned(440, LUT_AMPL_WIDTH - 1),
		32629 => to_unsigned(437, LUT_AMPL_WIDTH - 1),
		32630 => to_unsigned(434, LUT_AMPL_WIDTH - 1),
		32631 => to_unsigned(430, LUT_AMPL_WIDTH - 1),
		32632 => to_unsigned(427, LUT_AMPL_WIDTH - 1),
		32633 => to_unsigned(424, LUT_AMPL_WIDTH - 1),
		32634 => to_unsigned(421, LUT_AMPL_WIDTH - 1),
		32635 => to_unsigned(418, LUT_AMPL_WIDTH - 1),
		32636 => to_unsigned(415, LUT_AMPL_WIDTH - 1),
		32637 => to_unsigned(412, LUT_AMPL_WIDTH - 1),
		32638 => to_unsigned(408, LUT_AMPL_WIDTH - 1),
		32639 => to_unsigned(405, LUT_AMPL_WIDTH - 1),
		32640 => to_unsigned(402, LUT_AMPL_WIDTH - 1),
		32641 => to_unsigned(399, LUT_AMPL_WIDTH - 1),
		32642 => to_unsigned(396, LUT_AMPL_WIDTH - 1),
		32643 => to_unsigned(393, LUT_AMPL_WIDTH - 1),
		32644 => to_unsigned(390, LUT_AMPL_WIDTH - 1),
		32645 => to_unsigned(386, LUT_AMPL_WIDTH - 1),
		32646 => to_unsigned(383, LUT_AMPL_WIDTH - 1),
		32647 => to_unsigned(380, LUT_AMPL_WIDTH - 1),
		32648 => to_unsigned(377, LUT_AMPL_WIDTH - 1),
		32649 => to_unsigned(374, LUT_AMPL_WIDTH - 1),
		32650 => to_unsigned(371, LUT_AMPL_WIDTH - 1),
		32651 => to_unsigned(368, LUT_AMPL_WIDTH - 1),
		32652 => to_unsigned(364, LUT_AMPL_WIDTH - 1),
		32653 => to_unsigned(361, LUT_AMPL_WIDTH - 1),
		32654 => to_unsigned(358, LUT_AMPL_WIDTH - 1),
		32655 => to_unsigned(355, LUT_AMPL_WIDTH - 1),
		32656 => to_unsigned(352, LUT_AMPL_WIDTH - 1),
		32657 => to_unsigned(349, LUT_AMPL_WIDTH - 1),
		32658 => to_unsigned(346, LUT_AMPL_WIDTH - 1),
		32659 => to_unsigned(342, LUT_AMPL_WIDTH - 1),
		32660 => to_unsigned(339, LUT_AMPL_WIDTH - 1),
		32661 => to_unsigned(336, LUT_AMPL_WIDTH - 1),
		32662 => to_unsigned(333, LUT_AMPL_WIDTH - 1),
		32663 => to_unsigned(330, LUT_AMPL_WIDTH - 1),
		32664 => to_unsigned(327, LUT_AMPL_WIDTH - 1),
		32665 => to_unsigned(324, LUT_AMPL_WIDTH - 1),
		32666 => to_unsigned(320, LUT_AMPL_WIDTH - 1),
		32667 => to_unsigned(317, LUT_AMPL_WIDTH - 1),
		32668 => to_unsigned(314, LUT_AMPL_WIDTH - 1),
		32669 => to_unsigned(311, LUT_AMPL_WIDTH - 1),
		32670 => to_unsigned(308, LUT_AMPL_WIDTH - 1),
		32671 => to_unsigned(305, LUT_AMPL_WIDTH - 1),
		32672 => to_unsigned(302, LUT_AMPL_WIDTH - 1),
		32673 => to_unsigned(298, LUT_AMPL_WIDTH - 1),
		32674 => to_unsigned(295, LUT_AMPL_WIDTH - 1),
		32675 => to_unsigned(292, LUT_AMPL_WIDTH - 1),
		32676 => to_unsigned(289, LUT_AMPL_WIDTH - 1),
		32677 => to_unsigned(286, LUT_AMPL_WIDTH - 1),
		32678 => to_unsigned(283, LUT_AMPL_WIDTH - 1),
		32679 => to_unsigned(280, LUT_AMPL_WIDTH - 1),
		32680 => to_unsigned(276, LUT_AMPL_WIDTH - 1),
		32681 => to_unsigned(273, LUT_AMPL_WIDTH - 1),
		32682 => to_unsigned(270, LUT_AMPL_WIDTH - 1),
		32683 => to_unsigned(267, LUT_AMPL_WIDTH - 1),
		32684 => to_unsigned(264, LUT_AMPL_WIDTH - 1),
		32685 => to_unsigned(261, LUT_AMPL_WIDTH - 1),
		32686 => to_unsigned(258, LUT_AMPL_WIDTH - 1),
		32687 => to_unsigned(254, LUT_AMPL_WIDTH - 1),
		32688 => to_unsigned(251, LUT_AMPL_WIDTH - 1),
		32689 => to_unsigned(248, LUT_AMPL_WIDTH - 1),
		32690 => to_unsigned(245, LUT_AMPL_WIDTH - 1),
		32691 => to_unsigned(242, LUT_AMPL_WIDTH - 1),
		32692 => to_unsigned(239, LUT_AMPL_WIDTH - 1),
		32693 => to_unsigned(236, LUT_AMPL_WIDTH - 1),
		32694 => to_unsigned(232, LUT_AMPL_WIDTH - 1),
		32695 => to_unsigned(229, LUT_AMPL_WIDTH - 1),
		32696 => to_unsigned(226, LUT_AMPL_WIDTH - 1),
		32697 => to_unsigned(223, LUT_AMPL_WIDTH - 1),
		32698 => to_unsigned(220, LUT_AMPL_WIDTH - 1),
		32699 => to_unsigned(217, LUT_AMPL_WIDTH - 1),
		32700 => to_unsigned(214, LUT_AMPL_WIDTH - 1),
		32701 => to_unsigned(210, LUT_AMPL_WIDTH - 1),
		32702 => to_unsigned(207, LUT_AMPL_WIDTH - 1),
		32703 => to_unsigned(204, LUT_AMPL_WIDTH - 1),
		32704 => to_unsigned(201, LUT_AMPL_WIDTH - 1),
		32705 => to_unsigned(198, LUT_AMPL_WIDTH - 1),
		32706 => to_unsigned(195, LUT_AMPL_WIDTH - 1),
		32707 => to_unsigned(192, LUT_AMPL_WIDTH - 1),
		32708 => to_unsigned(188, LUT_AMPL_WIDTH - 1),
		32709 => to_unsigned(185, LUT_AMPL_WIDTH - 1),
		32710 => to_unsigned(182, LUT_AMPL_WIDTH - 1),
		32711 => to_unsigned(179, LUT_AMPL_WIDTH - 1),
		32712 => to_unsigned(176, LUT_AMPL_WIDTH - 1),
		32713 => to_unsigned(173, LUT_AMPL_WIDTH - 1),
		32714 => to_unsigned(170, LUT_AMPL_WIDTH - 1),
		32715 => to_unsigned(166, LUT_AMPL_WIDTH - 1),
		32716 => to_unsigned(163, LUT_AMPL_WIDTH - 1),
		32717 => to_unsigned(160, LUT_AMPL_WIDTH - 1),
		32718 => to_unsigned(157, LUT_AMPL_WIDTH - 1),
		32719 => to_unsigned(154, LUT_AMPL_WIDTH - 1),
		32720 => to_unsigned(151, LUT_AMPL_WIDTH - 1),
		32721 => to_unsigned(148, LUT_AMPL_WIDTH - 1),
		32722 => to_unsigned(145, LUT_AMPL_WIDTH - 1),
		32723 => to_unsigned(141, LUT_AMPL_WIDTH - 1),
		32724 => to_unsigned(138, LUT_AMPL_WIDTH - 1),
		32725 => to_unsigned(135, LUT_AMPL_WIDTH - 1),
		32726 => to_unsigned(132, LUT_AMPL_WIDTH - 1),
		32727 => to_unsigned(129, LUT_AMPL_WIDTH - 1),
		32728 => to_unsigned(126, LUT_AMPL_WIDTH - 1),
		32729 => to_unsigned(123, LUT_AMPL_WIDTH - 1),
		32730 => to_unsigned(119, LUT_AMPL_WIDTH - 1),
		32731 => to_unsigned(116, LUT_AMPL_WIDTH - 1),
		32732 => to_unsigned(113, LUT_AMPL_WIDTH - 1),
		32733 => to_unsigned(110, LUT_AMPL_WIDTH - 1),
		32734 => to_unsigned(107, LUT_AMPL_WIDTH - 1),
		32735 => to_unsigned(104, LUT_AMPL_WIDTH - 1),
		32736 => to_unsigned(101, LUT_AMPL_WIDTH - 1),
		32737 => to_unsigned(97, LUT_AMPL_WIDTH - 1),
		32738 => to_unsigned(94, LUT_AMPL_WIDTH - 1),
		32739 => to_unsigned(91, LUT_AMPL_WIDTH - 1),
		32740 => to_unsigned(88, LUT_AMPL_WIDTH - 1),
		32741 => to_unsigned(85, LUT_AMPL_WIDTH - 1),
		32742 => to_unsigned(82, LUT_AMPL_WIDTH - 1),
		32743 => to_unsigned(79, LUT_AMPL_WIDTH - 1),
		32744 => to_unsigned(75, LUT_AMPL_WIDTH - 1),
		32745 => to_unsigned(72, LUT_AMPL_WIDTH - 1),
		32746 => to_unsigned(69, LUT_AMPL_WIDTH - 1),
		32747 => to_unsigned(66, LUT_AMPL_WIDTH - 1),
		32748 => to_unsigned(63, LUT_AMPL_WIDTH - 1),
		32749 => to_unsigned(60, LUT_AMPL_WIDTH - 1),
		32750 => to_unsigned(57, LUT_AMPL_WIDTH - 1),
		32751 => to_unsigned(53, LUT_AMPL_WIDTH - 1),
		32752 => to_unsigned(50, LUT_AMPL_WIDTH - 1),
		32753 => to_unsigned(47, LUT_AMPL_WIDTH - 1),
		32754 => to_unsigned(44, LUT_AMPL_WIDTH - 1),
		32755 => to_unsigned(41, LUT_AMPL_WIDTH - 1),
		32756 => to_unsigned(38, LUT_AMPL_WIDTH - 1),
		32757 => to_unsigned(35, LUT_AMPL_WIDTH - 1),
		32758 => to_unsigned(31, LUT_AMPL_WIDTH - 1),
		32759 => to_unsigned(28, LUT_AMPL_WIDTH - 1),
		32760 => to_unsigned(25, LUT_AMPL_WIDTH - 1),
		32761 => to_unsigned(22, LUT_AMPL_WIDTH - 1),
		32762 => to_unsigned(19, LUT_AMPL_WIDTH - 1),
		32763 => to_unsigned(16, LUT_AMPL_WIDTH - 1),
		32764 => to_unsigned(13, LUT_AMPL_WIDTH - 1),
		32765 => to_unsigned(9, LUT_AMPL_WIDTH - 1),
		32766 => to_unsigned(6, LUT_AMPL_WIDTH - 1),
		32767 => to_unsigned(3, LUT_AMPL_WIDTH - 1),
		others => to_unsigned(0, LUT_AMPL_WIDTH - 1)
);
end package sine_lut_pkg;

package body sine_lut_pkg is
end package body sine_lut_pkg;
